magic
tech sky130A
magscale 1 2
timestamp 1608703685
<< metal1 >>
rect 58802 700952 58808 701004
rect 58860 700992 58866 701004
rect 202782 700992 202788 701004
rect 58860 700964 202788 700992
rect 58860 700952 58866 700964
rect 202782 700952 202788 700964
rect 202840 700952 202846 701004
rect 58710 700884 58716 700936
rect 58768 700924 58774 700936
rect 218974 700924 218980 700936
rect 58768 700896 218980 700924
rect 58768 700884 58774 700896
rect 218974 700884 218980 700896
rect 219032 700884 219038 700936
rect 58986 700816 58992 700868
rect 59044 700856 59050 700868
rect 267642 700856 267648 700868
rect 59044 700828 267648 700856
rect 59044 700816 59050 700828
rect 267642 700816 267648 700828
rect 267700 700816 267706 700868
rect 58894 700748 58900 700800
rect 58952 700788 58958 700800
rect 283834 700788 283840 700800
rect 58952 700760 283840 700788
rect 58952 700748 58958 700760
rect 283834 700748 283840 700760
rect 283892 700748 283898 700800
rect 59078 700680 59084 700732
rect 59136 700720 59142 700732
rect 332502 700720 332508 700732
rect 59136 700692 332508 700720
rect 59136 700680 59142 700692
rect 332502 700680 332508 700692
rect 332560 700680 332566 700732
rect 57698 700612 57704 700664
rect 57756 700652 57762 700664
rect 348786 700652 348792 700664
rect 57756 700624 348792 700652
rect 57756 700612 57762 700624
rect 348786 700612 348792 700624
rect 348844 700612 348850 700664
rect 59170 700544 59176 700596
rect 59228 700584 59234 700596
rect 397454 700584 397460 700596
rect 59228 700556 397460 700584
rect 59228 700544 59234 700556
rect 397454 700544 397460 700556
rect 397512 700544 397518 700596
rect 57790 700476 57796 700528
rect 57848 700516 57854 700528
rect 413646 700516 413652 700528
rect 57848 700488 413652 700516
rect 57848 700476 57854 700488
rect 413646 700476 413652 700488
rect 413704 700476 413710 700528
rect 57882 700408 57888 700460
rect 57940 700448 57946 700460
rect 478506 700448 478512 700460
rect 57940 700420 478512 700448
rect 57940 700408 57946 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 59262 700340 59268 700392
rect 59320 700380 59326 700392
rect 527174 700380 527180 700392
rect 59320 700352 527180 700380
rect 59320 700340 59326 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 59354 700272 59360 700324
rect 59412 700312 59418 700324
rect 543458 700312 543464 700324
rect 59412 700284 543464 700312
rect 59412 700272 59418 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 58526 700204 58532 700256
rect 58584 700244 58590 700256
rect 136634 700244 136640 700256
rect 58584 700216 136640 700244
rect 58584 700204 58590 700216
rect 136634 700204 136640 700216
rect 136692 700204 136698 700256
rect 137278 700204 137284 700256
rect 137336 700244 137342 700256
rect 235166 700244 235172 700256
rect 137336 700216 235172 700244
rect 137336 700204 137342 700216
rect 235166 700204 235172 700216
rect 235224 700204 235230 700256
rect 57606 700136 57612 700188
rect 57664 700176 57670 700188
rect 154114 700176 154120 700188
rect 57664 700148 154120 700176
rect 57664 700136 57670 700148
rect 154114 700136 154120 700148
rect 154172 700136 154178 700188
rect 57514 700068 57520 700120
rect 57572 700108 57578 700120
rect 89162 700108 89168 700120
rect 57572 700080 89168 700108
rect 57572 700068 57578 700080
rect 89162 700068 89168 700080
rect 89220 700068 89226 700120
rect 136634 700068 136640 700120
rect 136692 700108 136698 700120
rect 137830 700108 137836 700120
rect 136692 700080 137836 700108
rect 136692 700068 136698 700080
rect 137830 700068 137836 700080
rect 137888 700068 137894 700120
rect 58434 700000 58440 700052
rect 58492 700040 58498 700052
rect 72970 700040 72976 700052
rect 58492 700012 72976 700040
rect 58492 700000 58498 700012
rect 72970 700000 72976 700012
rect 73028 700000 73034 700052
rect 40494 699932 40500 699984
rect 40552 699972 40558 699984
rect 42058 699972 42064 699984
rect 40552 699944 42064 699972
rect 40552 699932 40558 699944
rect 42058 699932 42064 699944
rect 42116 699932 42122 699984
rect 8110 699660 8116 699712
rect 8168 699700 8174 699712
rect 10318 699700 10324 699712
rect 8168 699672 10324 699700
rect 8168 699660 8174 699672
rect 10318 699660 10324 699672
rect 10376 699660 10382 699712
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 104986 698232 104992 698284
rect 105044 698272 105050 698284
rect 105538 698272 105544 698284
rect 105044 698244 105544 698272
rect 105044 698232 105050 698244
rect 105538 698232 105544 698244
rect 105596 698232 105602 698284
rect 364426 698232 364432 698284
rect 364484 698272 364490 698284
rect 365070 698272 365076 698284
rect 364484 698244 365076 698272
rect 364484 698232 364490 698244
rect 365070 698232 365076 698244
rect 365128 698232 365134 698284
rect 560294 697280 560300 697332
rect 560352 697320 560358 697332
rect 565170 697320 565176 697332
rect 560352 697292 565176 697320
rect 560352 697280 560358 697292
rect 565170 697280 565176 697292
rect 565228 697280 565234 697332
rect 166902 697144 166908 697196
rect 166960 697184 166966 697196
rect 172422 697184 172428 697196
rect 166960 697156 172428 697184
rect 166960 697144 166966 697156
rect 172422 697144 172428 697156
rect 172480 697144 172486 697196
rect 540974 697144 540980 697196
rect 541032 697184 541038 697196
rect 548610 697184 548616 697196
rect 541032 697156 548616 697184
rect 541032 697144 541038 697156
rect 548610 697144 548616 697156
rect 548668 697144 548674 697196
rect 70302 697076 70308 697128
rect 70360 697116 70366 697128
rect 77202 697116 77208 697128
rect 70360 697088 77208 697116
rect 70360 697076 70366 697088
rect 77202 697076 77208 697088
rect 77260 697076 77266 697128
rect 89622 697076 89628 697128
rect 89680 697116 89686 697128
rect 96522 697116 96528 697128
rect 89680 697088 96528 697116
rect 89680 697076 89686 697088
rect 96522 697076 96528 697088
rect 96580 697076 96586 697128
rect 108942 697076 108948 697128
rect 109000 697116 109006 697128
rect 115842 697116 115848 697128
rect 109000 697088 115848 697116
rect 109000 697076 109006 697088
rect 115842 697076 115848 697088
rect 115900 697076 115906 697128
rect 128262 697076 128268 697128
rect 128320 697116 128326 697128
rect 135162 697116 135168 697128
rect 128320 697088 135168 697116
rect 128320 697076 128326 697088
rect 135162 697076 135168 697088
rect 135220 697076 135226 697128
rect 147582 697076 147588 697128
rect 147640 697116 147646 697128
rect 154482 697116 154488 697128
rect 147640 697088 154488 697116
rect 147640 697076 147646 697088
rect 154482 697076 154488 697088
rect 154540 697076 154546 697128
rect 186222 697076 186228 697128
rect 186280 697116 186286 697128
rect 193122 697116 193128 697128
rect 186280 697088 193128 697116
rect 186280 697076 186286 697088
rect 193122 697076 193128 697088
rect 193180 697076 193186 697128
rect 205542 697076 205548 697128
rect 205600 697116 205606 697128
rect 212442 697116 212448 697128
rect 205600 697088 212448 697116
rect 205600 697076 205606 697088
rect 212442 697076 212448 697088
rect 212500 697076 212506 697128
rect 224862 697076 224868 697128
rect 224920 697116 224926 697128
rect 231762 697116 231768 697128
rect 224920 697088 231768 697116
rect 224920 697076 224926 697088
rect 231762 697076 231768 697088
rect 231820 697076 231826 697128
rect 244182 697076 244188 697128
rect 244240 697116 244246 697128
rect 251082 697116 251088 697128
rect 244240 697088 251088 697116
rect 244240 697076 244246 697088
rect 251082 697076 251088 697088
rect 251140 697076 251146 697128
rect 263502 697076 263508 697128
rect 263560 697116 263566 697128
rect 270402 697116 270408 697128
rect 263560 697088 270408 697116
rect 263560 697076 263566 697088
rect 270402 697076 270408 697088
rect 270460 697076 270466 697128
rect 282822 697076 282828 697128
rect 282880 697116 282886 697128
rect 289722 697116 289728 697128
rect 282880 697088 289728 697116
rect 282880 697076 282886 697088
rect 289722 697076 289728 697088
rect 289780 697076 289786 697128
rect 302142 697076 302148 697128
rect 302200 697116 302206 697128
rect 309042 697116 309048 697128
rect 302200 697088 309048 697116
rect 302200 697076 302206 697088
rect 309042 697076 309048 697088
rect 309100 697076 309106 697128
rect 321462 697076 321468 697128
rect 321520 697116 321526 697128
rect 328362 697116 328368 697128
rect 321520 697088 328368 697116
rect 321520 697076 321526 697088
rect 328362 697076 328368 697088
rect 328420 697076 328426 697128
rect 169754 695444 169760 695496
rect 169812 695484 169818 695496
rect 170030 695484 170036 695496
rect 169812 695456 170036 695484
rect 169812 695444 169818 695456
rect 170030 695444 170036 695456
rect 170088 695444 170094 695496
rect 429194 692792 429200 692844
rect 429252 692832 429258 692844
rect 429930 692832 429936 692844
rect 429252 692804 429936 692832
rect 429252 692792 429258 692804
rect 429930 692792 429936 692804
rect 429988 692792 429994 692844
rect 494054 692792 494060 692844
rect 494112 692832 494118 692844
rect 494882 692832 494888 692844
rect 494112 692804 494888 692832
rect 494112 692792 494118 692804
rect 494882 692792 494888 692804
rect 494940 692792 494946 692844
rect 173894 686264 173900 686316
rect 173952 686304 173958 686316
rect 178770 686304 178776 686316
rect 173952 686276 178776 686304
rect 173952 686264 173958 686276
rect 178770 686264 178776 686276
rect 178828 686264 178834 686316
rect 367094 686264 367100 686316
rect 367152 686304 367158 686316
rect 371970 686304 371976 686316
rect 367152 686276 371976 686304
rect 367152 686264 367158 686276
rect 371970 686264 371976 686276
rect 372028 686264 372034 686316
rect 560294 686264 560300 686316
rect 560352 686304 560358 686316
rect 565170 686304 565176 686316
rect 560352 686276 565176 686304
rect 560352 686264 560358 686276
rect 565170 686264 565176 686276
rect 565228 686264 565234 686316
rect 154574 686128 154580 686180
rect 154632 686168 154638 686180
rect 162210 686168 162216 686180
rect 154632 686140 162216 686168
rect 154632 686128 154638 686140
rect 162210 686128 162216 686140
rect 162268 686128 162274 686180
rect 289814 686128 289820 686180
rect 289872 686168 289878 686180
rect 294506 686168 294512 686180
rect 289872 686140 294512 686168
rect 289872 686128 289878 686140
rect 294506 686128 294512 686140
rect 294564 686128 294570 686180
rect 347774 686128 347780 686180
rect 347832 686168 347838 686180
rect 355410 686168 355416 686180
rect 347832 686140 355416 686168
rect 347832 686128 347838 686140
rect 355410 686128 355416 686140
rect 355468 686128 355474 686180
rect 540974 686128 540980 686180
rect 541032 686168 541038 686180
rect 548610 686168 548616 686180
rect 541032 686140 548616 686168
rect 541032 686128 541038 686140
rect 548610 686128 548616 686140
rect 548668 686128 548674 686180
rect 169754 685856 169760 685908
rect 169812 685896 169818 685908
rect 169938 685896 169944 685908
rect 169812 685868 169944 685896
rect 169812 685856 169818 685868
rect 169938 685856 169944 685868
rect 169996 685856 170002 685908
rect 299566 685856 299572 685908
rect 299624 685896 299630 685908
rect 300118 685896 300124 685908
rect 299624 685868 300124 685896
rect 299624 685856 299630 685868
rect 300118 685856 300124 685868
rect 300176 685856 300182 685908
rect 559006 684496 559012 684548
rect 559064 684536 559070 684548
rect 559650 684536 559656 684548
rect 559064 684508 559656 684536
rect 559064 684496 559070 684508
rect 559650 684496 559656 684508
rect 559708 684496 559714 684548
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299658 684468 299664 684480
rect 299624 684440 299664 684468
rect 299624 684428 299630 684440
rect 299658 684428 299664 684440
rect 299716 684428 299722 684480
rect 2774 681708 2780 681760
rect 2832 681748 2838 681760
rect 5074 681748 5080 681760
rect 2832 681720 5080 681748
rect 2832 681708 2838 681720
rect 5074 681708 5080 681720
rect 5132 681708 5138 681760
rect 299658 679028 299664 679040
rect 299584 679000 299664 679028
rect 299584 678972 299612 679000
rect 299658 678988 299664 679000
rect 299716 678988 299722 679040
rect 299566 678920 299572 678972
rect 299624 678920 299630 678972
rect 429194 676132 429200 676184
rect 429252 676172 429258 676184
rect 429286 676172 429292 676184
rect 429252 676144 429292 676172
rect 429252 676132 429258 676144
rect 429286 676132 429292 676144
rect 429344 676132 429350 676184
rect 559006 674840 559012 674892
rect 559064 674880 559070 674892
rect 559374 674880 559380 674892
rect 559064 674852 559380 674880
rect 559064 674840 559070 674852
rect 559374 674840 559380 674852
rect 559432 674840 559438 674892
rect 173894 673888 173900 673940
rect 173952 673928 173958 673940
rect 178770 673928 178776 673940
rect 173952 673900 178776 673928
rect 173952 673888 173958 673900
rect 178770 673888 178776 673900
rect 178828 673888 178834 673940
rect 367094 673888 367100 673940
rect 367152 673928 367158 673940
rect 371970 673928 371976 673940
rect 367152 673900 371976 673928
rect 367152 673888 367158 673900
rect 371970 673888 371976 673900
rect 372028 673888 372034 673940
rect 560294 673888 560300 673940
rect 560352 673928 560358 673940
rect 565170 673928 565176 673940
rect 560352 673900 565176 673928
rect 560352 673888 560358 673900
rect 565170 673888 565176 673900
rect 565228 673888 565234 673940
rect 154574 673752 154580 673804
rect 154632 673792 154638 673804
rect 162210 673792 162216 673804
rect 154632 673764 162216 673792
rect 154632 673752 154638 673764
rect 162210 673752 162216 673764
rect 162268 673752 162274 673804
rect 289814 673752 289820 673804
rect 289872 673792 289878 673804
rect 292666 673792 292672 673804
rect 289872 673764 292672 673792
rect 289872 673752 289878 673764
rect 292666 673752 292672 673764
rect 292724 673752 292730 673804
rect 347774 673752 347780 673804
rect 347832 673792 347838 673804
rect 355410 673792 355416 673804
rect 347832 673764 355416 673792
rect 347832 673752 347838 673764
rect 355410 673752 355416 673764
rect 355468 673752 355474 673804
rect 540974 673752 540980 673804
rect 541032 673792 541038 673804
rect 548610 673792 548616 673804
rect 541032 673764 548616 673792
rect 541032 673752 541038 673764
rect 548610 673752 548616 673764
rect 548668 673752 548674 673804
rect 104894 673480 104900 673532
rect 104952 673520 104958 673532
rect 105078 673520 105084 673532
rect 104952 673492 105084 673520
rect 104952 673480 104958 673492
rect 105078 673480 105084 673492
rect 105136 673480 105142 673532
rect 494054 673480 494060 673532
rect 494112 673520 494118 673532
rect 494238 673520 494244 673532
rect 494112 673492 494244 673520
rect 494112 673480 494118 673492
rect 494238 673480 494244 673492
rect 494296 673480 494302 673532
rect 364426 669400 364432 669452
rect 364484 669400 364490 669452
rect 364444 669316 364472 669400
rect 364426 669264 364432 669316
rect 364484 669264 364490 669316
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 21358 667944 21364 667956
rect 3476 667916 21364 667944
rect 3476 667904 3482 667916
rect 21358 667904 21364 667916
rect 21416 667904 21422 667956
rect 299566 666544 299572 666596
rect 299624 666584 299630 666596
rect 299750 666584 299756 666596
rect 299624 666556 299756 666584
rect 299624 666544 299630 666556
rect 299750 666544 299756 666556
rect 299808 666544 299814 666596
rect 429286 666544 429292 666596
rect 429344 666584 429350 666596
rect 429378 666584 429384 666596
rect 429344 666556 429384 666584
rect 429344 666544 429350 666556
rect 429378 666544 429384 666556
rect 429436 666544 429442 666596
rect 559098 661716 559104 661768
rect 559156 661756 559162 661768
rect 559374 661756 559380 661768
rect 559156 661728 559380 661756
rect 559156 661716 559162 661728
rect 559374 661716 559380 661728
rect 559432 661716 559438 661768
rect 170030 659716 170036 659728
rect 169956 659688 170036 659716
rect 169956 659660 169984 659688
rect 170030 659676 170036 659688
rect 170088 659676 170094 659728
rect 299750 659716 299756 659728
rect 299584 659688 299756 659716
rect 299584 659660 299612 659688
rect 299750 659676 299756 659688
rect 299808 659676 299814 659728
rect 429378 659716 429384 659728
rect 429304 659688 429384 659716
rect 429304 659660 429332 659688
rect 429378 659676 429384 659688
rect 429436 659676 429442 659728
rect 169938 659608 169944 659660
rect 169996 659608 170002 659660
rect 299566 659608 299572 659660
rect 299624 659608 299630 659660
rect 429286 659608 429292 659660
rect 429344 659608 429350 659660
rect 559098 656888 559104 656940
rect 559156 656928 559162 656940
rect 559190 656928 559196 656940
rect 559156 656900 559196 656928
rect 559156 656888 559162 656900
rect 559190 656888 559196 656900
rect 559248 656888 559254 656940
rect 169754 655460 169760 655512
rect 169812 655500 169818 655512
rect 169938 655500 169944 655512
rect 169812 655472 169944 655500
rect 169812 655460 169818 655472
rect 169938 655460 169944 655472
rect 169996 655460 170002 655512
rect 104894 654100 104900 654152
rect 104952 654140 104958 654152
rect 105078 654140 105084 654152
rect 104952 654112 105084 654140
rect 104952 654100 104958 654112
rect 105078 654100 105084 654112
rect 105136 654100 105142 654152
rect 364334 654100 364340 654152
rect 364392 654140 364398 654152
rect 364518 654140 364524 654152
rect 364392 654112 364524 654140
rect 364392 654100 364398 654112
rect 364518 654100 364524 654112
rect 364576 654100 364582 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 507854 653352 507860 653404
rect 507912 653392 507918 653404
rect 513374 653392 513380 653404
rect 507912 653364 513380 653392
rect 507912 653352 507918 653364
rect 513374 653352 513380 653364
rect 513432 653352 513438 653404
rect 513374 652808 513380 652860
rect 513432 652848 513438 652860
rect 518894 652848 518900 652860
rect 513432 652820 518900 652848
rect 513432 652808 513438 652820
rect 518894 652808 518900 652820
rect 518952 652808 518958 652860
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 13078 652780 13084 652792
rect 3108 652752 13084 652780
rect 3108 652740 3114 652752
rect 13078 652740 13084 652752
rect 13136 652740 13142 652792
rect 129274 652740 129280 652792
rect 129332 652780 129338 652792
rect 133598 652780 133604 652792
rect 129332 652752 133604 652780
rect 129332 652740 129338 652752
rect 133598 652740 133604 652752
rect 133656 652780 133662 652792
rect 139578 652780 139584 652792
rect 133656 652752 139584 652780
rect 133656 652740 133662 652752
rect 139578 652740 139584 652752
rect 139636 652780 139642 652792
rect 259178 652780 259184 652792
rect 139636 652752 259184 652780
rect 139636 652740 139642 652752
rect 259178 652740 259184 652752
rect 259236 652780 259242 652792
rect 263778 652780 263784 652792
rect 259236 652752 263784 652780
rect 259236 652740 259242 652752
rect 263778 652740 263784 652752
rect 263836 652780 263842 652792
rect 269114 652780 269120 652792
rect 263836 652752 269120 652780
rect 263836 652740 263842 652752
rect 269114 652740 269120 652752
rect 269172 652780 269178 652792
rect 378502 652780 378508 652792
rect 269172 652752 378508 652780
rect 269172 652740 269178 652752
rect 378502 652740 378508 652752
rect 378560 652780 378566 652792
rect 383470 652780 383476 652792
rect 378560 652752 383476 652780
rect 378560 652740 378566 652752
rect 383470 652740 383476 652752
rect 383528 652780 383534 652792
rect 389358 652780 389364 652792
rect 383528 652752 389364 652780
rect 383528 652740 383534 652752
rect 389358 652740 389364 652752
rect 389416 652780 389422 652792
rect 507854 652780 507860 652792
rect 389416 652752 507860 652780
rect 389416 652740 389422 652752
rect 507854 652740 507860 652752
rect 507912 652740 507918 652792
rect 57422 650836 57428 650888
rect 57480 650876 57486 650888
rect 104894 650876 104900 650888
rect 57480 650848 104900 650876
rect 57480 650836 57486 650848
rect 104894 650836 104900 650848
rect 104952 650836 104958 650888
rect 59538 650768 59544 650820
rect 59596 650808 59602 650820
rect 364334 650808 364340 650820
rect 59596 650780 364340 650808
rect 59596 650768 59602 650780
rect 364334 650768 364340 650780
rect 364392 650768 364398 650820
rect 58342 650700 58348 650752
rect 58400 650740 58406 650752
rect 462314 650740 462320 650752
rect 58400 650712 462320 650740
rect 58400 650700 58406 650712
rect 462314 650700 462320 650712
rect 462372 650700 462378 650752
rect 59446 650632 59452 650684
rect 59504 650672 59510 650684
rect 494054 650672 494060 650684
rect 59504 650644 494060 650672
rect 59504 650632 59510 650644
rect 494054 650632 494060 650644
rect 494112 650632 494118 650684
rect 139394 650360 139400 650412
rect 139452 650400 139458 650412
rect 266354 650400 266360 650412
rect 139452 650372 266360 650400
rect 139452 650360 139458 650372
rect 266354 650360 266360 650372
rect 266412 650360 266418 650412
rect 281994 650360 282000 650412
rect 282052 650400 282058 650412
rect 389174 650400 389180 650412
rect 282052 650372 389180 650400
rect 282052 650360 282058 650372
rect 389174 650360 389180 650372
rect 389232 650400 389238 650412
rect 516410 650400 516416 650412
rect 389232 650372 516416 650400
rect 389232 650360 389238 650372
rect 516410 650360 516416 650372
rect 516468 650360 516474 650412
rect 58618 650292 58624 650344
rect 58676 650332 58682 650344
rect 580166 650332 580172 650344
rect 58676 650304 580172 650332
rect 58676 650292 58682 650304
rect 580166 650292 580172 650304
rect 580224 650292 580230 650344
rect 266354 650020 266360 650072
rect 266412 650060 266418 650072
rect 281534 650060 281540 650072
rect 266412 650032 281540 650060
rect 266412 650020 266418 650032
rect 281534 650020 281540 650032
rect 281592 650060 281598 650072
rect 281994 650060 282000 650072
rect 281592 650032 282000 650060
rect 281592 650020 281598 650032
rect 281994 650020 282000 650032
rect 282052 650020 282058 650072
rect 299566 649952 299572 650004
rect 299624 649992 299630 650004
rect 299750 649992 299756 650004
rect 299624 649964 299756 649992
rect 299624 649952 299630 649964
rect 299750 649952 299756 649964
rect 299808 649952 299814 650004
rect 429286 649952 429292 650004
rect 429344 649992 429350 650004
rect 429470 649992 429476 650004
rect 429344 649964 429476 649992
rect 429344 649952 429350 649964
rect 429470 649952 429476 649964
rect 429528 649952 429534 650004
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 142062 645872 142068 645924
rect 142120 645912 142126 645924
rect 187694 645912 187700 645924
rect 142120 645884 187700 645912
rect 142120 645872 142126 645884
rect 187694 645872 187700 645884
rect 187752 645872 187758 645924
rect 291930 645872 291936 645924
rect 291988 645912 291994 645924
rect 307386 645912 307392 645924
rect 291988 645884 307392 645912
rect 291988 645872 291994 645884
rect 307386 645872 307392 645884
rect 307444 645872 307450 645924
rect 399478 645872 399484 645924
rect 399536 645912 399542 645924
rect 437474 645912 437480 645924
rect 399536 645884 437480 645912
rect 399536 645872 399542 645884
rect 437474 645872 437480 645884
rect 437532 645872 437538 645924
rect 140682 644444 140688 644496
rect 140740 644484 140746 644496
rect 187694 644484 187700 644496
rect 140740 644456 187700 644484
rect 140740 644444 140746 644456
rect 187694 644444 187700 644456
rect 187752 644444 187758 644496
rect 290550 644444 290556 644496
rect 290608 644484 290614 644496
rect 307110 644484 307116 644496
rect 290608 644456 307116 644484
rect 290608 644444 290614 644456
rect 307110 644444 307116 644456
rect 307168 644444 307174 644496
rect 398098 644444 398104 644496
rect 398156 644484 398162 644496
rect 437474 644484 437480 644496
rect 398156 644456 437480 644484
rect 398156 644444 398162 644456
rect 437474 644444 437480 644456
rect 437532 644444 437538 644496
rect 137922 643084 137928 643136
rect 137980 643124 137986 643136
rect 187694 643124 187700 643136
rect 137980 643096 187700 643124
rect 137980 643084 137986 643096
rect 187694 643084 187700 643096
rect 187752 643084 187758 643136
rect 287698 643084 287704 643136
rect 287756 643124 287762 643136
rect 307110 643124 307116 643136
rect 287756 643096 307116 643124
rect 287756 643084 287762 643096
rect 307110 643084 307116 643096
rect 307168 643084 307174 643136
rect 395338 643084 395344 643136
rect 395396 643124 395402 643136
rect 437474 643124 437480 643136
rect 395396 643096 437480 643124
rect 395396 643084 395402 643096
rect 437474 643084 437480 643096
rect 437532 643084 437538 643136
rect 299474 642336 299480 642388
rect 299532 642376 299538 642388
rect 299750 642376 299756 642388
rect 299532 642348 299756 642376
rect 299532 642336 299538 642348
rect 299750 642336 299756 642348
rect 299808 642336 299814 642388
rect 160738 641724 160744 641776
rect 160796 641764 160802 641776
rect 187694 641764 187700 641776
rect 160796 641736 187700 641764
rect 160796 641724 160802 641736
rect 187694 641724 187700 641736
rect 187752 641724 187758 641776
rect 286318 641724 286324 641776
rect 286376 641764 286382 641776
rect 307662 641764 307668 641776
rect 286376 641736 307668 641764
rect 286376 641724 286382 641736
rect 307662 641724 307668 641736
rect 307720 641724 307726 641776
rect 393958 641724 393964 641776
rect 394016 641764 394022 641776
rect 437474 641764 437480 641776
rect 394016 641736 437480 641764
rect 394016 641724 394022 641736
rect 437474 641724 437480 641736
rect 437532 641724 437538 641776
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 159358 640296 159364 640348
rect 159416 640336 159422 640348
rect 187694 640336 187700 640348
rect 159416 640308 187700 640336
rect 159416 640296 159422 640308
rect 187694 640296 187700 640308
rect 187752 640296 187758 640348
rect 284938 640296 284944 640348
rect 284996 640336 285002 640348
rect 307662 640336 307668 640348
rect 284996 640308 307668 640336
rect 284996 640296 285002 640308
rect 307662 640296 307668 640308
rect 307720 640296 307726 640348
rect 392578 640296 392584 640348
rect 392636 640336 392642 640348
rect 437474 640336 437480 640348
rect 392636 640308 437480 640336
rect 392636 640296 392642 640308
rect 437474 640296 437480 640308
rect 437532 640296 437538 640348
rect 283558 638936 283564 638988
rect 283616 638976 283622 638988
rect 306650 638976 306656 638988
rect 283616 638948 306656 638976
rect 283616 638936 283622 638948
rect 306650 638936 306656 638948
rect 306708 638936 306714 638988
rect 391198 638936 391204 638988
rect 391256 638976 391262 638988
rect 437474 638976 437480 638988
rect 391256 638948 437480 638976
rect 391256 638936 391262 638948
rect 437474 638936 437480 638948
rect 437532 638936 437538 638988
rect 299474 637644 299480 637696
rect 299532 637684 299538 637696
rect 299532 637656 299704 637684
rect 299532 637644 299538 637656
rect 299676 637628 299704 637656
rect 425072 637656 429516 637684
rect 294598 637576 294604 637628
rect 294656 637616 294662 637628
rect 299566 637616 299572 637628
rect 294656 637588 299572 637616
rect 294656 637576 294662 637588
rect 299566 637576 299572 637588
rect 299624 637576 299630 637628
rect 299658 637576 299664 637628
rect 299716 637576 299722 637628
rect 388438 637576 388444 637628
rect 388496 637616 388502 637628
rect 425072 637616 425100 637656
rect 388496 637588 425100 637616
rect 429488 637616 429516 637656
rect 437474 637616 437480 637628
rect 429488 637588 437480 637616
rect 388496 637576 388502 637588
rect 437474 637576 437480 637588
rect 437532 637576 437538 637628
rect 429194 637508 429200 637560
rect 429252 637548 429258 637560
rect 429378 637548 429384 637560
rect 429252 637520 429384 637548
rect 429252 637508 429258 637520
rect 429378 637508 429384 637520
rect 429436 637508 429442 637560
rect 169662 636216 169668 636268
rect 169720 636256 169726 636268
rect 169938 636256 169944 636268
rect 169720 636228 169944 636256
rect 169720 636216 169726 636228
rect 169938 636216 169944 636228
rect 169996 636216 170002 636268
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 169662 627920 169668 627972
rect 169720 627960 169726 627972
rect 170030 627960 170036 627972
rect 169720 627932 170036 627960
rect 169720 627920 169726 627932
rect 170030 627920 170036 627932
rect 170088 627920 170094 627972
rect 299842 627920 299848 627972
rect 299900 627960 299906 627972
rect 300026 627960 300032 627972
rect 299900 627932 300032 627960
rect 299900 627920 299906 627932
rect 300026 627920 300032 627932
rect 300084 627920 300090 627972
rect 429194 627920 429200 627972
rect 429252 627960 429258 627972
rect 429562 627960 429568 627972
rect 429252 627932 429568 627960
rect 429252 627920 429258 627932
rect 429562 627920 429568 627932
rect 429620 627920 429626 627972
rect 3878 623772 3884 623824
rect 3936 623812 3942 623824
rect 5166 623812 5172 623824
rect 3936 623784 5172 623812
rect 3936 623772 3942 623784
rect 5166 623772 5172 623784
rect 5224 623772 5230 623824
rect 299842 621092 299848 621104
rect 299768 621064 299848 621092
rect 299768 620968 299796 621064
rect 299842 621052 299848 621064
rect 299900 621052 299906 621104
rect 429562 621092 429568 621104
rect 429488 621064 429568 621092
rect 429488 620968 429516 621064
rect 429562 621052 429568 621064
rect 429620 621052 429626 621104
rect 299750 620916 299756 620968
rect 299808 620916 299814 620968
rect 429470 620916 429476 620968
rect 429528 620916 429534 620968
rect 169846 618264 169852 618316
rect 169904 618304 169910 618316
rect 170030 618304 170036 618316
rect 169904 618276 170036 618304
rect 169904 618264 169910 618276
rect 170030 618264 170036 618276
rect 170088 618264 170094 618316
rect 169938 611396 169944 611448
rect 169996 611436 170002 611448
rect 169996 611408 170076 611436
rect 169996 611396 170002 611408
rect 170048 611244 170076 611408
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 170030 611192 170036 611244
rect 170088 611192 170094 611244
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 31018 610008 31024 610020
rect 3476 609980 31024 610008
rect 3476 609968 3482 609980
rect 31018 609968 31024 609980
rect 31076 609968 31082 610020
rect 299566 608540 299572 608592
rect 299624 608580 299630 608592
rect 299658 608580 299664 608592
rect 299624 608552 299664 608580
rect 299624 608540 299630 608552
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 429286 608540 429292 608592
rect 429344 608580 429350 608592
rect 429378 608580 429384 608592
rect 429344 608552 429384 608580
rect 429344 608540 429350 608552
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559006 608540 559012 608592
rect 559064 608580 559070 608592
rect 559098 608580 559104 608592
rect 559064 608552 559104 608580
rect 559064 608540 559070 608552
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 299566 601672 299572 601724
rect 299624 601712 299630 601724
rect 299842 601712 299848 601724
rect 299624 601684 299848 601712
rect 299624 601672 299630 601684
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 429286 601672 429292 601724
rect 429344 601712 429350 601724
rect 429562 601712 429568 601724
rect 429344 601684 429568 601712
rect 429344 601672 429350 601684
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559006 601672 559012 601724
rect 559064 601712 559070 601724
rect 559282 601712 559288 601724
rect 559064 601684 559288 601712
rect 559064 601672 559070 601684
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 169846 598952 169852 599004
rect 169904 598992 169910 599004
rect 170030 598992 170036 599004
rect 169904 598964 170036 598992
rect 169904 598952 169910 598964
rect 170030 598952 170036 598964
rect 170088 598952 170094 599004
rect 299658 598884 299664 598936
rect 299716 598924 299722 598936
rect 299842 598924 299848 598936
rect 299716 598896 299848 598924
rect 299716 598884 299722 598896
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 429378 598884 429384 598936
rect 429436 598924 429442 598936
rect 429562 598924 429568 598936
rect 429436 598896 429568 598924
rect 429436 598884 429442 598896
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559098 598884 559104 598936
rect 559156 598924 559162 598936
rect 559282 598924 559288 598936
rect 559156 598896 559288 598924
rect 559156 598884 559162 598896
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 14458 594844 14464 594856
rect 3292 594816 14464 594844
rect 3292 594804 3298 594816
rect 14458 594804 14464 594816
rect 14516 594804 14522 594856
rect 169938 592084 169944 592136
rect 169996 592124 170002 592136
rect 169996 592096 170076 592124
rect 169996 592084 170002 592096
rect 170048 591932 170076 592096
rect 170030 591880 170036 591932
rect 170088 591880 170094 591932
rect 299658 589296 299664 589348
rect 299716 589336 299722 589348
rect 299934 589336 299940 589348
rect 299716 589308 299940 589336
rect 299716 589296 299722 589308
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 429378 589296 429384 589348
rect 429436 589336 429442 589348
rect 429654 589336 429660 589348
rect 429436 589308 429660 589336
rect 429436 589296 429442 589308
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559098 589296 559104 589348
rect 559156 589336 559162 589348
rect 559374 589336 559380 589348
rect 559156 589308 559380 589336
rect 559156 589296 559162 589308
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 429654 582468 429660 582480
rect 429580 582440 429660 582468
rect 429580 582344 429608 582440
rect 429654 582428 429660 582440
rect 429712 582428 429718 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 429562 582292 429568 582344
rect 429620 582292 429626 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 270034 580252 270040 580304
rect 270092 580292 270098 580304
rect 281626 580292 281632 580304
rect 270092 580264 281632 580292
rect 270092 580252 270098 580264
rect 281626 580252 281632 580264
rect 281684 580252 281690 580304
rect 177942 579640 177948 579692
rect 178000 579680 178006 579692
rect 187694 579680 187700 579692
rect 178000 579652 187700 579680
rect 178000 579640 178006 579652
rect 187694 579640 187700 579652
rect 187752 579640 187758 579692
rect 285030 579640 285036 579692
rect 285088 579680 285094 579692
rect 306926 579680 306932 579692
rect 285088 579652 306932 579680
rect 285088 579640 285094 579652
rect 306926 579640 306932 579652
rect 306984 579640 306990 579692
rect 402238 579640 402244 579692
rect 402296 579680 402302 579692
rect 437474 579680 437480 579692
rect 402296 579652 437480 579680
rect 402296 579640 402302 579652
rect 437474 579640 437480 579652
rect 437532 579640 437538 579692
rect 170122 578212 170128 578264
rect 170180 578252 170186 578264
rect 170306 578252 170312 578264
rect 170180 578224 170312 578252
rect 170180 578212 170186 578224
rect 170306 578212 170312 578224
rect 170364 578212 170370 578264
rect 282178 578212 282184 578264
rect 282236 578252 282242 578264
rect 306374 578252 306380 578264
rect 282236 578224 306380 578252
rect 282236 578212 282242 578224
rect 306374 578212 306380 578224
rect 306432 578212 306438 578264
rect 170122 572704 170128 572756
rect 170180 572704 170186 572756
rect 170140 572620 170168 572704
rect 170122 572568 170128 572620
rect 170180 572568 170186 572620
rect 3970 567196 3976 567248
rect 4028 567236 4034 567248
rect 5258 567236 5264 567248
rect 4028 567208 5264 567236
rect 4028 567196 4034 567208
rect 5258 567196 5264 567208
rect 5316 567196 5322 567248
rect 170122 563156 170128 563168
rect 170048 563128 170128 563156
rect 170048 563032 170076 563128
rect 170122 563116 170128 563128
rect 170180 563116 170186 563168
rect 170030 562980 170036 563032
rect 170088 562980 170094 563032
rect 281718 561620 281724 561672
rect 281776 561660 281782 561672
rect 282178 561660 282184 561672
rect 281776 561632 282184 561660
rect 281776 561620 281782 561632
rect 282178 561620 282184 561632
rect 282236 561620 282242 561672
rect 59630 560872 59636 560924
rect 59688 560912 59694 560924
rect 188982 560912 188988 560924
rect 59688 560884 188988 560912
rect 59688 560872 59694 560884
rect 188982 560872 188988 560884
rect 189040 560912 189046 560924
rect 281718 560912 281724 560924
rect 189040 560884 281724 560912
rect 189040 560872 189046 560884
rect 281718 560872 281724 560884
rect 281776 560872 281782 560924
rect 306282 560872 306288 560924
rect 306340 560912 306346 560924
rect 438118 560912 438124 560924
rect 306340 560884 438124 560912
rect 306340 560872 306346 560884
rect 438118 560872 438124 560884
rect 438176 560872 438182 560924
rect 559006 560260 559012 560312
rect 559064 560300 559070 560312
rect 559098 560300 559104 560312
rect 559064 560272 559104 560300
rect 559064 560260 559070 560272
rect 559098 560260 559104 560272
rect 559156 560260 559162 560312
rect 79318 558832 79324 558884
rect 79376 558872 79382 558884
rect 81434 558872 81440 558884
rect 79376 558844 81440 558872
rect 79376 558832 79382 558844
rect 81434 558832 81440 558844
rect 81492 558832 81498 558884
rect 81526 558832 81532 558884
rect 81584 558872 81590 558884
rect 86862 558872 86868 558884
rect 81584 558844 86868 558872
rect 81584 558832 81590 558844
rect 86862 558832 86868 558844
rect 86920 558832 86926 558884
rect 90082 558872 90088 558884
rect 87800 558844 90088 558872
rect 80698 558764 80704 558816
rect 80756 558804 80762 558816
rect 87800 558804 87828 558844
rect 90082 558832 90088 558844
rect 90140 558872 90146 558884
rect 91002 558872 91008 558884
rect 90140 558844 91008 558872
rect 90140 558832 90146 558844
rect 91002 558832 91008 558844
rect 91060 558832 91066 558884
rect 335446 558832 335452 558884
rect 335504 558872 335510 558884
rect 344278 558872 344284 558884
rect 335504 558844 344284 558872
rect 335504 558832 335510 558844
rect 344278 558832 344284 558844
rect 344336 558832 344342 558884
rect 355318 558832 355324 558884
rect 355376 558872 355382 558884
rect 483014 558872 483020 558884
rect 355376 558844 483020 558872
rect 355376 558832 355382 558844
rect 483014 558832 483020 558844
rect 483072 558832 483078 558884
rect 80756 558776 87828 558804
rect 80756 558764 80762 558776
rect 87874 558764 87880 558816
rect 87932 558804 87938 558816
rect 96614 558804 96620 558816
rect 87932 558776 96620 558804
rect 87932 558764 87938 558776
rect 96614 558764 96620 558776
rect 96672 558764 96678 558816
rect 223574 558764 223580 558816
rect 223632 558804 223638 558816
rect 231946 558804 231952 558816
rect 223632 558776 231952 558804
rect 223632 558764 223638 558776
rect 231946 558764 231952 558776
rect 232004 558764 232010 558816
rect 343726 558764 343732 558816
rect 343784 558804 343790 558816
rect 351914 558804 351920 558816
rect 343784 558776 351920 558804
rect 343784 558764 343790 558776
rect 351914 558764 351920 558776
rect 351972 558764 351978 558816
rect 458818 558764 458824 558816
rect 458876 558804 458882 558816
rect 468018 558804 468024 558816
rect 458876 558776 468024 558804
rect 458876 558764 458882 558776
rect 468018 558764 468024 558776
rect 468076 558804 468082 558816
rect 477126 558804 477132 558816
rect 468076 558776 477132 558804
rect 468076 558764 468082 558776
rect 477126 558764 477132 558776
rect 477184 558804 477190 558816
rect 485774 558804 485780 558816
rect 477184 558776 485780 558804
rect 477184 558764 477190 558776
rect 485774 558764 485780 558776
rect 485832 558764 485838 558816
rect 79502 558696 79508 558748
rect 79560 558736 79566 558748
rect 88978 558736 88984 558748
rect 79560 558708 88984 558736
rect 79560 558696 79566 558708
rect 88978 558696 88984 558708
rect 89036 558696 89042 558748
rect 100294 558736 100300 558748
rect 93504 558708 100300 558736
rect 77386 558628 77392 558680
rect 77444 558668 77450 558680
rect 81526 558668 81532 558680
rect 77444 558640 81532 558668
rect 77444 558628 77450 558640
rect 81526 558628 81532 558640
rect 81584 558628 81590 558680
rect 81618 558628 81624 558680
rect 81676 558668 81682 558680
rect 91370 558668 91376 558680
rect 81676 558640 91376 558668
rect 81676 558628 81682 558640
rect 91370 558628 91376 558640
rect 91428 558668 91434 558680
rect 93504 558668 93532 558708
rect 100294 558696 100300 558708
rect 100352 558696 100358 558748
rect 216766 558696 216772 558748
rect 216824 558736 216830 558748
rect 225782 558736 225788 558748
rect 216824 558708 225788 558736
rect 216824 558696 216830 558708
rect 225782 558696 225788 558708
rect 225840 558696 225846 558748
rect 226334 558696 226340 558748
rect 226392 558736 226398 558748
rect 227162 558736 227168 558748
rect 226392 558708 227168 558736
rect 226392 558696 226398 558708
rect 227162 558696 227168 558708
rect 227220 558736 227226 558748
rect 235994 558736 236000 558748
rect 227220 558708 236000 558736
rect 227220 558696 227226 558708
rect 235994 558696 236000 558708
rect 236052 558696 236058 558748
rect 344278 558696 344284 558748
rect 344336 558736 344342 558748
rect 353294 558736 353300 558748
rect 344336 558708 353300 558736
rect 344336 558696 344342 558708
rect 353294 558696 353300 558708
rect 353352 558696 353358 558748
rect 460658 558696 460664 558748
rect 460716 558736 460722 558748
rect 468570 558736 468576 558748
rect 460716 558708 468576 558736
rect 460716 558696 460722 558708
rect 468570 558696 468576 558708
rect 468628 558696 468634 558748
rect 475562 558696 475568 558748
rect 475620 558736 475626 558748
rect 484394 558736 484400 558748
rect 475620 558708 484400 558736
rect 475620 558696 475626 558708
rect 484394 558696 484400 558708
rect 484452 558696 484458 558748
rect 91428 558640 93532 558668
rect 91428 558628 91434 558640
rect 95326 558628 95332 558680
rect 95384 558668 95390 558680
rect 105354 558668 105360 558680
rect 95384 558640 105360 558668
rect 95384 558628 95390 558640
rect 105354 558628 105360 558640
rect 105412 558668 105418 558680
rect 106090 558668 106096 558680
rect 105412 558640 106096 558668
rect 105412 558628 105418 558640
rect 106090 558628 106096 558640
rect 106148 558628 106154 558680
rect 215294 558628 215300 558680
rect 215352 558668 215358 558680
rect 224402 558668 224408 558680
rect 215352 558640 224408 558668
rect 215352 558628 215358 558640
rect 224402 558628 224408 558640
rect 224460 558668 224466 558680
rect 233234 558668 233240 558680
rect 224460 558640 233240 558668
rect 224460 558628 224466 558640
rect 233234 558628 233240 558640
rect 233292 558628 233298 558680
rect 338942 558628 338948 558680
rect 339000 558668 339006 558680
rect 348326 558668 348332 558680
rect 339000 558640 348332 558668
rect 339000 558628 339006 558640
rect 348326 558628 348332 558640
rect 348384 558668 348390 558680
rect 357434 558668 357440 558680
rect 348384 558640 357440 558668
rect 348384 558628 348390 558640
rect 357434 558628 357440 558640
rect 357492 558628 357498 558680
rect 484486 558668 484492 558680
rect 357544 558640 484492 558668
rect 75730 558560 75736 558612
rect 75788 558600 75794 558612
rect 84286 558600 84292 558612
rect 75788 558572 84292 558600
rect 75788 558560 75794 558572
rect 84286 558560 84292 558572
rect 84344 558600 84350 558612
rect 93578 558600 93584 558612
rect 84344 558572 93584 558600
rect 84344 558560 84350 558572
rect 93578 558560 93584 558572
rect 93636 558560 93642 558612
rect 108574 558560 108580 558612
rect 108632 558600 108638 558612
rect 211338 558600 211344 558612
rect 108632 558572 211344 558600
rect 108632 558560 108638 558572
rect 211338 558560 211344 558572
rect 211396 558560 211402 558612
rect 212534 558560 212540 558612
rect 212592 558600 212598 558612
rect 213178 558600 213184 558612
rect 212592 558572 213184 558600
rect 212592 558560 212598 558572
rect 213178 558560 213184 558572
rect 213236 558600 213242 558612
rect 222286 558600 222292 558612
rect 213236 558572 222292 558600
rect 213236 558560 213242 558572
rect 222286 558560 222292 558572
rect 222344 558600 222350 558612
rect 231854 558600 231860 558612
rect 222344 558572 231860 558600
rect 222344 558560 222350 558572
rect 231854 558560 231860 558572
rect 231912 558560 231918 558612
rect 336642 558560 336648 558612
rect 336700 558600 336706 558612
rect 346302 558600 346308 558612
rect 336700 558572 346308 558600
rect 336700 558560 336706 558572
rect 346302 558560 346308 558572
rect 346360 558560 346366 558612
rect 346946 558600 346952 558612
rect 346859 558572 346952 558600
rect 346946 558560 346952 558572
rect 347004 558600 347010 558612
rect 356054 558600 356060 558612
rect 347004 558572 356060 558600
rect 347004 558560 347010 558572
rect 356054 558560 356060 558572
rect 356112 558560 356118 558612
rect 356790 558560 356796 558612
rect 356848 558600 356854 558612
rect 357544 558600 357572 558640
rect 484486 558628 484492 558640
rect 484544 558628 484550 558680
rect 356848 558572 357572 558600
rect 356848 558560 356854 558572
rect 453482 558560 453488 558612
rect 453540 558600 453546 558612
rect 462958 558600 462964 558612
rect 453540 558572 462964 558600
rect 453540 558560 453546 558572
rect 462958 558560 462964 558572
rect 463016 558600 463022 558612
rect 463602 558600 463608 558612
rect 463016 558572 463608 558600
rect 463016 558560 463022 558572
rect 463602 558560 463608 558572
rect 463660 558560 463666 558612
rect 464338 558560 464344 558612
rect 464396 558600 464402 558612
rect 473538 558600 473544 558612
rect 464396 558572 473544 558600
rect 464396 558560 464402 558572
rect 473538 558560 473544 558572
rect 473596 558600 473602 558612
rect 483014 558600 483020 558612
rect 473596 558572 483020 558600
rect 473596 558560 473602 558572
rect 483014 558560 483020 558572
rect 483072 558560 483078 558612
rect 72418 558492 72424 558544
rect 72476 558532 72482 558544
rect 81618 558532 81624 558544
rect 72476 558504 81624 558532
rect 72476 558492 72482 558504
rect 81618 558492 81624 558504
rect 81676 558492 81682 558544
rect 86862 558492 86868 558544
rect 86920 558532 86926 558544
rect 95326 558532 95332 558544
rect 86920 558504 95332 558532
rect 86920 558492 86926 558504
rect 95326 558492 95332 558504
rect 95384 558492 95390 558544
rect 96614 558492 96620 558544
rect 96672 558532 96678 558544
rect 106274 558532 106280 558544
rect 96672 558504 106280 558532
rect 96672 558492 96678 558504
rect 106274 558492 106280 558504
rect 106332 558532 106338 558544
rect 107470 558532 107476 558544
rect 106332 558504 107476 558532
rect 106332 558492 106338 558504
rect 107470 558492 107476 558504
rect 107528 558492 107534 558544
rect 107838 558492 107844 558544
rect 107896 558532 107902 558544
rect 209774 558532 209780 558544
rect 107896 558504 209780 558532
rect 107896 558492 107902 558504
rect 209774 558492 209780 558504
rect 209832 558492 209838 558544
rect 211154 558492 211160 558544
rect 211212 558532 211218 558544
rect 211890 558532 211896 558544
rect 211212 558504 211896 558532
rect 211212 558492 211218 558504
rect 211890 558492 211896 558504
rect 211948 558532 211954 558544
rect 221090 558532 221096 558544
rect 211948 558504 221096 558532
rect 211948 558492 211954 558504
rect 221090 558492 221096 558504
rect 221148 558532 221154 558544
rect 230474 558532 230480 558544
rect 221148 558504 230480 558532
rect 221148 558492 221154 558504
rect 230474 558492 230480 558504
rect 230532 558492 230538 558544
rect 337378 558492 337384 558544
rect 337436 558532 337442 558544
rect 346964 558532 346992 558560
rect 337436 558504 346992 558532
rect 337436 558492 337442 558504
rect 460382 558492 460388 558544
rect 460440 558532 460446 558544
rect 460842 558532 460848 558544
rect 460440 558504 460848 558532
rect 460440 558492 460446 558504
rect 460842 558492 460848 558504
rect 460900 558532 460906 558544
rect 470042 558532 470048 558544
rect 460900 558504 470048 558532
rect 460900 558492 460906 558504
rect 470042 558492 470048 558504
rect 470100 558532 470106 558544
rect 479426 558532 479432 558544
rect 470100 558504 479432 558532
rect 470100 558492 470106 558504
rect 479426 558492 479432 558504
rect 479484 558532 479490 558544
rect 488534 558532 488540 558544
rect 479484 558504 488540 558532
rect 479484 558492 479490 558504
rect 488534 558492 488540 558504
rect 488592 558492 488598 558544
rect 76006 558424 76012 558476
rect 76064 558464 76070 558476
rect 85390 558464 85396 558476
rect 76064 558436 85396 558464
rect 76064 558424 76070 558436
rect 85390 558424 85396 558436
rect 85448 558464 85454 558476
rect 94590 558464 94596 558476
rect 85448 558436 94596 558464
rect 85448 558424 85454 558436
rect 94590 558424 94596 558436
rect 94648 558464 94654 558476
rect 103974 558464 103980 558476
rect 94648 558436 103980 558464
rect 94648 558424 94654 558436
rect 103974 558424 103980 558436
rect 104032 558464 104038 558476
rect 104710 558464 104716 558476
rect 104032 558436 104716 558464
rect 104032 558424 104038 558436
rect 104710 558424 104716 558436
rect 104768 558424 104774 558476
rect 166902 558424 166908 558476
rect 166960 558464 166966 558476
rect 201494 558464 201500 558476
rect 166960 558436 201500 558464
rect 166960 558424 166966 558436
rect 201494 558424 201500 558436
rect 201552 558424 201558 558476
rect 331306 558424 331312 558476
rect 331364 558464 331370 558476
rect 331766 558464 331772 558476
rect 331364 558436 331772 558464
rect 331364 558424 331370 558436
rect 331766 558424 331772 558436
rect 331824 558464 331830 558476
rect 340966 558464 340972 558476
rect 331824 558436 340972 558464
rect 331824 558424 331830 558436
rect 340966 558424 340972 558436
rect 341024 558464 341030 558476
rect 350534 558464 350540 558476
rect 341024 558436 350540 558464
rect 341024 558424 341030 558436
rect 350534 558424 350540 558436
rect 350592 558424 350598 558476
rect 453298 558424 453304 558476
rect 453356 558464 453362 558476
rect 461762 558464 461768 558476
rect 453356 558436 461768 558464
rect 453356 558424 453362 558436
rect 461762 558424 461768 558436
rect 461820 558464 461826 558476
rect 471238 558464 471244 558476
rect 461820 558436 471244 558464
rect 461820 558424 461826 558436
rect 471238 558424 471244 558436
rect 471296 558464 471302 558476
rect 480438 558464 480444 558476
rect 471296 558436 480444 558464
rect 471296 558424 471302 558436
rect 480438 558424 480444 558436
rect 480496 558424 480502 558476
rect 73706 558356 73712 558408
rect 73764 558396 73770 558408
rect 82906 558396 82912 558408
rect 73764 558368 82912 558396
rect 73764 558356 73770 558368
rect 82906 558356 82912 558368
rect 82964 558396 82970 558408
rect 92474 558396 92480 558408
rect 82964 558368 92480 558396
rect 82964 558356 82970 558368
rect 92474 558356 92480 558368
rect 92532 558396 92538 558408
rect 100754 558396 100760 558408
rect 92532 558368 100760 558396
rect 92532 558356 92538 558368
rect 100754 558356 100760 558368
rect 100812 558356 100818 558408
rect 165522 558356 165528 558408
rect 165580 558396 165586 558408
rect 200206 558396 200212 558408
rect 165580 558368 200212 558396
rect 165580 558356 165586 558368
rect 200206 558356 200212 558368
rect 200264 558356 200270 558408
rect 218054 558356 218060 558408
rect 218112 558396 218118 558408
rect 218882 558396 218888 558408
rect 218112 558368 218888 558396
rect 218112 558356 218118 558368
rect 218882 558356 218888 558368
rect 218940 558396 218946 558408
rect 227714 558396 227720 558408
rect 218940 558368 227720 558396
rect 218940 558356 218946 558368
rect 227714 558356 227720 558368
rect 227772 558356 227778 558408
rect 227806 558356 227812 558408
rect 227864 558396 227870 558408
rect 229462 558396 229468 558408
rect 227864 558368 229468 558396
rect 227864 558356 227870 558368
rect 229462 558356 229468 558368
rect 229520 558396 229526 558408
rect 238754 558396 238760 558408
rect 229520 558368 238760 558396
rect 229520 558356 229526 558368
rect 238754 558356 238760 558368
rect 238812 558356 238818 558408
rect 332686 558356 332692 558408
rect 332744 558396 332750 558408
rect 342530 558396 342536 558408
rect 332744 558368 342536 558396
rect 332744 558356 332750 558368
rect 342530 558356 342536 558368
rect 342588 558396 342594 558408
rect 347958 558396 347964 558408
rect 342588 558368 347964 558396
rect 342588 558356 342594 558368
rect 347958 558356 347964 558368
rect 348016 558356 348022 558408
rect 358170 558356 358176 558408
rect 358228 558396 358234 558408
rect 455414 558396 455420 558408
rect 358228 558368 455420 558396
rect 358228 558356 358234 558368
rect 455414 558356 455420 558368
rect 455472 558356 455478 558408
rect 463602 558356 463608 558408
rect 463660 558396 463666 558408
rect 472250 558396 472256 558408
rect 463660 558368 472256 558396
rect 463660 558356 463666 558368
rect 472250 558356 472256 558368
rect 472308 558396 472314 558408
rect 481634 558396 481640 558408
rect 472308 558368 481640 558396
rect 472308 558356 472314 558368
rect 481634 558356 481640 558368
rect 481692 558356 481698 558408
rect 75822 558288 75828 558340
rect 75880 558328 75886 558340
rect 80054 558328 80060 558340
rect 75880 558300 80060 558328
rect 75880 558288 75886 558300
rect 80054 558288 80060 558300
rect 80112 558288 80118 558340
rect 88978 558288 88984 558340
rect 89036 558328 89042 558340
rect 98270 558328 98276 558340
rect 89036 558300 98276 558328
rect 89036 558288 89042 558300
rect 98270 558288 98276 558300
rect 98328 558328 98334 558340
rect 107838 558328 107844 558340
rect 98328 558300 107844 558328
rect 98328 558288 98334 558300
rect 107838 558288 107844 558300
rect 107896 558288 107902 558340
rect 162762 558288 162768 558340
rect 162820 558328 162826 558340
rect 198734 558328 198740 558340
rect 162820 558300 198740 558328
rect 162820 558288 162826 558300
rect 198734 558288 198740 558300
rect 198792 558288 198798 558340
rect 213914 558288 213920 558340
rect 213972 558328 213978 558340
rect 223574 558328 223580 558340
rect 213972 558300 223580 558328
rect 213972 558288 213978 558300
rect 223574 558288 223580 558300
rect 223632 558288 223638 558340
rect 225782 558288 225788 558340
rect 225840 558328 225846 558340
rect 234614 558328 234620 558340
rect 225840 558300 234620 558328
rect 225840 558288 225846 558300
rect 234614 558288 234620 558300
rect 234672 558288 234678 558340
rect 339862 558288 339868 558340
rect 339920 558328 339926 558340
rect 349522 558328 349528 558340
rect 339920 558300 349528 558328
rect 339920 558288 339926 558300
rect 349522 558288 349528 558300
rect 349580 558328 349586 558340
rect 357710 558328 357716 558340
rect 349580 558300 357716 558328
rect 349580 558288 349586 558300
rect 357710 558288 357716 558300
rect 357768 558288 357774 558340
rect 359458 558288 359464 558340
rect 359516 558328 359522 558340
rect 456794 558328 456800 558340
rect 359516 558300 456800 558328
rect 359516 558288 359522 558300
rect 456794 558288 456800 558300
rect 456852 558288 456858 558340
rect 465166 558288 465172 558340
rect 465224 558328 465230 558340
rect 474826 558328 474832 558340
rect 465224 558300 474832 558328
rect 465224 558288 465230 558300
rect 474826 558288 474832 558300
rect 474884 558288 474890 558340
rect 477586 558288 477592 558340
rect 477644 558328 477650 558340
rect 478322 558328 478328 558340
rect 477644 558300 478328 558328
rect 477644 558288 477650 558300
rect 478322 558288 478328 558300
rect 478380 558328 478386 558340
rect 487154 558328 487160 558340
rect 478380 558300 487160 558328
rect 478380 558288 478386 558300
rect 487154 558288 487160 558300
rect 487212 558288 487218 558340
rect 78490 558220 78496 558272
rect 78548 558260 78554 558272
rect 87874 558260 87880 558272
rect 78548 558232 87880 558260
rect 78548 558220 78554 558232
rect 87874 558220 87880 558232
rect 87932 558220 87938 558272
rect 91002 558220 91008 558272
rect 91060 558260 91066 558272
rect 99558 558260 99564 558272
rect 91060 558232 99564 558260
rect 91060 558220 91066 558232
rect 99558 558220 99564 558232
rect 99616 558260 99622 558272
rect 108574 558260 108580 558272
rect 99616 558232 108580 558260
rect 99616 558220 99622 558232
rect 108574 558220 108580 558232
rect 108632 558220 108638 558272
rect 161382 558220 161388 558272
rect 161440 558260 161446 558272
rect 197354 558260 197360 558272
rect 161440 558232 197360 558260
rect 161440 558220 161446 558232
rect 197354 558220 197360 558232
rect 197412 558220 197418 558272
rect 216674 558220 216680 558272
rect 216732 558260 216738 558272
rect 217594 558260 217600 558272
rect 216732 558232 217600 558260
rect 216732 558220 216738 558232
rect 217594 558220 217600 558232
rect 217652 558260 217658 558272
rect 226334 558260 226340 558272
rect 217652 558232 226340 558260
rect 217652 558220 217658 558232
rect 226334 558220 226340 558232
rect 226392 558220 226398 558272
rect 227714 558220 227720 558272
rect 227772 558260 227778 558272
rect 237374 558260 237380 558272
rect 227772 558232 237380 558260
rect 227772 558220 227778 558232
rect 237374 558220 237380 558232
rect 237432 558220 237438 558272
rect 291838 558220 291844 558272
rect 291896 558260 291902 558272
rect 329834 558260 329840 558272
rect 291896 558232 329840 558260
rect 291896 558220 291902 558232
rect 329834 558220 329840 558232
rect 329892 558220 329898 558272
rect 334066 558220 334072 558272
rect 334124 558260 334130 558272
rect 343726 558260 343732 558272
rect 334124 558232 343732 558260
rect 334124 558220 334130 558232
rect 343726 558220 343732 558232
rect 343784 558220 343790 558272
rect 346302 558220 346308 558272
rect 346360 558260 346366 558272
rect 354674 558260 354680 558272
rect 346360 558232 354680 558260
rect 346360 558220 346366 558232
rect 354674 558220 354680 558232
rect 354732 558220 354738 558272
rect 359550 558220 359556 558272
rect 359608 558260 359614 558272
rect 458174 558260 458180 558272
rect 359608 558232 458180 558260
rect 359608 558220 359614 558232
rect 458174 558220 458180 558232
rect 458232 558220 458238 558272
rect 467098 558220 467104 558272
rect 467156 558260 467162 558272
rect 488534 558260 488540 558272
rect 467156 558232 488540 558260
rect 467156 558220 467162 558232
rect 488534 558220 488540 558232
rect 488592 558220 488598 558272
rect 64322 558152 64328 558204
rect 64380 558192 64386 558204
rect 193766 558192 193772 558204
rect 64380 558164 193772 558192
rect 64380 558152 64386 558164
rect 193766 558152 193772 558164
rect 193824 558192 193830 558204
rect 313734 558192 313740 558204
rect 193824 558164 313740 558192
rect 193824 558152 193830 558164
rect 313734 558152 313740 558164
rect 313792 558192 313798 558204
rect 443086 558192 443092 558204
rect 313792 558164 443092 558192
rect 313792 558152 313798 558164
rect 443086 558152 443092 558164
rect 443144 558152 443150 558204
rect 443638 558152 443644 558204
rect 443696 558192 443702 558204
rect 459554 558192 459560 558204
rect 443696 558164 459560 558192
rect 443696 558152 443702 558164
rect 459554 558152 459560 558164
rect 459612 558152 459618 558204
rect 465718 558152 465724 558204
rect 465776 558192 465782 558204
rect 487154 558192 487160 558204
rect 465776 558164 487160 558192
rect 465776 558152 465782 558164
rect 487154 558152 487160 558164
rect 487212 558152 487218 558204
rect 128262 558084 128268 558136
rect 128320 558124 128326 558136
rect 195974 558124 195980 558136
rect 128320 558096 195980 558124
rect 128320 558084 128326 558096
rect 195974 558084 195980 558096
rect 196032 558084 196038 558136
rect 204898 558084 204904 558136
rect 204956 558124 204962 558136
rect 213914 558124 213920 558136
rect 204956 558096 213920 558124
rect 204956 558084 204962 558096
rect 213914 558084 213920 558096
rect 213972 558084 213978 558136
rect 290458 558084 290464 558136
rect 290516 558124 290522 558136
rect 331214 558124 331220 558136
rect 290516 558096 331220 558124
rect 290516 558084 290522 558096
rect 331214 558084 331220 558096
rect 331272 558084 331278 558136
rect 349798 558084 349804 558136
rect 349856 558124 349862 558136
rect 452654 558124 452660 558136
rect 349856 558096 452660 558124
rect 349856 558084 349862 558096
rect 452654 558084 452660 558096
rect 452712 558084 452718 558136
rect 454678 558084 454684 558136
rect 454736 558124 454742 558136
rect 464246 558124 464252 558136
rect 454736 558096 464252 558124
rect 454736 558084 454742 558096
rect 464246 558084 464252 558096
rect 464304 558084 464310 558136
rect 464338 558084 464344 558136
rect 464396 558124 464402 558136
rect 485774 558124 485780 558136
rect 464396 558096 485780 558124
rect 464396 558084 464402 558096
rect 485774 558084 485780 558096
rect 485832 558084 485838 558136
rect 80698 558016 80704 558068
rect 80756 558056 80762 558068
rect 82814 558056 82820 558068
rect 80756 558028 82820 558056
rect 80756 558016 80762 558028
rect 82814 558016 82820 558028
rect 82872 558016 82878 558068
rect 100754 558016 100760 558068
rect 100812 558056 100818 558068
rect 101858 558056 101864 558068
rect 100812 558028 101864 558056
rect 100812 558016 100818 558028
rect 101858 558016 101864 558028
rect 101916 558056 101922 558068
rect 198734 558056 198740 558068
rect 101916 558028 198740 558056
rect 101916 558016 101922 558028
rect 198734 558016 198740 558028
rect 198792 558016 198798 558068
rect 206278 558016 206284 558068
rect 206336 558056 206342 558068
rect 215294 558056 215300 558068
rect 206336 558028 215300 558056
rect 206336 558016 206342 558028
rect 215294 558016 215300 558028
rect 215352 558016 215358 558068
rect 322198 558016 322204 558068
rect 322256 558056 322262 558068
rect 328454 558056 328460 558068
rect 322256 558028 328460 558056
rect 322256 558016 322262 558028
rect 328454 558016 328460 558028
rect 328512 558016 328518 558068
rect 329098 558016 329104 558068
rect 329156 558056 329162 558068
rect 337378 558056 337384 558068
rect 329156 558028 337384 558056
rect 329156 558016 329162 558028
rect 337378 558016 337384 558028
rect 337436 558016 337442 558068
rect 352558 558016 352564 558068
rect 352616 558056 352622 558068
rect 476114 558056 476120 558068
rect 352616 558028 476120 558056
rect 352616 558016 352622 558028
rect 476114 558016 476120 558028
rect 476172 558016 476178 558068
rect 100294 557948 100300 558000
rect 100352 557988 100358 558000
rect 197354 557988 197360 558000
rect 100352 557960 197360 557988
rect 100352 557948 100358 557960
rect 197354 557948 197360 557960
rect 197412 557948 197418 558000
rect 209222 557948 209228 558000
rect 209280 557988 209286 558000
rect 216674 557988 216680 558000
rect 209280 557960 216680 557988
rect 209280 557948 209286 557960
rect 216674 557948 216680 557960
rect 216732 557948 216738 558000
rect 327718 557948 327724 558000
rect 327776 557988 327782 558000
rect 336642 557988 336648 558000
rect 327776 557960 336648 557988
rect 327776 557948 327782 557960
rect 336642 557948 336648 557960
rect 336700 557948 336706 558000
rect 352650 557948 352656 558000
rect 352708 557988 352714 558000
rect 477494 557988 477500 558000
rect 352708 557960 477500 557988
rect 352708 557948 352714 557960
rect 477494 557948 477500 557960
rect 477552 557948 477558 558000
rect 71682 557880 71688 557932
rect 71740 557920 71746 557932
rect 78674 557920 78680 557932
rect 71740 557892 78680 557920
rect 71740 557880 71746 557892
rect 78674 557880 78680 557892
rect 78732 557880 78738 557932
rect 202138 557880 202144 557932
rect 202196 557920 202202 557932
rect 211154 557920 211160 557932
rect 202196 557892 211160 557920
rect 202196 557880 202202 557892
rect 211154 557880 211160 557892
rect 211212 557880 211218 557932
rect 322290 557880 322296 557932
rect 322348 557920 322354 557932
rect 331306 557920 331312 557932
rect 322348 557892 331312 557920
rect 322348 557880 322354 557892
rect 331306 557880 331312 557892
rect 331364 557880 331370 557932
rect 352742 557880 352748 557932
rect 352800 557920 352806 557932
rect 478874 557920 478880 557932
rect 352800 557892 478880 557920
rect 352800 557880 352806 557892
rect 478874 557880 478880 557892
rect 478932 557880 478938 557932
rect 70302 557812 70308 557864
rect 70360 557852 70366 557864
rect 77294 557852 77300 557864
rect 70360 557824 77300 557852
rect 70360 557812 70366 557824
rect 77294 557812 77300 557824
rect 77352 557812 77358 557864
rect 93578 557812 93584 557864
rect 93636 557852 93642 557864
rect 102686 557852 102692 557864
rect 93636 557824 102692 557852
rect 93636 557812 93642 557824
rect 102686 557812 102692 557824
rect 102744 557852 102750 557864
rect 201494 557852 201500 557864
rect 102744 557824 201500 557852
rect 102744 557812 102750 557824
rect 201494 557812 201500 557824
rect 201552 557812 201558 557864
rect 203518 557812 203524 557864
rect 203576 557852 203582 557864
rect 212534 557852 212540 557864
rect 203576 557824 212540 557852
rect 203576 557812 203582 557824
rect 212534 557812 212540 557824
rect 212592 557812 212598 557864
rect 302878 557812 302884 557864
rect 302936 557852 302942 557864
rect 322934 557852 322940 557864
rect 302936 557824 322940 557852
rect 302936 557812 302942 557824
rect 322934 557812 322940 557824
rect 322992 557812 322998 557864
rect 323670 557812 323676 557864
rect 323728 557852 323734 557864
rect 332686 557852 332692 557864
rect 323728 557824 332692 557852
rect 323728 557812 323734 557824
rect 332686 557812 332692 557824
rect 332744 557812 332750 557864
rect 353938 557812 353944 557864
rect 353996 557852 354002 557864
rect 480530 557852 480536 557864
rect 353996 557824 480536 557852
rect 353996 557812 354002 557824
rect 480530 557812 480536 557824
rect 480588 557812 480594 557864
rect 66162 557744 66168 557796
rect 66220 557784 66226 557796
rect 74534 557784 74540 557796
rect 66220 557756 74540 557784
rect 66220 557744 66226 557756
rect 74534 557744 74540 557756
rect 74592 557744 74598 557796
rect 106090 557744 106096 557796
rect 106148 557784 106154 557796
rect 205634 557784 205640 557796
rect 106148 557756 205640 557784
rect 106148 557744 106154 557756
rect 205634 557744 205640 557756
rect 205692 557744 205698 557796
rect 287790 557744 287796 557796
rect 287848 557784 287854 557796
rect 317414 557784 317420 557796
rect 287848 557756 317420 557784
rect 287848 557744 287854 557756
rect 317414 557744 317420 557756
rect 317472 557744 317478 557796
rect 324958 557744 324964 557796
rect 325016 557784 325022 557796
rect 334066 557784 334072 557796
rect 325016 557756 334072 557784
rect 325016 557744 325022 557756
rect 334066 557744 334072 557756
rect 334124 557744 334130 557796
rect 356698 557744 356704 557796
rect 356756 557784 356762 557796
rect 483014 557784 483020 557796
rect 356756 557756 483020 557784
rect 356756 557744 356762 557756
rect 483014 557744 483020 557756
rect 483072 557744 483078 557796
rect 67450 557676 67456 557728
rect 67508 557716 67514 557728
rect 75914 557716 75920 557728
rect 67508 557688 75920 557716
rect 67508 557676 67514 557688
rect 75914 557676 75920 557688
rect 75972 557676 75978 557728
rect 107470 557676 107476 557728
rect 107528 557716 107534 557728
rect 207014 557716 207020 557728
rect 107528 557688 207020 557716
rect 107528 557676 107534 557688
rect 207014 557676 207020 557688
rect 207072 557676 207078 557728
rect 207658 557676 207664 557728
rect 207716 557716 207722 557728
rect 216766 557716 216772 557728
rect 207716 557688 216772 557716
rect 207716 557676 207722 557688
rect 216766 557676 216772 557688
rect 216824 557676 216830 557728
rect 286410 557676 286416 557728
rect 286468 557716 286474 557728
rect 320174 557716 320180 557728
rect 286468 557688 320180 557716
rect 286468 557676 286474 557688
rect 320174 557676 320180 557688
rect 320232 557676 320238 557728
rect 326338 557676 326344 557728
rect 326396 557716 326402 557728
rect 335446 557716 335452 557728
rect 326396 557688 335452 557716
rect 326396 557676 326402 557688
rect 335446 557676 335452 557688
rect 335504 557676 335510 557728
rect 354030 557676 354036 557728
rect 354088 557716 354094 557728
rect 481634 557716 481640 557728
rect 354088 557688 481640 557716
rect 354088 557676 354094 557688
rect 481634 557676 481640 557688
rect 481692 557676 481698 557728
rect 63402 557608 63408 557660
rect 63460 557648 63466 557660
rect 73154 557648 73160 557660
rect 63460 557620 73160 557648
rect 63460 557608 63466 557620
rect 73154 557608 73160 557620
rect 73212 557608 73218 557660
rect 104710 557608 104716 557660
rect 104768 557648 104774 557660
rect 202874 557648 202880 557660
rect 104768 557620 202880 557648
rect 104768 557608 104774 557620
rect 202874 557608 202880 557620
rect 202932 557608 202938 557660
rect 209038 557608 209044 557660
rect 209096 557648 209102 557660
rect 218054 557648 218060 557660
rect 209096 557620 218060 557648
rect 209096 557608 209102 557620
rect 218054 557608 218060 557620
rect 218112 557608 218118 557660
rect 329282 557608 329288 557660
rect 329340 557648 329346 557660
rect 338942 557648 338948 557660
rect 329340 557620 338948 557648
rect 329340 557608 329346 557620
rect 338942 557608 338948 557620
rect 339000 557608 339006 557660
rect 358078 557608 358084 557660
rect 358136 557648 358142 557660
rect 454034 557648 454040 557660
rect 358136 557620 454040 557648
rect 358136 557608 358142 557620
rect 454034 557608 454040 557620
rect 454092 557608 454098 557660
rect 456058 557608 456064 557660
rect 456116 557648 456122 557660
rect 465166 557648 465172 557660
rect 456116 557620 465172 557648
rect 456116 557608 456122 557620
rect 465166 557608 465172 557620
rect 465224 557608 465230 557660
rect 468570 557608 468576 557660
rect 468628 557648 468634 557660
rect 477586 557648 477592 557660
rect 468628 557620 477592 557648
rect 468628 557608 468634 557620
rect 477586 557608 477592 557620
rect 477644 557608 477650 557660
rect 62022 557540 62028 557592
rect 62080 557580 62086 557592
rect 71774 557580 71780 557592
rect 62080 557552 71780 557580
rect 62080 557540 62086 557552
rect 71774 557540 71780 557552
rect 71832 557540 71838 557592
rect 74442 557540 74448 557592
rect 74500 557580 74506 557592
rect 78674 557580 78680 557592
rect 74500 557552 78680 557580
rect 74500 557540 74506 557552
rect 78674 557540 78680 557552
rect 78732 557540 78738 557592
rect 210418 557540 210424 557592
rect 210476 557580 210482 557592
rect 220078 557580 220084 557592
rect 210476 557552 220084 557580
rect 210476 557540 210482 557552
rect 220078 557540 220084 557552
rect 220136 557580 220142 557592
rect 227806 557580 227812 557592
rect 220136 557552 227812 557580
rect 220136 557540 220142 557552
rect 227806 557540 227812 557552
rect 227864 557540 227870 557592
rect 330478 557540 330484 557592
rect 330536 557580 330542 557592
rect 339862 557580 339868 557592
rect 330536 557552 339868 557580
rect 330536 557540 330542 557552
rect 339862 557540 339868 557552
rect 339920 557540 339926 557592
rect 450538 557540 450544 557592
rect 450596 557580 450602 557592
rect 451366 557580 451372 557592
rect 450596 557552 451372 557580
rect 450596 557540 450602 557552
rect 451366 557540 451372 557552
rect 451424 557540 451430 557592
rect 457438 557540 457444 557592
rect 457496 557580 457502 557592
rect 466546 557580 466552 557592
rect 457496 557552 466552 557580
rect 457496 557540 457502 557552
rect 466546 557540 466552 557552
rect 466604 557580 466610 557592
rect 474642 557580 474648 557592
rect 466604 557552 474648 557580
rect 466604 557540 466610 557552
rect 474642 557540 474648 557552
rect 474700 557540 474706 557592
rect 474826 557540 474832 557592
rect 474884 557580 474890 557592
rect 483014 557580 483020 557592
rect 474884 557552 483020 557580
rect 474884 557540 474890 557552
rect 483014 557540 483020 557552
rect 483072 557540 483078 557592
rect 58250 556180 58256 556232
rect 58308 556220 58314 556232
rect 579614 556220 579620 556232
rect 58308 556192 579620 556220
rect 58308 556180 58314 556192
rect 579614 556180 579620 556192
rect 579672 556180 579678 556232
rect 169846 553392 169852 553444
rect 169904 553432 169910 553444
rect 170030 553432 170036 553444
rect 169904 553404 170036 553432
rect 169904 553392 169910 553404
rect 170030 553392 170036 553404
rect 170088 553392 170094 553444
rect 57330 545096 57336 545148
rect 57388 545136 57394 545148
rect 580166 545136 580172 545148
rect 57388 545108 580172 545136
rect 57388 545096 57394 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 56778 543668 56784 543720
rect 56836 543708 56842 543720
rect 146018 543708 146024 543720
rect 56836 543680 146024 543708
rect 56836 543668 56842 543680
rect 146018 543668 146024 543680
rect 146076 543668 146082 543720
rect 206922 543668 206928 543720
rect 206980 543708 206986 543720
rect 220722 543708 220728 543720
rect 206980 543680 220728 543708
rect 206980 543668 206986 543680
rect 220722 543668 220728 543680
rect 220780 543668 220786 543720
rect 229002 543668 229008 543720
rect 229060 543708 229066 543720
rect 260190 543708 260196 543720
rect 229060 543680 260196 543708
rect 229060 543668 229066 543680
rect 260190 543668 260196 543680
rect 260248 543668 260254 543720
rect 56870 543600 56876 543652
rect 56928 543640 56934 543652
rect 148134 543640 148140 543652
rect 56928 543612 148140 543640
rect 56928 543600 56934 543612
rect 148134 543600 148140 543612
rect 148192 543600 148198 543652
rect 205542 543600 205548 543652
rect 205600 543640 205606 543652
rect 218698 543640 218704 543652
rect 205600 543612 218704 543640
rect 205600 543600 205606 543612
rect 218698 543600 218704 543612
rect 218756 543600 218762 543652
rect 227622 543600 227628 543652
rect 227680 543640 227686 543652
rect 258074 543640 258080 543652
rect 227680 543612 258080 543640
rect 227680 543600 227686 543612
rect 258074 543600 258080 543612
rect 258132 543600 258138 543652
rect 61010 543532 61016 543584
rect 61068 543572 61074 543584
rect 62022 543572 62028 543584
rect 61068 543544 62028 543572
rect 61068 543532 61074 543544
rect 62022 543532 62028 543544
rect 62080 543532 62086 543584
rect 150158 543572 150164 543584
rect 62132 543544 150164 543572
rect 56962 543464 56968 543516
rect 57020 543504 57026 543516
rect 62132 543504 62160 543544
rect 150158 543532 150164 543544
rect 150216 543532 150222 543584
rect 164694 543532 164700 543584
rect 164752 543572 164758 543584
rect 165522 543572 165528 543584
rect 164752 543544 165528 543572
rect 164752 543532 164758 543544
rect 165522 543532 165528 543544
rect 165580 543532 165586 543584
rect 177206 543532 177212 543584
rect 177264 543572 177270 543584
rect 177942 543572 177948 543584
rect 177264 543544 177948 543572
rect 177264 543532 177270 543544
rect 177942 543532 177948 543544
rect 178000 543532 178006 543584
rect 208302 543532 208308 543584
rect 208360 543572 208366 543584
rect 222838 543572 222844 543584
rect 208360 543544 222844 543572
rect 208360 543532 208366 543544
rect 222838 543532 222844 543544
rect 222896 543532 222902 543584
rect 231762 543532 231768 543584
rect 231820 543572 231826 543584
rect 264330 543572 264336 543584
rect 231820 543544 264336 543572
rect 231820 543532 231826 543544
rect 264330 543532 264336 543544
rect 264388 543532 264394 543584
rect 152274 543504 152280 543516
rect 57020 543476 62160 543504
rect 62224 543476 152280 543504
rect 57020 543464 57026 543476
rect 57054 543396 57060 543448
rect 57112 543436 57118 543448
rect 62224 543436 62252 543476
rect 152274 543464 152280 543476
rect 152332 543464 152338 543516
rect 160554 543464 160560 543516
rect 160612 543504 160618 543516
rect 161382 543504 161388 543516
rect 160612 543476 161388 543504
rect 160612 543464 160618 543476
rect 161382 543464 161388 543476
rect 161440 543464 161446 543516
rect 193766 543464 193772 543516
rect 193824 543504 193830 543516
rect 209038 543504 209044 543516
rect 193824 543476 209044 543504
rect 193824 543464 193830 543476
rect 209038 543464 209044 543476
rect 209096 543464 209102 543516
rect 209682 543464 209688 543516
rect 209740 543504 209746 543516
rect 224862 543504 224868 543516
rect 209740 543476 224868 543504
rect 209740 543464 209746 543476
rect 224862 543464 224868 543476
rect 224920 543464 224926 543516
rect 230382 543464 230388 543516
rect 230440 543504 230446 543516
rect 262214 543504 262220 543516
rect 230440 543476 262220 543504
rect 230440 543464 230446 543476
rect 262214 543464 262220 543476
rect 262272 543464 262278 543516
rect 154390 543436 154396 543448
rect 57112 543408 62252 543436
rect 62316 543408 154396 543436
rect 57112 543396 57118 543408
rect 57146 543328 57152 543380
rect 57204 543368 57210 543380
rect 62316 543368 62344 543408
rect 154390 543396 154396 543408
rect 154448 543396 154454 543448
rect 195882 543396 195888 543448
rect 195940 543436 195946 543448
rect 210418 543436 210424 543448
rect 195940 543408 210424 543436
rect 195940 543396 195946 543408
rect 210418 543396 210424 543408
rect 210476 543396 210482 543448
rect 210970 543396 210976 543448
rect 211028 543436 211034 543448
rect 226978 543436 226984 543448
rect 211028 543408 226984 543436
rect 211028 543396 211034 543408
rect 226978 543396 226984 543408
rect 227036 543396 227042 543448
rect 233050 543396 233056 543448
rect 233108 543436 233114 543448
rect 266446 543436 266452 543448
rect 233108 543408 266452 543436
rect 233108 543396 233114 543408
rect 266446 543396 266452 543408
rect 266504 543396 266510 543448
rect 156414 543368 156420 543380
rect 57204 543340 62344 543368
rect 62408 543340 156420 543368
rect 57204 543328 57210 543340
rect 57238 543260 57244 543312
rect 57296 543300 57302 543312
rect 62408 543300 62436 543340
rect 156414 543328 156420 543340
rect 156472 543328 156478 543380
rect 189626 543328 189632 543380
rect 189684 543368 189690 543380
rect 207658 543368 207664 543380
rect 189684 543340 207664 543368
rect 189684 543328 189690 543340
rect 207658 543328 207664 543340
rect 207716 543328 207722 543380
rect 212442 543328 212448 543380
rect 212500 543368 212506 543380
rect 231118 543368 231124 543380
rect 212500 543340 231124 543368
rect 212500 543328 212506 543340
rect 231118 543328 231124 543340
rect 231176 543328 231182 543380
rect 233142 543328 233148 543380
rect 233200 543368 233206 543380
rect 268470 543368 268476 543380
rect 233200 543340 268476 543368
rect 233200 543328 233206 543340
rect 268470 543328 268476 543340
rect 268528 543328 268534 543380
rect 57296 543272 62436 543300
rect 57296 543260 57302 543272
rect 65150 543260 65156 543312
rect 65208 543300 65214 543312
rect 66162 543300 66168 543312
rect 65208 543272 66168 543300
rect 65208 543260 65214 543272
rect 66162 543260 66168 543272
rect 66220 543260 66226 543312
rect 73430 543260 73436 543312
rect 73488 543300 73494 543312
rect 74442 543300 74448 543312
rect 73488 543272 74448 543300
rect 73488 543260 73494 543272
rect 74442 543260 74448 543272
rect 74500 543260 74506 543312
rect 77570 543260 77576 543312
rect 77628 543300 77634 543312
rect 79318 543300 79324 543312
rect 77628 543272 79324 543300
rect 77628 543260 77634 543272
rect 79318 543260 79324 543272
rect 79376 543260 79382 543312
rect 79686 543260 79692 543312
rect 79744 543300 79750 543312
rect 80698 543300 80704 543312
rect 79744 543272 80704 543300
rect 79744 543260 79750 543272
rect 80698 543260 80704 543272
rect 80756 543260 80762 543312
rect 80790 543260 80796 543312
rect 80848 543300 80854 543312
rect 168834 543300 168840 543312
rect 80848 543272 168840 543300
rect 80848 543260 80854 543272
rect 168834 543260 168840 543272
rect 168892 543260 168898 543312
rect 191742 543260 191748 543312
rect 191800 543300 191806 543312
rect 209222 543300 209228 543312
rect 191800 543272 209228 543300
rect 191800 543260 191806 543272
rect 209222 543260 209228 543272
rect 209280 543260 209286 543312
rect 211062 543260 211068 543312
rect 211120 543300 211126 543312
rect 229094 543300 229100 543312
rect 211120 543272 229100 543300
rect 211120 543260 211126 543272
rect 229094 543260 229100 543272
rect 229152 543260 229158 543312
rect 234522 543260 234528 543312
rect 234580 543300 234586 543312
rect 270586 543300 270592 543312
rect 234580 543272 270592 543300
rect 234580 543260 234586 543272
rect 270586 543260 270592 543272
rect 270644 543260 270650 543312
rect 70118 543192 70124 543244
rect 70176 543232 70182 543244
rect 170950 543232 170956 543244
rect 70176 543204 170956 543232
rect 70176 543192 70182 543204
rect 170950 543192 170956 543204
rect 171008 543192 171014 543244
rect 187510 543192 187516 543244
rect 187568 543232 187574 543244
rect 206278 543232 206284 543244
rect 187568 543204 206284 543232
rect 187568 543192 187574 543204
rect 206278 543192 206284 543204
rect 206336 543192 206342 543244
rect 213822 543192 213828 543244
rect 213880 543232 213886 543244
rect 233234 543232 233240 543244
rect 213880 543204 233240 543232
rect 213880 543192 213886 543204
rect 233234 543192 233240 543204
rect 233292 543192 233298 543244
rect 235902 543192 235908 543244
rect 235960 543232 235966 543244
rect 272610 543232 272616 543244
rect 235960 543204 272616 543232
rect 235960 543192 235966 543204
rect 272610 543192 272616 543204
rect 272668 543192 272674 543244
rect 70210 543124 70216 543176
rect 70268 543164 70274 543176
rect 173066 543164 173072 543176
rect 70268 543136 173072 543164
rect 70268 543124 70274 543136
rect 173066 543124 173072 543136
rect 173124 543124 173130 543176
rect 185486 543124 185492 543176
rect 185544 543164 185550 543176
rect 204898 543164 204904 543176
rect 185544 543136 204904 543164
rect 185544 543124 185550 543136
rect 204898 543124 204904 543136
rect 204956 543124 204962 543176
rect 216582 543124 216588 543176
rect 216640 543164 216646 543176
rect 237374 543164 237380 543176
rect 216640 543136 237380 543164
rect 216640 543124 216646 543136
rect 237374 543124 237380 543136
rect 237432 543124 237438 543176
rect 238662 543124 238668 543176
rect 238720 543164 238726 543176
rect 276750 543164 276756 543176
rect 238720 543136 276756 543164
rect 238720 543124 238726 543136
rect 276750 543124 276756 543136
rect 276808 543124 276814 543176
rect 71590 543056 71596 543108
rect 71648 543096 71654 543108
rect 175090 543096 175096 543108
rect 71648 543068 175096 543096
rect 71648 543056 71654 543068
rect 175090 543056 175096 543068
rect 175148 543056 175154 543108
rect 183370 543056 183376 543108
rect 183428 543096 183434 543108
rect 203518 543096 203524 543108
rect 183428 543068 203524 543096
rect 183428 543056 183434 543068
rect 203518 543056 203524 543068
rect 203576 543056 203582 543108
rect 215202 543056 215208 543108
rect 215260 543096 215266 543108
rect 235258 543096 235264 543108
rect 215260 543068 235264 543096
rect 215260 543056 215266 543068
rect 235258 543056 235264 543068
rect 235316 543056 235322 543108
rect 237282 543056 237288 543108
rect 237340 543096 237346 543108
rect 274726 543096 274732 543108
rect 237340 543068 274732 543096
rect 237340 543056 237346 543068
rect 274726 543056 274732 543068
rect 274784 543056 274790 543108
rect 56686 542988 56692 543040
rect 56744 543028 56750 543040
rect 179230 543028 179236 543040
rect 56744 543000 179236 543028
rect 56744 542988 56750 543000
rect 179230 542988 179236 543000
rect 179288 542988 179294 543040
rect 181346 542988 181352 543040
rect 181404 543028 181410 543040
rect 202138 543028 202144 543040
rect 181404 543000 202144 543028
rect 181404 542988 181410 543000
rect 202138 542988 202144 543000
rect 202196 542988 202202 543040
rect 202782 542988 202788 543040
rect 202840 543028 202846 543040
rect 214558 543028 214564 543040
rect 202840 543000 214564 543028
rect 202840 542988 202846 543000
rect 214558 542988 214564 543000
rect 214616 542988 214622 543040
rect 217962 542988 217968 543040
rect 218020 543028 218026 543040
rect 239398 543028 239404 543040
rect 218020 543000 239404 543028
rect 218020 542988 218026 543000
rect 239398 542988 239404 543000
rect 239456 542988 239462 543040
rect 240042 542988 240048 543040
rect 240100 543028 240106 543040
rect 278866 543028 278872 543040
rect 240100 543000 278872 543028
rect 240100 542988 240106 543000
rect 278866 542988 278872 543000
rect 278924 542988 278930 543040
rect 67542 542920 67548 542972
rect 67600 542960 67606 542972
rect 143994 542960 144000 542972
rect 67600 542932 144000 542960
rect 67600 542920 67606 542932
rect 143994 542920 144000 542932
rect 144052 542920 144058 542972
rect 204162 542920 204168 542972
rect 204220 542960 204226 542972
rect 216582 542960 216588 542972
rect 204220 542932 216588 542960
rect 204220 542920 204226 542932
rect 216582 542920 216588 542932
rect 216640 542920 216646 542972
rect 226242 542920 226248 542972
rect 226300 542960 226306 542972
rect 256050 542960 256056 542972
rect 226300 542932 256056 542960
rect 226300 542920 226306 542932
rect 256050 542920 256056 542932
rect 256108 542920 256114 542972
rect 68922 542852 68928 542904
rect 68980 542892 68986 542904
rect 80790 542892 80796 542904
rect 68980 542864 80796 542892
rect 68980 542852 68986 542864
rect 80790 542852 80796 542864
rect 80848 542852 80854 542904
rect 91002 542852 91008 542904
rect 91060 542892 91066 542904
rect 92106 542892 92112 542904
rect 91060 542864 92112 542892
rect 91060 542852 91066 542864
rect 92106 542852 92112 542864
rect 92164 542852 92170 542904
rect 92382 542852 92388 542904
rect 92440 542892 92446 542904
rect 94130 542892 94136 542904
rect 92440 542864 94136 542892
rect 92440 542852 92446 542864
rect 94130 542852 94136 542864
rect 94188 542852 94194 542904
rect 100662 542852 100668 542904
rect 100720 542892 100726 542904
rect 108666 542892 108672 542904
rect 100720 542864 108672 542892
rect 100720 542852 100726 542864
rect 108666 542852 108672 542864
rect 108724 542852 108730 542904
rect 108942 542852 108948 542904
rect 109000 542892 109006 542904
rect 123202 542892 123208 542904
rect 109000 542864 123208 542892
rect 109000 542852 109006 542864
rect 123202 542852 123208 542864
rect 123260 542852 123266 542904
rect 127342 542852 127348 542904
rect 127400 542892 127406 542904
rect 128262 542892 128268 542904
rect 127400 542864 128268 542892
rect 127400 542852 127406 542864
rect 128262 542852 128268 542864
rect 128320 542852 128326 542904
rect 129458 542852 129464 542904
rect 129516 542892 129522 542904
rect 188430 542892 188436 542904
rect 129516 542864 188436 542892
rect 129516 542852 129522 542864
rect 188430 542852 188436 542864
rect 188488 542852 188494 542904
rect 226150 542852 226156 542904
rect 226208 542892 226214 542904
rect 253934 542892 253940 542904
rect 226208 542864 253940 542892
rect 226208 542852 226214 542864
rect 253934 542852 253940 542864
rect 253992 542852 253998 542904
rect 93670 542784 93676 542836
rect 93728 542824 93734 542836
rect 96246 542824 96252 542836
rect 93728 542796 96252 542824
rect 93728 542784 93734 542796
rect 96246 542784 96252 542796
rect 96304 542784 96310 542836
rect 99282 542784 99288 542836
rect 99340 542824 99346 542836
rect 106642 542824 106648 542836
rect 99340 542796 106648 542824
rect 99340 542784 99346 542796
rect 106642 542784 106648 542796
rect 106700 542784 106706 542836
rect 110322 542784 110328 542836
rect 110380 542824 110386 542836
rect 125318 542824 125324 542836
rect 110380 542796 125324 542824
rect 110380 542784 110386 542796
rect 125318 542784 125324 542796
rect 125376 542784 125382 542836
rect 131482 542784 131488 542836
rect 131540 542824 131546 542836
rect 188338 542824 188344 542836
rect 131540 542796 188344 542824
rect 131540 542784 131546 542796
rect 188338 542784 188344 542796
rect 188396 542784 188402 542836
rect 223482 542784 223488 542836
rect 223540 542824 223546 542836
rect 249794 542824 249800 542836
rect 223540 542796 249800 542824
rect 223540 542784 223546 542796
rect 249794 542784 249800 542796
rect 249852 542784 249858 542836
rect 93762 542716 93768 542768
rect 93820 542756 93826 542768
rect 98362 542756 98368 542768
rect 93820 542728 98368 542756
rect 93820 542716 93826 542728
rect 98362 542716 98368 542728
rect 98420 542716 98426 542768
rect 107562 542716 107568 542768
rect 107620 542756 107626 542768
rect 121178 542756 121184 542768
rect 107620 542728 121184 542756
rect 107620 542716 107626 542728
rect 121178 542716 121184 542728
rect 121236 542716 121242 542768
rect 139854 542716 139860 542768
rect 139912 542756 139918 542768
rect 140682 542756 140688 542768
rect 139912 542728 140688 542756
rect 139912 542716 139918 542728
rect 140682 542716 140688 542728
rect 140740 542716 140746 542768
rect 140774 542716 140780 542768
rect 140832 542756 140838 542768
rect 159358 542756 159364 542768
rect 140832 542728 159364 542756
rect 140832 542716 140838 542728
rect 159358 542716 159364 542728
rect 159416 542716 159422 542768
rect 224678 542716 224684 542768
rect 224736 542756 224742 542768
rect 251910 542756 251916 542768
rect 224736 542728 251916 542756
rect 224736 542716 224742 542728
rect 251910 542716 251916 542728
rect 251968 542716 251974 542768
rect 69290 542648 69296 542700
rect 69348 542688 69354 542700
rect 70302 542688 70308 542700
rect 69348 542660 70308 542688
rect 69348 542648 69354 542660
rect 70302 542648 70308 542660
rect 70360 542648 70366 542700
rect 96522 542648 96528 542700
rect 96580 542688 96586 542700
rect 102502 542688 102508 542700
rect 96580 542660 102508 542688
rect 96580 542648 96586 542660
rect 102502 542648 102508 542660
rect 102560 542648 102566 542700
rect 104526 542688 104532 542700
rect 102612 542660 104532 542688
rect 83826 542580 83832 542632
rect 83884 542620 83890 542632
rect 85666 542620 85672 542632
rect 83884 542592 85672 542620
rect 83884 542580 83890 542592
rect 85666 542580 85672 542592
rect 85724 542580 85730 542632
rect 97902 542580 97908 542632
rect 97960 542620 97966 542632
rect 102612 542620 102640 542660
rect 104526 542648 104532 542660
rect 104584 542648 104590 542700
rect 106182 542648 106188 542700
rect 106240 542688 106246 542700
rect 119062 542688 119068 542700
rect 106240 542660 119068 542688
rect 106240 542648 106246 542660
rect 119062 542648 119068 542660
rect 119120 542648 119126 542700
rect 135714 542648 135720 542700
rect 135772 542688 135778 542700
rect 160738 542688 160744 542700
rect 135772 542660 160744 542688
rect 135772 542648 135778 542660
rect 160738 542648 160744 542660
rect 160796 542648 160802 542700
rect 220538 542648 220544 542700
rect 220596 542688 220602 542700
rect 245654 542688 245660 542700
rect 220596 542660 245660 542688
rect 220596 542648 220602 542660
rect 245654 542648 245660 542660
rect 245712 542648 245718 542700
rect 97960 542592 102640 542620
rect 97960 542580 97966 542592
rect 103422 542580 103428 542632
rect 103480 542620 103486 542632
rect 114922 542620 114928 542632
rect 103480 542592 114928 542620
rect 103480 542580 103486 542592
rect 114922 542580 114928 542592
rect 114980 542580 114986 542632
rect 222102 542580 222108 542632
rect 222160 542620 222166 542632
rect 247770 542620 247776 542632
rect 222160 542592 247776 542620
rect 222160 542580 222166 542592
rect 247770 542580 247776 542592
rect 247828 542580 247834 542632
rect 81710 542512 81716 542564
rect 81768 542552 81774 542564
rect 84194 542552 84200 542564
rect 81768 542524 84200 542552
rect 81768 542512 81774 542524
rect 84194 542512 84200 542524
rect 84252 542512 84258 542564
rect 104802 542512 104808 542564
rect 104860 542552 104866 542564
rect 117038 542552 117044 542564
rect 104860 542524 117044 542552
rect 104860 542512 104866 542524
rect 117038 542512 117044 542524
rect 117096 542512 117102 542564
rect 133598 542512 133604 542564
rect 133656 542552 133662 542564
rect 140774 542552 140780 542564
rect 133656 542524 140780 542552
rect 133656 542512 133662 542524
rect 140774 542512 140780 542524
rect 140832 542512 140838 542564
rect 217870 542512 217876 542564
rect 217928 542552 217934 542564
rect 241514 542552 241520 542564
rect 217928 542524 241520 542552
rect 217928 542512 217934 542524
rect 241514 542512 241520 542524
rect 241572 542512 241578 542564
rect 95142 542444 95148 542496
rect 95200 542484 95206 542496
rect 100386 542484 100392 542496
rect 95200 542456 100392 542484
rect 95200 542444 95206 542456
rect 100386 542444 100392 542456
rect 100444 542444 100450 542496
rect 101950 542444 101956 542496
rect 102008 542484 102014 542496
rect 112806 542484 112812 542496
rect 102008 542456 112812 542484
rect 102008 542444 102014 542456
rect 112806 542444 112812 542456
rect 112864 542444 112870 542496
rect 219342 542444 219348 542496
rect 219400 542484 219406 542496
rect 243538 542484 243544 542496
rect 219400 542456 243544 542484
rect 219400 542444 219406 542456
rect 243538 542444 243544 542456
rect 243596 542444 243602 542496
rect 102042 542376 102048 542428
rect 102100 542416 102106 542428
rect 110782 542416 110788 542428
rect 102100 542388 110788 542416
rect 102100 542376 102106 542388
rect 110782 542376 110788 542388
rect 110840 542376 110846 542428
rect 211154 540948 211160 541000
rect 211212 540988 211218 541000
rect 211430 540988 211436 541000
rect 211212 540960 211436 540988
rect 211212 540948 211218 540960
rect 211430 540948 211436 540960
rect 211488 540948 211494 541000
rect 56778 540268 56784 540320
rect 56836 540308 56842 540320
rect 137278 540308 137284 540320
rect 56836 540280 137284 540308
rect 56836 540268 56842 540280
rect 137278 540268 137284 540280
rect 137336 540268 137342 540320
rect 56686 540200 56692 540252
rect 56744 540240 56750 540252
rect 170030 540240 170036 540252
rect 56744 540212 170036 540240
rect 56744 540200 56750 540212
rect 170030 540200 170036 540212
rect 170088 540200 170094 540252
rect 56870 539180 56876 539232
rect 56928 539220 56934 539232
rect 299750 539220 299756 539232
rect 56928 539192 299756 539220
rect 56928 539180 56934 539192
rect 299750 539180 299756 539192
rect 299808 539180 299814 539232
rect 59722 539112 59728 539164
rect 59780 539152 59786 539164
rect 429470 539152 429476 539164
rect 59780 539124 429476 539152
rect 59780 539112 59786 539124
rect 429470 539112 429476 539124
rect 429528 539112 429534 539164
rect 59630 539044 59636 539096
rect 59688 539084 59694 539096
rect 559190 539084 559196 539096
rect 59688 539056 559196 539084
rect 59688 539044 59694 539056
rect 559190 539044 559196 539056
rect 559248 539044 559254 539096
rect 57974 538976 57980 539028
rect 58032 539016 58038 539028
rect 580350 539016 580356 539028
rect 58032 538988 580356 539016
rect 58032 538976 58038 538988
rect 580350 538976 580356 538988
rect 580408 538976 580414 539028
rect 58066 538908 58072 538960
rect 58124 538948 58130 538960
rect 580626 538948 580632 538960
rect 58124 538920 580632 538948
rect 58124 538908 58130 538920
rect 580626 538908 580632 538920
rect 580684 538908 580690 538960
rect 57054 538840 57060 538892
rect 57112 538880 57118 538892
rect 580534 538880 580540 538892
rect 57112 538852 580540 538880
rect 57112 538840 57118 538852
rect 580534 538840 580540 538852
rect 580592 538840 580598 538892
rect 2958 538364 2964 538416
rect 3016 538404 3022 538416
rect 5350 538404 5356 538416
rect 3016 538376 5356 538404
rect 3016 538364 3022 538376
rect 5350 538364 5356 538376
rect 5408 538364 5414 538416
rect 60734 538364 60740 538416
rect 60792 538404 60798 538416
rect 541618 538404 541624 538416
rect 60792 538376 541624 538404
rect 60792 538364 60798 538376
rect 541618 538364 541624 538376
rect 541676 538364 541682 538416
rect 59998 538296 60004 538348
rect 60056 538336 60062 538348
rect 563698 538336 563704 538348
rect 60056 538308 563704 538336
rect 60056 538296 60062 538308
rect 563698 538296 563704 538308
rect 563756 538296 563762 538348
rect 19978 538228 19984 538280
rect 20036 538268 20042 538280
rect 57238 538268 57244 538280
rect 20036 538240 57244 538268
rect 20036 538228 20042 538240
rect 57238 538228 57244 538240
rect 57296 538228 57302 538280
rect 58158 538228 58164 538280
rect 58216 538268 58222 538280
rect 579798 538268 579804 538280
rect 58216 538240 579804 538268
rect 58216 538228 58222 538240
rect 579798 538228 579804 538240
rect 579856 538228 579862 538280
rect 57146 537888 57152 537940
rect 57204 537928 57210 537940
rect 580258 537928 580264 537940
rect 57204 537900 580264 537928
rect 57204 537888 57210 537900
rect 580258 537888 580264 537900
rect 580316 537888 580322 537940
rect 48958 536800 48964 536852
rect 49016 536840 49022 536852
rect 57238 536840 57244 536852
rect 49016 536812 57244 536840
rect 49016 536800 49022 536812
rect 57238 536800 57244 536812
rect 57296 536800 57302 536852
rect 60090 536800 60096 536852
rect 60148 536840 60154 536852
rect 60734 536840 60740 536852
rect 60148 536812 60740 536840
rect 60148 536800 60154 536812
rect 60734 536800 60740 536812
rect 60792 536800 60798 536852
rect 282822 536732 282828 536784
rect 282880 536772 282886 536784
rect 467098 536772 467104 536784
rect 282880 536744 467104 536772
rect 282880 536732 282886 536744
rect 467098 536732 467104 536744
rect 467156 536732 467162 536784
rect 282822 535372 282828 535424
rect 282880 535412 282886 535424
rect 465718 535412 465724 535424
rect 282880 535384 465724 535412
rect 282880 535372 282886 535384
rect 465718 535372 465724 535384
rect 465776 535372 465782 535424
rect 4798 534080 4804 534132
rect 4856 534120 4862 534132
rect 57238 534120 57244 534132
rect 4856 534092 57244 534120
rect 4856 534080 4862 534092
rect 57238 534080 57244 534092
rect 57296 534080 57302 534132
rect 282822 532652 282828 532704
rect 282880 532692 282886 532704
rect 464338 532692 464344 532704
rect 282880 532664 464344 532692
rect 282880 532652 282886 532664
rect 464338 532652 464344 532664
rect 464396 532652 464402 532704
rect 53098 531360 53104 531412
rect 53156 531400 53162 531412
rect 57238 531400 57244 531412
rect 53156 531372 57244 531400
rect 53156 531360 53162 531372
rect 57238 531360 57244 531372
rect 57296 531360 57302 531412
rect 282822 531224 282828 531276
rect 282880 531264 282886 531276
rect 356790 531264 356796 531276
rect 282880 531236 356796 531264
rect 282880 531224 282886 531236
rect 356790 531224 356796 531236
rect 356848 531224 356854 531276
rect 541618 530544 541624 530596
rect 541676 530584 541682 530596
rect 556154 530584 556160 530596
rect 541676 530556 556160 530584
rect 541676 530544 541682 530556
rect 556154 530544 556160 530556
rect 556212 530544 556218 530596
rect 563698 530000 563704 530052
rect 563756 530040 563762 530052
rect 563756 530012 565860 530040
rect 563756 530000 563762 530012
rect 46198 529932 46204 529984
rect 46256 529972 46262 529984
rect 57238 529972 57244 529984
rect 46256 529944 57244 529972
rect 46256 529932 46262 529944
rect 57238 529932 57244 529944
rect 57296 529932 57302 529984
rect 565832 529904 565860 530012
rect 569218 529904 569224 529916
rect 565832 529876 569224 529904
rect 569218 529864 569224 529876
rect 569276 529864 569282 529916
rect 556154 529184 556160 529236
rect 556212 529224 556218 529236
rect 568482 529224 568488 529236
rect 556212 529196 568488 529224
rect 556212 529184 556218 529196
rect 568482 529184 568488 529196
rect 568540 529184 568546 529236
rect 282822 528504 282828 528556
rect 282880 528544 282886 528556
rect 356698 528544 356704 528556
rect 282880 528516 356704 528544
rect 282880 528504 282886 528516
rect 356698 528504 356704 528516
rect 356756 528504 356762 528556
rect 4890 527144 4896 527196
rect 4948 527184 4954 527196
rect 57238 527184 57244 527196
rect 4948 527156 57244 527184
rect 4948 527144 4954 527156
rect 57238 527144 57244 527156
rect 57296 527144 57302 527196
rect 17218 525784 17224 525836
rect 17276 525824 17282 525836
rect 57238 525824 57244 525836
rect 17276 525796 57244 525824
rect 17276 525784 17282 525796
rect 57238 525784 57244 525796
rect 57296 525784 57302 525836
rect 568482 525784 568488 525836
rect 568540 525824 568546 525836
rect 568540 525796 568620 525824
rect 568540 525784 568546 525796
rect 282822 525716 282828 525768
rect 282880 525756 282886 525768
rect 355318 525756 355324 525768
rect 282880 525728 355324 525756
rect 282880 525716 282886 525728
rect 355318 525716 355324 525728
rect 355376 525716 355382 525768
rect 568592 525756 568620 525796
rect 571978 525756 571984 525768
rect 568592 525728 571984 525756
rect 571978 525716 571984 525728
rect 572036 525716 572042 525768
rect 282822 524356 282828 524408
rect 282880 524396 282886 524408
rect 354030 524396 354036 524408
rect 282880 524368 354036 524396
rect 282880 524356 282886 524368
rect 354030 524356 354036 524368
rect 354088 524356 354094 524408
rect 43438 522996 43444 523048
rect 43496 523036 43502 523048
rect 57238 523036 57244 523048
rect 43496 523008 57244 523036
rect 43496 522996 43502 523008
rect 57238 522996 57244 523008
rect 57296 522996 57302 523048
rect 4982 521636 4988 521688
rect 5040 521676 5046 521688
rect 57238 521676 57244 521688
rect 5040 521648 57244 521676
rect 5040 521636 5046 521648
rect 57238 521636 57244 521648
rect 57296 521636 57302 521688
rect 282822 521568 282828 521620
rect 282880 521608 282886 521620
rect 353938 521608 353944 521620
rect 282880 521580 353944 521608
rect 282880 521568 282886 521580
rect 353938 521568 353944 521580
rect 353996 521568 354002 521620
rect 569218 521568 569224 521620
rect 569276 521608 569282 521620
rect 570966 521608 570972 521620
rect 569276 521580 570972 521608
rect 569276 521568 569282 521580
rect 570966 521568 570972 521580
rect 571024 521568 571030 521620
rect 282822 520208 282828 520260
rect 282880 520248 282886 520260
rect 352742 520248 352748 520260
rect 282880 520220 352748 520248
rect 282880 520208 282886 520220
rect 352742 520208 352748 520220
rect 352800 520208 352806 520260
rect 51718 518916 51724 518968
rect 51776 518956 51782 518968
rect 57238 518956 57244 518968
rect 51776 518928 57244 518956
rect 51776 518916 51782 518928
rect 57238 518916 57244 518928
rect 57296 518916 57302 518968
rect 35158 517488 35164 517540
rect 35216 517528 35222 517540
rect 57238 517528 57244 517540
rect 35216 517500 57244 517528
rect 35216 517488 35222 517500
rect 57238 517488 57244 517500
rect 57296 517488 57302 517540
rect 570966 517488 570972 517540
rect 571024 517528 571030 517540
rect 571024 517500 571380 517528
rect 571024 517488 571030 517500
rect 281902 517420 281908 517472
rect 281960 517460 281966 517472
rect 352650 517460 352656 517472
rect 281960 517432 352656 517460
rect 281960 517420 281966 517432
rect 352650 517420 352656 517432
rect 352708 517420 352714 517472
rect 571352 517460 571380 517500
rect 573358 517460 573364 517472
rect 571352 517432 573364 517460
rect 573358 517420 573364 517432
rect 573416 517420 573422 517472
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 57238 514808 57244 514820
rect 3476 514780 57244 514808
rect 3476 514768 3482 514780
rect 57238 514768 57244 514780
rect 57296 514768 57302 514820
rect 282822 514700 282828 514752
rect 282880 514740 282886 514752
rect 352558 514740 352564 514752
rect 282880 514712 352564 514740
rect 282880 514700 282886 514712
rect 352558 514700 352564 514712
rect 352616 514700 352622 514752
rect 50338 513340 50344 513392
rect 50396 513380 50402 513392
rect 57238 513380 57244 513392
rect 50396 513352 57244 513380
rect 50396 513340 50402 513352
rect 57238 513340 57244 513352
rect 57296 513340 57302 513392
rect 282086 513272 282092 513324
rect 282144 513312 282150 513324
rect 476206 513312 476212 513324
rect 282144 513284 476212 513312
rect 282144 513272 282150 513284
rect 476206 513272 476212 513284
rect 476264 513272 476270 513324
rect 571978 513272 571984 513324
rect 572036 513312 572042 513324
rect 574738 513312 574744 513324
rect 572036 513284 574744 513312
rect 572036 513272 572042 513284
rect 574738 513272 574744 513284
rect 574796 513272 574802 513324
rect 33778 510620 33784 510672
rect 33836 510660 33842 510672
rect 57238 510660 57244 510672
rect 33836 510632 57244 510660
rect 33836 510620 33842 510632
rect 57238 510620 57244 510632
rect 57296 510620 57302 510672
rect 282822 510552 282828 510604
rect 282880 510592 282886 510604
rect 474734 510592 474740 510604
rect 282880 510564 474740 510592
rect 282880 510552 282886 510564
rect 474734 510552 474740 510564
rect 474792 510552 474798 510604
rect 2774 509532 2780 509584
rect 2832 509572 2838 509584
rect 5442 509572 5448 509584
rect 2832 509544 5448 509572
rect 2832 509532 2838 509544
rect 5442 509532 5448 509544
rect 5500 509532 5506 509584
rect 3510 509260 3516 509312
rect 3568 509300 3574 509312
rect 57238 509300 57244 509312
rect 3568 509272 57244 509300
rect 3568 509260 3574 509272
rect 57238 509260 57244 509272
rect 57296 509260 57302 509312
rect 282270 509192 282276 509244
rect 282328 509232 282334 509244
rect 473354 509232 473360 509244
rect 282328 509204 473360 509232
rect 282328 509192 282334 509204
rect 473354 509192 473360 509204
rect 473412 509192 473418 509244
rect 574738 507764 574744 507816
rect 574796 507804 574802 507816
rect 577958 507804 577964 507816
rect 574796 507776 577964 507804
rect 574796 507764 574802 507776
rect 577958 507764 577964 507776
rect 578016 507764 578022 507816
rect 39390 506472 39396 506524
rect 39448 506512 39454 506524
rect 57238 506512 57244 506524
rect 39448 506484 57244 506512
rect 39448 506472 39454 506484
rect 57238 506472 57244 506484
rect 57296 506472 57302 506524
rect 281902 506404 281908 506456
rect 281960 506444 281966 506456
rect 471974 506444 471980 506456
rect 281960 506416 471980 506444
rect 281960 506404 281966 506416
rect 471974 506404 471980 506416
rect 472032 506404 472038 506456
rect 577958 506268 577964 506320
rect 578016 506308 578022 506320
rect 580258 506308 580264 506320
rect 578016 506280 580264 506308
rect 578016 506268 578022 506280
rect 580258 506268 580264 506280
rect 580316 506268 580322 506320
rect 28258 505112 28264 505164
rect 28316 505152 28322 505164
rect 57238 505152 57244 505164
rect 28316 505124 57244 505152
rect 28316 505112 28322 505124
rect 57238 505112 57244 505124
rect 57296 505112 57302 505164
rect 282822 503616 282828 503668
rect 282880 503656 282886 503668
rect 470594 503656 470600 503668
rect 282880 503628 470600 503656
rect 282880 503616 282886 503628
rect 470594 503616 470600 503628
rect 470652 503616 470658 503668
rect 3602 502324 3608 502376
rect 3660 502364 3666 502376
rect 57238 502364 57244 502376
rect 3660 502336 57244 502364
rect 3660 502324 3666 502336
rect 57238 502324 57244 502336
rect 57296 502324 57302 502376
rect 282086 502256 282092 502308
rect 282144 502296 282150 502308
rect 469214 502296 469220 502308
rect 282144 502268 469220 502296
rect 282144 502256 282150 502268
rect 469214 502256 469220 502268
rect 469272 502256 469278 502308
rect 37918 500964 37924 501016
rect 37976 501004 37982 501016
rect 57238 501004 57244 501016
rect 37976 500976 57244 501004
rect 37976 500964 37982 500976
rect 57238 500964 57244 500976
rect 57296 500964 57302 501016
rect 573358 499536 573364 499588
rect 573416 499576 573422 499588
rect 573416 499548 574140 499576
rect 573416 499536 573422 499548
rect 282822 499468 282828 499520
rect 282880 499508 282886 499520
rect 467926 499508 467932 499520
rect 282880 499480 467932 499508
rect 282880 499468 282886 499480
rect 467926 499468 467932 499480
rect 467984 499468 467990 499520
rect 574112 499508 574140 499548
rect 576762 499508 576768 499520
rect 574112 499480 576768 499508
rect 576762 499468 576768 499480
rect 576820 499468 576826 499520
rect 20070 498176 20076 498228
rect 20128 498216 20134 498228
rect 57238 498216 57244 498228
rect 20128 498188 57244 498216
rect 20128 498176 20134 498188
rect 57238 498176 57244 498188
rect 57296 498176 57302 498228
rect 282270 498108 282276 498160
rect 282328 498148 282334 498160
rect 467834 498148 467840 498160
rect 282328 498120 467840 498148
rect 282328 498108 282334 498120
rect 467834 498108 467840 498120
rect 467892 498108 467898 498160
rect 281902 495388 281908 495440
rect 281960 495428 281966 495440
rect 466454 495428 466460 495440
rect 281960 495400 466460 495428
rect 281960 495388 281966 495400
rect 466454 495388 466460 495400
rect 466512 495388 466518 495440
rect 32398 494028 32404 494080
rect 32456 494068 32462 494080
rect 57238 494068 57244 494080
rect 32456 494040 57244 494068
rect 32456 494028 32462 494040
rect 57238 494028 57244 494040
rect 57296 494028 57302 494080
rect 282454 493960 282460 494012
rect 282512 494000 282518 494012
rect 465074 494000 465080 494012
rect 282512 493972 465080 494000
rect 282512 493960 282518 493972
rect 465074 493960 465080 493972
rect 465132 493960 465138 494012
rect 576854 493824 576860 493876
rect 576912 493864 576918 493876
rect 578878 493864 578884 493876
rect 576912 493836 578884 493864
rect 576912 493824 576918 493836
rect 578878 493824 578884 493836
rect 578936 493824 578942 493876
rect 17310 491308 17316 491360
rect 17368 491348 17374 491360
rect 57238 491348 57244 491360
rect 17368 491320 57244 491348
rect 17368 491308 17374 491320
rect 57238 491308 57244 491320
rect 57296 491308 57302 491360
rect 282086 491240 282092 491292
rect 282144 491280 282150 491292
rect 463694 491280 463700 491292
rect 282144 491252 463700 491280
rect 282144 491240 282150 491252
rect 463694 491240 463700 491252
rect 463752 491240 463758 491292
rect 56962 491172 56968 491224
rect 57020 491212 57026 491224
rect 57238 491212 57244 491224
rect 57020 491184 57244 491212
rect 57020 491172 57026 491184
rect 57238 491172 57244 491184
rect 57296 491172 57302 491224
rect 282822 488452 282828 488504
rect 282880 488492 282886 488504
rect 462314 488492 462320 488504
rect 282880 488464 462320 488492
rect 282880 488452 282886 488464
rect 462314 488452 462320 488464
rect 462372 488452 462378 488504
rect 3694 487160 3700 487212
rect 3752 487200 3758 487212
rect 56594 487200 56600 487212
rect 3752 487172 56600 487200
rect 3752 487160 3758 487172
rect 56594 487160 56600 487172
rect 56652 487160 56658 487212
rect 282822 487092 282828 487144
rect 282880 487132 282886 487144
rect 461026 487132 461032 487144
rect 282880 487104 461032 487132
rect 282880 487092 282886 487104
rect 461026 487092 461032 487104
rect 461084 487092 461090 487144
rect 15838 485800 15844 485852
rect 15896 485840 15902 485852
rect 56594 485840 56600 485852
rect 15896 485812 56600 485840
rect 15896 485800 15902 485812
rect 56594 485800 56600 485812
rect 56652 485800 56658 485852
rect 282822 484304 282828 484356
rect 282880 484344 282886 484356
rect 460934 484344 460940 484356
rect 282880 484316 460940 484344
rect 282880 484304 282886 484316
rect 460934 484304 460940 484316
rect 460992 484304 460998 484356
rect 3786 483012 3792 483064
rect 3844 483052 3850 483064
rect 56594 483052 56600 483064
rect 3844 483024 56600 483052
rect 3844 483012 3850 483024
rect 56594 483012 56600 483024
rect 56652 483012 56658 483064
rect 282454 482944 282460 482996
rect 282512 482984 282518 482996
rect 443638 482984 443644 482996
rect 282512 482956 443644 482984
rect 282512 482944 282518 482956
rect 443638 482944 443644 482956
rect 443696 482944 443702 482996
rect 4062 481652 4068 481704
rect 4120 481692 4126 481704
rect 56594 481692 56600 481704
rect 4120 481664 56600 481692
rect 4120 481652 4126 481664
rect 56594 481652 56600 481664
rect 56652 481652 56658 481704
rect 3234 480632 3240 480684
rect 3292 480672 3298 480684
rect 5534 480672 5540 480684
rect 3292 480644 5540 480672
rect 3292 480632 3298 480644
rect 5534 480632 5540 480644
rect 5592 480632 5598 480684
rect 282086 480156 282092 480208
rect 282144 480196 282150 480208
rect 359550 480196 359556 480208
rect 282144 480168 359556 480196
rect 282144 480156 282150 480168
rect 359550 480156 359556 480168
rect 359608 480156 359614 480208
rect 3970 478864 3976 478916
rect 4028 478904 4034 478916
rect 56594 478904 56600 478916
rect 4028 478876 56600 478904
rect 4028 478864 4034 478876
rect 56594 478864 56600 478876
rect 56652 478864 56658 478916
rect 282822 477436 282828 477488
rect 282880 477476 282886 477488
rect 359458 477476 359464 477488
rect 282880 477448 359464 477476
rect 282880 477436 282886 477448
rect 359458 477436 359464 477448
rect 359516 477436 359522 477488
rect 3326 476008 3332 476060
rect 3384 476048 3390 476060
rect 56594 476048 56600 476060
rect 3384 476020 56600 476048
rect 3384 476008 3390 476020
rect 56594 476008 56600 476020
rect 56652 476008 56658 476060
rect 282546 476008 282552 476060
rect 282604 476048 282610 476060
rect 358170 476048 358176 476060
rect 282604 476020 358176 476048
rect 282604 476008 282610 476020
rect 358170 476008 358176 476020
rect 358228 476008 358234 476060
rect 5534 474648 5540 474700
rect 5592 474688 5598 474700
rect 56594 474688 56600 474700
rect 5592 474660 56600 474688
rect 5592 474648 5598 474660
rect 56594 474648 56600 474660
rect 56652 474648 56658 474700
rect 282086 473288 282092 473340
rect 282144 473328 282150 473340
rect 358078 473328 358084 473340
rect 282144 473300 358084 473328
rect 282144 473288 282150 473300
rect 358078 473288 358084 473300
rect 358136 473288 358142 473340
rect 5442 471928 5448 471980
rect 5500 471968 5506 471980
rect 56594 471968 56600 471980
rect 5500 471940 56600 471968
rect 5500 471928 5506 471940
rect 56594 471928 56600 471940
rect 56652 471928 56658 471980
rect 282454 471928 282460 471980
rect 282512 471968 282518 471980
rect 349798 471968 349804 471980
rect 282512 471940 349804 471968
rect 282512 471928 282518 471940
rect 349798 471928 349804 471940
rect 349856 471928 349862 471980
rect 3878 470500 3884 470552
rect 3936 470540 3942 470552
rect 56502 470540 56508 470552
rect 3936 470512 56508 470540
rect 3936 470500 3942 470512
rect 56502 470500 56508 470512
rect 56560 470500 56566 470552
rect 282086 469140 282092 469192
rect 282144 469180 282150 469192
rect 452746 469180 452752 469192
rect 282144 469152 452752 469180
rect 282144 469140 282150 469152
rect 452746 469140 452752 469152
rect 452804 469140 452810 469192
rect 5350 467780 5356 467832
rect 5408 467820 5414 467832
rect 56502 467820 56508 467832
rect 5408 467792 56508 467820
rect 5408 467780 5414 467792
rect 56502 467780 56508 467792
rect 56560 467780 56566 467832
rect 5258 466352 5264 466404
rect 5316 466392 5322 466404
rect 56502 466392 56508 466404
rect 5316 466364 56508 466392
rect 5316 466352 5322 466364
rect 56502 466352 56508 466364
rect 56560 466352 56566 466404
rect 282822 466352 282828 466404
rect 282880 466392 282886 466404
rect 330478 466392 330484 466404
rect 282880 466364 330484 466392
rect 282880 466352 282886 466364
rect 330478 466352 330484 466364
rect 330536 466352 330542 466404
rect 282270 464992 282276 465044
rect 282328 465032 282334 465044
rect 329282 465032 329288 465044
rect 282328 465004 329288 465032
rect 282328 464992 282334 465004
rect 329282 464992 329288 465004
rect 329340 464992 329346 465044
rect 31018 463632 31024 463684
rect 31076 463672 31082 463684
rect 56502 463672 56508 463684
rect 31076 463644 56508 463672
rect 31076 463632 31082 463644
rect 56502 463632 56508 463644
rect 56560 463632 56566 463684
rect 14458 462272 14464 462324
rect 14516 462312 14522 462324
rect 56502 462312 56508 462324
rect 14516 462284 56508 462312
rect 14516 462272 14522 462284
rect 56502 462272 56508 462284
rect 56560 462272 56566 462324
rect 282822 462272 282828 462324
rect 282880 462312 282886 462324
rect 329098 462312 329104 462324
rect 282880 462284 329104 462312
rect 282880 462272 282886 462284
rect 329098 462272 329104 462284
rect 329156 462272 329162 462324
rect 576854 462000 576860 462052
rect 576912 462040 576918 462052
rect 579982 462040 579988 462052
rect 576912 462012 579988 462040
rect 576912 462000 576918 462012
rect 579982 462000 579988 462012
rect 580040 462000 580046 462052
rect 282454 460844 282460 460896
rect 282512 460884 282518 460896
rect 327718 460884 327724 460896
rect 282512 460856 327724 460884
rect 282512 460844 282518 460856
rect 327718 460844 327724 460856
rect 327776 460844 327782 460896
rect 571794 459552 571800 459604
rect 571852 459592 571858 459604
rect 576854 459592 576860 459604
rect 571852 459564 576860 459592
rect 571852 459552 571858 459564
rect 576854 459552 576860 459564
rect 576912 459552 576918 459604
rect 5166 459484 5172 459536
rect 5224 459524 5230 459536
rect 56594 459524 56600 459536
rect 5224 459496 56600 459524
rect 5224 459484 5230 459496
rect 56594 459484 56600 459496
rect 56652 459484 56658 459536
rect 282086 458124 282092 458176
rect 282144 458164 282150 458176
rect 326338 458164 326344 458176
rect 282144 458136 326344 458164
rect 282144 458124 282150 458136
rect 326338 458124 326344 458136
rect 326396 458124 326402 458176
rect 21358 456696 21364 456748
rect 21416 456736 21422 456748
rect 56594 456736 56600 456748
rect 21416 456708 56600 456736
rect 21416 456696 21422 456708
rect 56594 456696 56600 456708
rect 56652 456696 56658 456748
rect 566458 456016 566464 456068
rect 566516 456056 566522 456068
rect 571794 456056 571800 456068
rect 566516 456028 571800 456056
rect 566516 456016 566522 456028
rect 571794 456016 571800 456028
rect 571852 456016 571858 456068
rect 13078 455336 13084 455388
rect 13136 455376 13142 455388
rect 56594 455376 56600 455388
rect 13136 455348 56600 455376
rect 13136 455336 13142 455348
rect 56594 455336 56600 455348
rect 56652 455336 56658 455388
rect 282822 455336 282828 455388
rect 282880 455376 282886 455388
rect 324958 455376 324964 455388
rect 282880 455348 324964 455376
rect 282880 455336 282886 455348
rect 324958 455336 324964 455348
rect 325016 455336 325022 455388
rect 282822 453976 282828 454028
rect 282880 454016 282886 454028
rect 323670 454016 323676 454028
rect 282880 453988 323676 454016
rect 282880 453976 282886 453988
rect 323670 453976 323676 453988
rect 323728 453976 323734 454028
rect 5074 452480 5080 452532
rect 5132 452520 5138 452532
rect 56594 452520 56600 452532
rect 5132 452492 56600 452520
rect 5132 452480 5138 452492
rect 56594 452480 56600 452492
rect 56652 452480 56658 452532
rect 3326 452344 3332 452396
rect 3384 452384 3390 452396
rect 56502 452384 56508 452396
rect 3384 452356 56508 452384
rect 3384 452344 3390 452356
rect 56502 452344 56508 452356
rect 56560 452344 56566 452396
rect 24762 451188 24768 451240
rect 24820 451228 24826 451240
rect 56594 451228 56600 451240
rect 24820 451200 56600 451228
rect 24820 451188 24826 451200
rect 56594 451188 56600 451200
rect 56652 451188 56658 451240
rect 282822 451188 282828 451240
rect 282880 451228 282886 451240
rect 322290 451228 322296 451240
rect 282880 451200 322296 451228
rect 282880 451188 282886 451200
rect 322290 451188 322296 451200
rect 322348 451188 322354 451240
rect 282454 449828 282460 449880
rect 282512 449868 282518 449880
rect 460382 449868 460388 449880
rect 282512 449840 460388 449868
rect 282512 449828 282518 449840
rect 460382 449828 460388 449840
rect 460440 449828 460446 449880
rect 56594 448604 56600 448656
rect 56652 448644 56658 448656
rect 57514 448644 57520 448656
rect 56652 448616 57520 448644
rect 56652 448604 56658 448616
rect 57514 448604 57520 448616
rect 57572 448604 57578 448656
rect 10318 448468 10324 448520
rect 10376 448508 10382 448520
rect 57514 448508 57520 448520
rect 10376 448480 57520 448508
rect 10376 448468 10382 448480
rect 57514 448468 57520 448480
rect 57572 448468 57578 448520
rect 42058 447040 42064 447092
rect 42116 447080 42122 447092
rect 57514 447080 57520 447092
rect 42116 447052 57520 447080
rect 42116 447040 42122 447052
rect 57514 447040 57520 447052
rect 57572 447040 57578 447092
rect 282822 447040 282828 447092
rect 282880 447080 282886 447092
rect 460198 447080 460204 447092
rect 282880 447052 460204 447080
rect 282880 447040 282886 447052
rect 460198 447040 460204 447052
rect 460256 447040 460262 447092
rect 566458 445788 566464 445800
rect 564452 445760 566464 445788
rect 563238 445680 563244 445732
rect 563296 445720 563302 445732
rect 564452 445720 564480 445760
rect 566458 445748 566464 445760
rect 566516 445748 566522 445800
rect 563296 445692 564480 445720
rect 563296 445680 563302 445692
rect 282822 444320 282828 444372
rect 282880 444360 282886 444372
rect 458818 444360 458824 444372
rect 282880 444332 458824 444360
rect 282880 444320 282886 444332
rect 458818 444320 458824 444332
rect 458876 444320 458882 444372
rect 282822 442892 282828 442944
rect 282880 442932 282886 442944
rect 457438 442932 457444 442944
rect 282880 442904 457444 442932
rect 282880 442892 282886 442904
rect 457438 442892 457444 442904
rect 457496 442892 457502 442944
rect 562410 442144 562416 442196
rect 562468 442184 562474 442196
rect 563238 442184 563244 442196
rect 562468 442156 563244 442184
rect 562468 442144 562474 442156
rect 563238 442144 563244 442156
rect 563296 442144 563302 442196
rect 578602 440240 578608 440292
rect 578660 440280 578666 440292
rect 580258 440280 580264 440292
rect 578660 440252 580264 440280
rect 578660 440240 578666 440252
rect 580258 440240 580264 440252
rect 580316 440240 580322 440292
rect 282822 440172 282828 440224
rect 282880 440212 282886 440224
rect 456058 440212 456064 440224
rect 282880 440184 456064 440212
rect 282880 440172 282886 440184
rect 456058 440172 456064 440184
rect 456116 440172 456122 440224
rect 560938 438880 560944 438932
rect 560996 438920 561002 438932
rect 562410 438920 562416 438932
rect 560996 438892 562416 438920
rect 560996 438880 561002 438892
rect 562410 438880 562416 438892
rect 562468 438880 562474 438932
rect 576118 438880 576124 438932
rect 576176 438920 576182 438932
rect 578602 438920 578608 438932
rect 576176 438892 578608 438920
rect 576176 438880 576182 438892
rect 578602 438880 578608 438892
rect 578660 438880 578666 438932
rect 282454 438812 282460 438864
rect 282512 438852 282518 438864
rect 454678 438852 454684 438864
rect 282512 438824 454684 438852
rect 282512 438812 282518 438824
rect 454678 438812 454684 438824
rect 454736 438812 454742 438864
rect 577958 437588 577964 437640
rect 578016 437628 578022 437640
rect 579614 437628 579620 437640
rect 578016 437600 579620 437628
rect 578016 437588 578022 437600
rect 579614 437588 579620 437600
rect 579672 437588 579678 437640
rect 282822 436024 282828 436076
rect 282880 436064 282886 436076
rect 453482 436064 453488 436076
rect 282880 436036 453488 436064
rect 282880 436024 282886 436036
rect 453482 436024 453488 436036
rect 453540 436024 453546 436076
rect 575842 435480 575848 435532
rect 575900 435520 575906 435532
rect 577958 435520 577964 435532
rect 575900 435492 577964 435520
rect 575900 435480 575906 435492
rect 577958 435480 577964 435492
rect 578016 435480 578022 435532
rect 57606 433984 57612 434036
rect 57664 434024 57670 434036
rect 60090 434024 60096 434036
rect 57664 433996 60096 434024
rect 57664 433984 57670 433996
rect 60090 433984 60096 433996
rect 60148 433984 60154 434036
rect 282822 433236 282828 433288
rect 282880 433276 282886 433288
rect 453298 433276 453304 433288
rect 282880 433248 453304 433276
rect 282880 433236 282886 433248
rect 453298 433236 453304 433248
rect 453356 433236 453362 433288
rect 574738 432488 574744 432540
rect 574796 432528 574802 432540
rect 575842 432528 575848 432540
rect 574796 432500 575848 432528
rect 574796 432488 574802 432500
rect 575842 432488 575848 432500
rect 575900 432488 575906 432540
rect 282822 431876 282828 431928
rect 282880 431916 282886 431928
rect 291930 431916 291936 431928
rect 282880 431888 291936 431916
rect 282880 431876 282886 431888
rect 291930 431876 291936 431888
rect 291988 431876 291994 431928
rect 58710 429156 58716 429208
rect 58768 429196 58774 429208
rect 59998 429196 60004 429208
rect 58768 429168 60004 429196
rect 58768 429156 58774 429168
rect 59998 429156 60004 429168
rect 60056 429156 60062 429208
rect 282822 429088 282828 429140
rect 282880 429128 282886 429140
rect 290550 429128 290556 429140
rect 282880 429100 290556 429128
rect 282880 429088 282886 429100
rect 290550 429088 290556 429100
rect 290608 429088 290614 429140
rect 570598 426776 570604 426828
rect 570656 426816 570662 426828
rect 576118 426816 576124 426828
rect 570656 426788 576124 426816
rect 570656 426776 570662 426788
rect 576118 426776 576124 426788
rect 576176 426776 576182 426828
rect 282822 426572 282828 426624
rect 282880 426612 282886 426624
rect 287698 426612 287704 426624
rect 282880 426584 287704 426612
rect 282880 426572 282886 426584
rect 287698 426572 287704 426584
rect 287756 426572 287762 426624
rect 282454 425008 282460 425060
rect 282512 425048 282518 425060
rect 286318 425048 286324 425060
rect 282512 425020 286324 425048
rect 282512 425008 282518 425020
rect 286318 425008 286324 425020
rect 286376 425008 286382 425060
rect 570782 422696 570788 422748
rect 570840 422736 570846 422748
rect 574738 422736 574744 422748
rect 570840 422708 574744 422736
rect 570840 422696 570846 422708
rect 574738 422696 574744 422708
rect 574796 422696 574802 422748
rect 282086 422220 282092 422272
rect 282144 422260 282150 422272
rect 284938 422260 284944 422272
rect 282144 422232 284944 422260
rect 282144 422220 282150 422232
rect 284938 422220 284944 422232
rect 284996 422220 285002 422272
rect 281718 420792 281724 420844
rect 281776 420832 281782 420844
rect 283558 420832 283564 420844
rect 281776 420804 283564 420832
rect 281776 420792 281782 420804
rect 283558 420792 283564 420804
rect 283616 420792 283622 420844
rect 567838 419500 567844 419552
rect 567896 419540 567902 419552
rect 570782 419540 570788 419552
rect 567896 419512 570788 419540
rect 567896 419500 567902 419512
rect 570782 419500 570788 419512
rect 570840 419500 570846 419552
rect 558178 418140 558184 418192
rect 558236 418180 558242 418192
rect 560938 418180 560944 418192
rect 558236 418152 560944 418180
rect 558236 418140 558242 418152
rect 560938 418140 560944 418152
rect 560996 418140 561002 418192
rect 282822 418072 282828 418124
rect 282880 418112 282886 418124
rect 294598 418112 294604 418124
rect 282880 418084 294604 418112
rect 282880 418072 282886 418084
rect 294598 418072 294604 418084
rect 294656 418072 294662 418124
rect 282822 416712 282828 416764
rect 282880 416752 282886 416764
rect 316034 416752 316040 416764
rect 282880 416724 316040 416752
rect 282880 416712 282886 416724
rect 316034 416712 316040 416724
rect 316092 416712 316098 416764
rect 57698 413924 57704 413976
rect 57756 413964 57762 413976
rect 58710 413964 58716 413976
rect 57756 413936 58716 413964
rect 57756 413924 57762 413936
rect 58710 413924 58716 413936
rect 58768 413924 58774 413976
rect 281902 413924 281908 413976
rect 281960 413964 281966 413976
rect 399478 413964 399484 413976
rect 281960 413936 399484 413964
rect 281960 413924 281966 413936
rect 399478 413924 399484 413936
rect 399536 413924 399542 413976
rect 282822 411204 282828 411256
rect 282880 411244 282886 411256
rect 398098 411244 398104 411256
rect 282880 411216 398104 411244
rect 282880 411204 282886 411216
rect 398098 411204 398104 411216
rect 398156 411204 398162 411256
rect 282086 409776 282092 409828
rect 282144 409816 282150 409828
rect 395338 409816 395344 409828
rect 282144 409788 395344 409816
rect 282144 409776 282150 409788
rect 395338 409776 395344 409788
rect 395396 409776 395402 409828
rect 282822 407056 282828 407108
rect 282880 407096 282886 407108
rect 393958 407096 393964 407108
rect 282880 407068 393964 407096
rect 282880 407056 282886 407068
rect 393958 407056 393964 407068
rect 394016 407056 394022 407108
rect 578970 405696 578976 405748
rect 579028 405736 579034 405748
rect 580258 405736 580264 405748
rect 579028 405708 580264 405736
rect 579028 405696 579034 405708
rect 580258 405696 580264 405708
rect 580316 405696 580322 405748
rect 282822 405628 282828 405680
rect 282880 405668 282886 405680
rect 392578 405668 392584 405680
rect 282880 405640 392584 405668
rect 282880 405628 282886 405640
rect 392578 405628 392584 405640
rect 392636 405628 392642 405680
rect 577590 403520 577596 403572
rect 577648 403560 577654 403572
rect 578970 403560 578976 403572
rect 577648 403532 578976 403560
rect 577648 403520 577654 403532
rect 578970 403520 578976 403532
rect 579028 403520 579034 403572
rect 281902 402908 281908 402960
rect 281960 402948 281966 402960
rect 391198 402948 391204 402960
rect 281960 402920 391204 402948
rect 281960 402908 281966 402920
rect 391198 402908 391204 402920
rect 391256 402908 391262 402960
rect 577498 400188 577504 400240
rect 577556 400228 577562 400240
rect 580902 400228 580908 400240
rect 577556 400200 580908 400228
rect 577556 400188 577562 400200
rect 580902 400188 580908 400200
rect 580960 400188 580966 400240
rect 282822 400120 282828 400172
rect 282880 400160 282886 400172
rect 388438 400160 388444 400172
rect 282880 400132 388444 400160
rect 282880 400120 282886 400132
rect 388438 400120 388444 400132
rect 388496 400120 388502 400172
rect 556798 399644 556804 399696
rect 556856 399684 556862 399696
rect 558178 399684 558184 399696
rect 556856 399656 558184 399684
rect 556856 399644 556862 399656
rect 558178 399644 558184 399656
rect 558236 399644 558242 399696
rect 282086 398760 282092 398812
rect 282144 398800 282150 398812
rect 445754 398800 445760 398812
rect 282144 398772 445760 398800
rect 282144 398760 282150 398772
rect 445754 398760 445760 398772
rect 445812 398760 445818 398812
rect 282086 395836 282092 395888
rect 282144 395876 282150 395888
rect 285030 395876 285036 395888
rect 282144 395848 285036 395876
rect 282144 395836 282150 395848
rect 285030 395836 285036 395848
rect 285088 395836 285094 395888
rect 282270 394612 282276 394664
rect 282328 394652 282334 394664
rect 402238 394652 402244 394664
rect 282328 394624 402244 394652
rect 282328 394612 282334 394624
rect 402238 394612 402244 394624
rect 402296 394612 402302 394664
rect 569218 394612 569224 394664
rect 569276 394652 569282 394664
rect 570598 394652 570604 394664
rect 569276 394624 570604 394652
rect 569276 394612 569282 394624
rect 570598 394612 570604 394624
rect 570656 394612 570662 394664
rect 566550 391960 566556 392012
rect 566608 392000 566614 392012
rect 567838 392000 567844 392012
rect 566608 391972 567844 392000
rect 566608 391960 566614 391972
rect 567838 391960 567844 391972
rect 567896 391960 567902 392012
rect 577866 391960 577872 392012
rect 577924 392000 577930 392012
rect 579614 392000 579620 392012
rect 577924 391972 579620 392000
rect 577924 391960 577930 391972
rect 579614 391960 579620 391972
rect 579672 391960 579678 392012
rect 281902 391892 281908 391944
rect 281960 391932 281966 391944
rect 320266 391932 320272 391944
rect 281960 391904 320272 391932
rect 281960 391892 281966 391904
rect 320266 391892 320272 391904
rect 320324 391892 320330 391944
rect 574094 390600 574100 390652
rect 574152 390640 574158 390652
rect 577590 390640 577596 390652
rect 574152 390612 577596 390640
rect 574152 390600 574158 390612
rect 577590 390600 577596 390612
rect 577648 390600 577654 390652
rect 282454 389784 282460 389836
rect 282512 389824 282518 389836
rect 286410 389824 286416 389836
rect 282512 389796 286416 389824
rect 282512 389784 282518 389796
rect 286410 389784 286416 389796
rect 286468 389784 286474 389836
rect 282086 387744 282092 387796
rect 282144 387784 282150 387796
rect 318794 387784 318800 387796
rect 282144 387756 318800 387784
rect 282144 387744 282150 387756
rect 318794 387744 318800 387756
rect 318852 387744 318858 387796
rect 555418 387744 555424 387796
rect 555476 387784 555482 387796
rect 556798 387784 556804 387796
rect 555476 387756 556804 387784
rect 555476 387744 555482 387756
rect 556798 387744 556804 387756
rect 556856 387744 556862 387796
rect 571978 387132 571984 387184
rect 572036 387172 572042 387184
rect 574094 387172 574100 387184
rect 572036 387144 574100 387172
rect 572036 387132 572042 387144
rect 574094 387132 574100 387144
rect 574152 387132 574158 387184
rect 576210 385024 576216 385076
rect 576268 385064 576274 385076
rect 577866 385064 577872 385076
rect 576268 385036 577872 385064
rect 576268 385024 576274 385036
rect 577866 385024 577872 385036
rect 577924 385024 577930 385076
rect 282822 384616 282828 384668
rect 282880 384656 282886 384668
rect 287790 384656 287796 384668
rect 282880 384628 287796 384656
rect 282880 384616 282886 384628
rect 287790 384616 287796 384628
rect 287848 384616 287854 384668
rect 282822 383596 282828 383648
rect 282880 383636 282886 383648
rect 450538 383636 450544 383648
rect 282880 383608 450544 383636
rect 282880 383596 282886 383608
rect 450538 383596 450544 383608
rect 450596 383596 450602 383648
rect 567378 382236 567384 382288
rect 567436 382276 567442 382288
rect 571978 382276 571984 382288
rect 567436 382248 571984 382276
rect 567436 382236 567442 382248
rect 571978 382236 571984 382248
rect 572036 382236 572042 382288
rect 574094 382236 574100 382288
rect 574152 382276 574158 382288
rect 576210 382276 576216 382288
rect 574152 382248 576216 382276
rect 574152 382236 574158 382248
rect 576210 382236 576216 382248
rect 576268 382236 576274 382288
rect 282822 380808 282828 380860
rect 282880 380848 282886 380860
rect 449158 380848 449164 380860
rect 282880 380820 449164 380848
rect 282880 380808 282886 380820
rect 449158 380808 449164 380820
rect 449216 380808 449222 380860
rect 282454 379448 282460 379500
rect 282512 379488 282518 379500
rect 447778 379488 447784 379500
rect 282512 379460 447784 379488
rect 282512 379448 282518 379460
rect 447778 379448 447784 379460
rect 447836 379448 447842 379500
rect 566642 377680 566648 377732
rect 566700 377720 566706 377732
rect 567378 377720 567384 377732
rect 566700 377692 567384 377720
rect 566700 377680 566706 377692
rect 567378 377680 567384 377692
rect 567436 377680 567442 377732
rect 282086 376660 282092 376712
rect 282144 376700 282150 376712
rect 446398 376700 446404 376712
rect 282144 376672 446404 376700
rect 282144 376660 282150 376672
rect 446398 376660 446404 376672
rect 446456 376660 446462 376712
rect 570966 376320 570972 376372
rect 571024 376360 571030 376372
rect 574094 376360 574100 376372
rect 571024 376332 574100 376360
rect 571024 376320 571030 376332
rect 574094 376320 574100 376332
rect 574152 376320 574158 376372
rect 282822 373940 282828 373992
rect 282880 373980 282886 373992
rect 358814 373980 358820 373992
rect 282880 373952 358820 373980
rect 282880 373940 282886 373952
rect 358814 373940 358820 373952
rect 358872 373940 358878 373992
rect 282546 372512 282552 372564
rect 282604 372552 282610 372564
rect 357434 372552 357440 372564
rect 282604 372524 357440 372552
rect 282604 372512 282610 372524
rect 357434 372512 357440 372524
rect 357492 372512 357498 372564
rect 566458 371696 566464 371748
rect 566516 371736 566522 371748
rect 569218 371736 569224 371748
rect 566516 371708 569224 371736
rect 566516 371696 566522 371708
rect 569218 371696 569224 371708
rect 569276 371696 569282 371748
rect 568758 371560 568764 371612
rect 568816 371600 568822 371612
rect 570966 371600 570972 371612
rect 568816 371572 570972 371600
rect 568816 371560 568822 371572
rect 570966 371560 570972 371572
rect 571024 371560 571030 371612
rect 565262 369860 565268 369912
rect 565320 369900 565326 369912
rect 566642 369900 566648 369912
rect 565320 369872 566648 369900
rect 565320 369860 565326 369872
rect 566642 369860 566648 369872
rect 566700 369860 566706 369912
rect 568758 369900 568764 369912
rect 566752 369872 568764 369900
rect 282822 369792 282828 369844
rect 282880 369832 282886 369844
rect 356054 369832 356060 369844
rect 282880 369804 356060 369832
rect 282880 369792 282886 369804
rect 356054 369792 356060 369804
rect 356112 369792 356118 369844
rect 564066 369792 564072 369844
rect 564124 369832 564130 369844
rect 566752 369832 566780 369872
rect 568758 369860 568764 369872
rect 568816 369860 568822 369912
rect 564124 369804 566780 369832
rect 564124 369792 564130 369804
rect 282454 368432 282460 368484
rect 282512 368472 282518 368484
rect 354766 368472 354772 368484
rect 282512 368444 354772 368472
rect 282512 368432 282518 368444
rect 354766 368432 354772 368444
rect 354824 368432 354830 368484
rect 563698 368432 563704 368484
rect 563756 368472 563762 368484
rect 566550 368472 566556 368484
rect 563756 368444 566556 368472
rect 563756 368432 563762 368444
rect 566550 368432 566556 368444
rect 566608 368432 566614 368484
rect 563790 368024 563796 368076
rect 563848 368064 563854 368076
rect 565262 368064 565268 368076
rect 563848 368036 565268 368064
rect 563848 368024 563854 368036
rect 565262 368024 565268 368036
rect 565320 368024 565326 368076
rect 560938 367072 560944 367124
rect 560996 367112 561002 367124
rect 564066 367112 564072 367124
rect 560996 367084 564072 367112
rect 560996 367072 561002 367084
rect 564066 367072 564072 367084
rect 564124 367072 564130 367124
rect 577590 367072 577596 367124
rect 577648 367112 577654 367124
rect 579522 367112 579528 367124
rect 577648 367084 579528 367112
rect 577648 367072 577654 367084
rect 579522 367072 579528 367084
rect 579580 367072 579586 367124
rect 2958 367004 2964 367056
rect 3016 367044 3022 367056
rect 15838 367044 15844 367056
rect 3016 367016 15844 367044
rect 3016 367004 3022 367016
rect 15838 367004 15844 367016
rect 15896 367004 15902 367056
rect 282086 365644 282092 365696
rect 282144 365684 282150 365696
rect 353294 365684 353300 365696
rect 282144 365656 353300 365684
rect 282144 365644 282150 365656
rect 353294 365644 353300 365656
rect 353352 365644 353358 365696
rect 282822 362856 282828 362908
rect 282880 362896 282886 362908
rect 352006 362896 352012 362908
rect 282880 362868 352012 362896
rect 282880 362856 282886 362868
rect 352006 362856 352012 362868
rect 352064 362856 352070 362908
rect 282546 361496 282552 361548
rect 282604 361536 282610 361548
rect 352190 361536 352196 361548
rect 282604 361508 352196 361536
rect 282604 361496 282610 361508
rect 352190 361496 352196 361508
rect 352248 361496 352254 361548
rect 553302 360816 553308 360868
rect 553360 360856 553366 360868
rect 563790 360856 563796 360868
rect 553360 360828 563796 360856
rect 553360 360816 553366 360828
rect 563790 360816 563796 360828
rect 563848 360816 563854 360868
rect 282822 358708 282828 358760
rect 282880 358748 282886 358760
rect 350534 358748 350540 358760
rect 282880 358720 350540 358748
rect 282880 358708 282886 358720
rect 350534 358708 350540 358720
rect 350592 358708 350598 358760
rect 282454 357348 282460 357400
rect 282512 357388 282518 357400
rect 349154 357388 349160 357400
rect 282512 357360 349160 357388
rect 282512 357348 282518 357360
rect 349154 357348 349160 357360
rect 349212 357348 349218 357400
rect 562410 357008 562416 357060
rect 562468 357048 562474 357060
rect 563698 357048 563704 357060
rect 562468 357020 563704 357048
rect 562468 357008 562474 357020
rect 563698 357008 563704 357020
rect 563756 357008 563762 357060
rect 551278 356600 551284 356652
rect 551336 356640 551342 356652
rect 553302 356640 553308 356652
rect 551336 356612 553308 356640
rect 551336 356600 551342 356612
rect 553302 356600 553308 356612
rect 553360 356600 553366 356652
rect 576854 356056 576860 356108
rect 576912 356096 576918 356108
rect 579522 356096 579528 356108
rect 576912 356068 579528 356096
rect 576912 356056 576918 356068
rect 579522 356056 579528 356068
rect 579580 356056 579586 356108
rect 574738 354696 574744 354748
rect 574796 354736 574802 354748
rect 577498 354736 577504 354748
rect 574796 354708 577504 354736
rect 574796 354696 574802 354708
rect 577498 354696 577504 354708
rect 577556 354696 577562 354748
rect 282086 354628 282092 354680
rect 282144 354668 282150 354680
rect 347774 354668 347780 354680
rect 282144 354640 347780 354668
rect 282144 354628 282150 354640
rect 347774 354628 347780 354640
rect 347832 354628 347838 354680
rect 571978 353404 571984 353456
rect 572036 353444 572042 353456
rect 576854 353444 576860 353456
rect 572036 353416 576860 353444
rect 572036 353404 572042 353416
rect 576854 353404 576860 353416
rect 576912 353404 576918 353456
rect 549254 351908 549260 351960
rect 549312 351948 549318 351960
rect 551278 351948 551284 351960
rect 549312 351920 551284 351948
rect 549312 351908 549318 351920
rect 551278 351908 551284 351920
rect 551336 351908 551342 351960
rect 554038 351908 554044 351960
rect 554096 351948 554102 351960
rect 555418 351948 555424 351960
rect 554096 351920 555424 351948
rect 554096 351908 554102 351920
rect 555418 351908 555424 351920
rect 555476 351908 555482 351960
rect 282822 351840 282828 351892
rect 282880 351880 282886 351892
rect 346394 351880 346400 351892
rect 282880 351852 346400 351880
rect 282880 351840 282886 351852
rect 346394 351840 346400 351852
rect 346452 351840 346458 351892
rect 561030 350548 561036 350600
rect 561088 350588 561094 350600
rect 562410 350588 562416 350600
rect 561088 350560 562416 350588
rect 561088 350548 561094 350560
rect 562410 350548 562416 350560
rect 562468 350548 562474 350600
rect 282546 350480 282552 350532
rect 282604 350520 282610 350532
rect 345014 350520 345020 350532
rect 282604 350492 345020 350520
rect 282604 350480 282610 350492
rect 345014 350480 345020 350492
rect 345072 350480 345078 350532
rect 564434 349800 564440 349852
rect 564492 349840 564498 349852
rect 571978 349840 571984 349852
rect 564492 349812 571984 349840
rect 564492 349800 564498 349812
rect 571978 349800 571984 349812
rect 572036 349800 572042 349852
rect 559558 348372 559564 348424
rect 559616 348412 559622 348424
rect 560938 348412 560944 348424
rect 559616 348384 560944 348412
rect 559616 348372 559622 348384
rect 560938 348372 560944 348384
rect 560996 348372 561002 348424
rect 282822 347692 282828 347744
rect 282880 347732 282886 347744
rect 343726 347732 343732 347744
rect 282880 347704 343732 347732
rect 282880 347692 282886 347704
rect 343726 347692 343732 347704
rect 343784 347692 343790 347744
rect 561674 347420 561680 347472
rect 561732 347460 561738 347472
rect 564434 347460 564440 347472
rect 561732 347432 564440 347460
rect 561732 347420 561738 347432
rect 564434 347420 564440 347432
rect 564492 347420 564498 347472
rect 573358 347420 573364 347472
rect 573416 347460 573422 347472
rect 574738 347460 574744 347472
rect 573416 347432 574744 347460
rect 573416 347420 573422 347432
rect 574738 347420 574744 347432
rect 574796 347420 574802 347472
rect 282454 346332 282460 346384
rect 282512 346372 282518 346384
rect 343634 346372 343640 346384
rect 282512 346344 343640 346372
rect 282512 346332 282518 346344
rect 343634 346332 343640 346344
rect 343692 346332 343698 346384
rect 548518 345856 548524 345908
rect 548576 345896 548582 345908
rect 549254 345896 549260 345908
rect 548576 345868 549260 345896
rect 548576 345856 548582 345868
rect 549254 345856 549260 345868
rect 549312 345856 549318 345908
rect 574094 345040 574100 345092
rect 574152 345080 574158 345092
rect 577590 345080 577596 345092
rect 574152 345052 577596 345080
rect 574152 345040 574158 345052
rect 577590 345040 577596 345052
rect 577648 345040 577654 345092
rect 559650 343612 559656 343664
rect 559708 343652 559714 343664
rect 561030 343652 561036 343664
rect 559708 343624 561036 343652
rect 559708 343612 559714 343624
rect 561030 343612 561036 343624
rect 561088 343612 561094 343664
rect 561674 343652 561680 343664
rect 561140 343624 561680 343652
rect 282822 343544 282828 343596
rect 282880 343584 282886 343596
rect 342254 343584 342260 343596
rect 282880 343556 342260 343584
rect 282880 343544 282886 343556
rect 342254 343544 342260 343556
rect 342312 343544 342318 343596
rect 558454 343544 558460 343596
rect 558512 343584 558518 343596
rect 561140 343584 561168 343624
rect 561674 343612 561680 343624
rect 561732 343612 561738 343664
rect 558512 343556 561168 343584
rect 558512 343544 558518 343556
rect 552658 342252 552664 342304
rect 552716 342292 552722 342304
rect 554038 342292 554044 342304
rect 552716 342264 554044 342292
rect 552716 342252 552722 342264
rect 554038 342252 554044 342264
rect 554096 342252 554102 342304
rect 553394 340892 553400 340944
rect 553452 340932 553458 340944
rect 558454 340932 558460 340944
rect 553452 340904 558460 340932
rect 553452 340892 553458 340904
rect 558454 340892 558460 340904
rect 558512 340892 558518 340944
rect 571426 340892 571432 340944
rect 571484 340932 571490 340944
rect 574094 340932 574100 340944
rect 571484 340904 574100 340932
rect 571484 340892 571490 340904
rect 574094 340892 574100 340904
rect 574152 340892 574158 340944
rect 282822 340824 282828 340876
rect 282880 340864 282886 340876
rect 340874 340864 340880 340876
rect 282880 340836 340880 340864
rect 282880 340824 282886 340836
rect 340874 340824 340880 340836
rect 340932 340824 340938 340876
rect 578878 340144 578884 340196
rect 578936 340184 578942 340196
rect 580166 340184 580172 340196
rect 578936 340156 580172 340184
rect 578936 340144 578942 340156
rect 580166 340144 580172 340156
rect 580224 340144 580230 340196
rect 57054 339396 57060 339448
rect 57112 339436 57118 339448
rect 58710 339436 58716 339448
rect 57112 339408 58716 339436
rect 57112 339396 57118 339408
rect 58710 339396 58716 339408
rect 58768 339396 58774 339448
rect 282822 339396 282828 339448
rect 282880 339436 282886 339448
rect 339494 339436 339500 339448
rect 282880 339408 339500 339436
rect 282880 339396 282886 339408
rect 339494 339396 339500 339408
rect 339552 339396 339558 339448
rect 563422 338648 563428 338700
rect 563480 338688 563486 338700
rect 566458 338688 566464 338700
rect 563480 338660 566464 338688
rect 563480 338648 563486 338660
rect 566458 338648 566464 338660
rect 566516 338648 566522 338700
rect 551370 338104 551376 338156
rect 551428 338144 551434 338156
rect 553394 338144 553400 338156
rect 551428 338116 553400 338144
rect 551428 338104 551434 338116
rect 553394 338104 553400 338116
rect 553452 338104 553458 338156
rect 3326 338036 3332 338088
rect 3384 338076 3390 338088
rect 56962 338076 56968 338088
rect 3384 338048 56968 338076
rect 3384 338036 3390 338048
rect 56962 338036 56968 338048
rect 57020 338036 57026 338088
rect 57698 336676 57704 336728
rect 57756 336716 57762 336728
rect 58618 336716 58624 336728
rect 57756 336688 58624 336716
rect 57756 336676 57762 336688
rect 58618 336676 58624 336688
rect 58676 336676 58682 336728
rect 282822 336676 282828 336728
rect 282880 336716 282886 336728
rect 338114 336716 338120 336728
rect 282880 336688 338120 336716
rect 282880 336676 282886 336688
rect 338114 336676 338120 336688
rect 338172 336676 338178 336728
rect 561766 336608 561772 336660
rect 561824 336648 561830 336660
rect 563422 336648 563428 336660
rect 561824 336620 563428 336648
rect 561824 336608 561830 336620
rect 563422 336608 563428 336620
rect 563480 336608 563486 336660
rect 570966 336336 570972 336388
rect 571024 336376 571030 336388
rect 571426 336376 571432 336388
rect 571024 336348 571432 336376
rect 571024 336336 571030 336348
rect 571426 336336 571432 336348
rect 571484 336336 571490 336388
rect 282362 335248 282368 335300
rect 282420 335288 282426 335300
rect 336826 335288 336832 335300
rect 282420 335260 336832 335288
rect 282420 335248 282426 335260
rect 336826 335248 336832 335260
rect 336884 335248 336890 335300
rect 551278 333956 551284 334008
rect 551336 333996 551342 334008
rect 552658 333996 552664 334008
rect 551336 333968 552664 333996
rect 551336 333956 551342 333968
rect 552658 333956 552664 333968
rect 552716 333956 552722 334008
rect 558822 333956 558828 334008
rect 558880 333996 558886 334008
rect 561766 333996 561772 334008
rect 558880 333968 561772 333996
rect 558880 333956 558886 333968
rect 561766 333956 561772 333968
rect 561824 333956 561830 334008
rect 282822 332528 282828 332580
rect 282880 332568 282886 332580
rect 336734 332568 336740 332580
rect 282880 332540 336740 332568
rect 282880 332528 282886 332540
rect 336734 332528 336740 332540
rect 336792 332528 336798 332580
rect 57146 331576 57152 331628
rect 57204 331616 57210 331628
rect 58802 331616 58808 331628
rect 57204 331588 58808 331616
rect 57204 331576 57210 331588
rect 58802 331576 58808 331588
rect 58860 331576 58866 331628
rect 556798 331440 556804 331492
rect 556856 331480 556862 331492
rect 558822 331480 558828 331492
rect 556856 331452 558828 331480
rect 556856 331440 556862 331452
rect 558822 331440 558828 331452
rect 558880 331440 558886 331492
rect 567838 331304 567844 331356
rect 567896 331344 567902 331356
rect 570966 331344 570972 331356
rect 567896 331316 570972 331344
rect 567896 331304 567902 331316
rect 570966 331304 570972 331316
rect 571024 331304 571030 331356
rect 546494 331168 546500 331220
rect 546552 331208 546558 331220
rect 548518 331208 548524 331220
rect 546552 331180 548524 331208
rect 546552 331168 546558 331180
rect 548518 331168 548524 331180
rect 548576 331168 548582 331220
rect 57330 330488 57336 330540
rect 57388 330528 57394 330540
rect 57698 330528 57704 330540
rect 57388 330500 57704 330528
rect 57388 330488 57394 330500
rect 57698 330488 57704 330500
rect 57756 330488 57762 330540
rect 565078 330080 565084 330132
rect 565136 330120 565142 330132
rect 567838 330120 567844 330132
rect 565136 330092 567844 330120
rect 565136 330080 565142 330092
rect 567838 330080 567844 330092
rect 567896 330080 567902 330132
rect 282822 329740 282828 329792
rect 282880 329780 282886 329792
rect 335354 329780 335360 329792
rect 282880 329752 335360 329780
rect 282880 329740 282886 329752
rect 335354 329740 335360 329752
rect 335412 329740 335418 329792
rect 57422 328380 57428 328432
rect 57480 328420 57486 328432
rect 58894 328420 58900 328432
rect 57480 328392 58900 328420
rect 57480 328380 57486 328392
rect 58894 328380 58900 328392
rect 58952 328380 58958 328432
rect 282822 328380 282828 328432
rect 282880 328420 282886 328432
rect 333974 328420 333980 328432
rect 282880 328392 333980 328420
rect 282880 328380 282886 328392
rect 333974 328380 333980 328392
rect 334032 328380 334038 328432
rect 576854 328380 576860 328432
rect 576912 328420 576918 328432
rect 578878 328420 578884 328432
rect 576912 328392 578884 328420
rect 576912 328380 576918 328392
rect 578878 328380 578884 328392
rect 578936 328380 578942 328432
rect 549346 328108 549352 328160
rect 549404 328148 549410 328160
rect 551370 328148 551376 328160
rect 549404 328120 551376 328148
rect 549404 328108 549410 328120
rect 551370 328108 551376 328120
rect 551428 328108 551434 328160
rect 549254 327700 549260 327752
rect 549312 327740 549318 327752
rect 559650 327740 559656 327752
rect 549312 327712 559656 327740
rect 549312 327700 549318 327712
rect 559650 327700 559656 327712
rect 559708 327700 559714 327752
rect 57698 327020 57704 327072
rect 57756 327060 57762 327072
rect 58986 327060 58992 327072
rect 57756 327032 58992 327060
rect 57756 327020 57762 327032
rect 58986 327020 58992 327032
rect 59044 327020 59050 327072
rect 546494 325700 546500 325712
rect 545132 325672 546500 325700
rect 282822 325592 282828 325644
rect 282880 325632 282886 325644
rect 332594 325632 332600 325644
rect 282880 325604 332600 325632
rect 282880 325592 282886 325604
rect 332594 325592 332600 325604
rect 332652 325592 332658 325644
rect 543734 325592 543740 325644
rect 543792 325632 543798 325644
rect 545132 325632 545160 325672
rect 546494 325660 546500 325672
rect 546552 325660 546558 325712
rect 543792 325604 545160 325632
rect 543792 325592 543798 325604
rect 552658 325320 552664 325372
rect 552716 325360 552722 325372
rect 559558 325360 559564 325372
rect 552716 325332 559564 325360
rect 552716 325320 552722 325332
rect 559558 325320 559564 325332
rect 559616 325320 559622 325372
rect 545114 324300 545120 324352
rect 545172 324340 545178 324352
rect 549346 324340 549352 324352
rect 545172 324312 549352 324340
rect 545172 324300 545178 324312
rect 549346 324300 549352 324312
rect 549404 324300 549410 324352
rect 553394 324300 553400 324352
rect 553452 324340 553458 324352
rect 556798 324340 556804 324352
rect 553452 324312 556804 324340
rect 553452 324300 553458 324312
rect 556798 324300 556804 324312
rect 556856 324300 556862 324352
rect 3050 324232 3056 324284
rect 3108 324272 3114 324284
rect 32398 324272 32404 324284
rect 3108 324244 32404 324272
rect 3108 324232 3114 324244
rect 32398 324232 32404 324244
rect 32456 324232 32462 324284
rect 282362 324232 282368 324284
rect 282420 324272 282426 324284
rect 290458 324272 290464 324284
rect 282420 324244 290464 324272
rect 282420 324232 282426 324244
rect 290458 324232 290464 324244
rect 290516 324232 290522 324284
rect 535454 323552 535460 323604
rect 535512 323592 535518 323604
rect 543734 323592 543740 323604
rect 535512 323564 543740 323592
rect 535512 323552 535518 323564
rect 543734 323552 543740 323564
rect 543792 323552 543798 323604
rect 57790 322940 57796 322992
rect 57848 322980 57854 322992
rect 59078 322980 59084 322992
rect 57848 322952 59084 322980
rect 57848 322940 57854 322952
rect 59078 322940 59084 322952
rect 59136 322940 59142 322992
rect 549162 322940 549168 322992
rect 549220 322980 549226 322992
rect 552658 322980 552664 322992
rect 549220 322952 552664 322980
rect 549220 322940 549226 322952
rect 552658 322940 552664 322952
rect 552716 322940 552722 322992
rect 57606 322056 57612 322108
rect 57664 322096 57670 322108
rect 59262 322096 59268 322108
rect 57664 322068 59268 322096
rect 57664 322056 57670 322068
rect 59262 322056 59268 322068
rect 59320 322056 59326 322108
rect 532878 321580 532884 321632
rect 532936 321620 532942 321632
rect 535454 321620 535460 321632
rect 532936 321592 535460 321620
rect 532936 321580 532942 321592
rect 535454 321580 535460 321592
rect 535512 321580 535518 321632
rect 549254 321620 549260 321632
rect 546512 321592 549260 321620
rect 282822 321512 282828 321564
rect 282880 321552 282886 321564
rect 329926 321552 329932 321564
rect 282880 321524 329932 321552
rect 282880 321512 282886 321524
rect 329926 321512 329932 321524
rect 329984 321512 329990 321564
rect 544102 321444 544108 321496
rect 544160 321484 544166 321496
rect 546512 321484 546540 321592
rect 549254 321580 549260 321592
rect 549312 321580 549318 321632
rect 544160 321456 546540 321484
rect 544160 321444 544166 321456
rect 548518 320696 548524 320748
rect 548576 320736 548582 320748
rect 551278 320736 551284 320748
rect 548576 320708 551284 320736
rect 548576 320696 548582 320708
rect 551278 320696 551284 320708
rect 551336 320696 551342 320748
rect 542998 320152 543004 320204
rect 543056 320192 543062 320204
rect 545114 320192 545120 320204
rect 543056 320164 545120 320192
rect 543056 320152 543062 320164
rect 545114 320152 545120 320164
rect 545172 320152 545178 320204
rect 56594 320084 56600 320136
rect 56652 320124 56658 320136
rect 58526 320124 58532 320136
rect 56652 320096 58532 320124
rect 56652 320084 56658 320096
rect 58526 320084 58532 320096
rect 58584 320084 58590 320136
rect 546494 319744 546500 319796
rect 546552 319784 546558 319796
rect 549162 319784 549168 319796
rect 546552 319756 549168 319784
rect 546552 319744 546558 319756
rect 549162 319744 549168 319756
rect 549220 319744 549226 319796
rect 549898 319472 549904 319524
rect 549956 319512 549962 319524
rect 553394 319512 553400 319524
rect 549956 319484 553400 319512
rect 549956 319472 549962 319484
rect 553394 319472 553400 319484
rect 553452 319472 553458 319524
rect 529566 319200 529572 319252
rect 529624 319240 529630 319252
rect 532878 319240 532884 319252
rect 529624 319212 532884 319240
rect 529624 319200 529630 319212
rect 532878 319200 532884 319212
rect 532936 319200 532942 319252
rect 574830 318792 574836 318844
rect 574888 318832 574894 318844
rect 576762 318832 576768 318844
rect 574888 318804 576768 318832
rect 574888 318792 574894 318804
rect 576762 318792 576768 318804
rect 576820 318792 576826 318844
rect 282822 318724 282828 318776
rect 282880 318764 282886 318776
rect 291838 318764 291844 318776
rect 282880 318736 291844 318764
rect 282880 318724 282886 318736
rect 291838 318724 291844 318736
rect 291896 318724 291902 318776
rect 57790 317880 57796 317892
rect 57440 317852 57796 317880
rect 57440 317268 57468 317852
rect 57790 317840 57796 317852
rect 57848 317840 57854 317892
rect 57514 317364 57520 317416
rect 57572 317404 57578 317416
rect 58434 317404 58440 317416
rect 57572 317376 58440 317404
rect 57572 317364 57578 317376
rect 58434 317364 58440 317376
rect 58492 317364 58498 317416
rect 282822 317364 282828 317416
rect 282880 317404 282886 317416
rect 322198 317404 322204 317416
rect 282880 317376 322204 317404
rect 282880 317364 282886 317376
rect 322198 317364 322204 317376
rect 322256 317364 322262 317416
rect 57514 317268 57520 317280
rect 57440 317240 57520 317268
rect 57514 317228 57520 317240
rect 57572 317228 57578 317280
rect 572714 317024 572720 317076
rect 572772 317064 572778 317076
rect 574830 317064 574836 317076
rect 572772 317036 574836 317064
rect 572772 317024 572778 317036
rect 574830 317024 574836 317036
rect 574888 317024 574894 317076
rect 542078 316956 542084 317008
rect 542136 316996 542142 317008
rect 544102 316996 544108 317008
rect 542136 316968 544108 316996
rect 542136 316956 542142 316968
rect 544102 316956 544108 316968
rect 544160 316956 544166 317008
rect 545206 316616 545212 316668
rect 545264 316656 545270 316668
rect 546494 316656 546500 316668
rect 545264 316628 546500 316656
rect 545264 316616 545270 316628
rect 546494 316616 546500 316628
rect 546552 316616 546558 316668
rect 529566 316044 529572 316056
rect 524432 316016 529572 316044
rect 56594 315936 56600 315988
rect 56652 315976 56658 315988
rect 57514 315976 57520 315988
rect 56652 315948 57520 315976
rect 56652 315936 56658 315948
rect 57514 315936 57520 315948
rect 57572 315936 57578 315988
rect 523494 315936 523500 315988
rect 523552 315976 523558 315988
rect 524432 315976 524460 316016
rect 529566 316004 529572 316016
rect 529624 316004 529630 316056
rect 523552 315948 524460 315976
rect 523552 315936 523558 315948
rect 57698 315800 57704 315852
rect 57756 315840 57762 315852
rect 57974 315840 57980 315852
rect 57756 315812 57980 315840
rect 57756 315800 57762 315812
rect 57974 315800 57980 315812
rect 58032 315800 58038 315852
rect 59078 314644 59084 314696
rect 59136 314684 59142 314696
rect 59998 314684 60004 314696
rect 59136 314656 60004 314684
rect 59136 314644 59142 314656
rect 59998 314644 60004 314656
rect 60056 314644 60062 314696
rect 560938 314644 560944 314696
rect 560996 314684 561002 314696
rect 565078 314684 565084 314696
rect 560996 314656 565084 314684
rect 560996 314644 561002 314656
rect 565078 314644 565084 314656
rect 565136 314644 565142 314696
rect 282822 314576 282828 314628
rect 282880 314616 282886 314628
rect 327074 314616 327080 314628
rect 282880 314588 327080 314616
rect 282880 314576 282886 314588
rect 327074 314576 327080 314588
rect 327132 314576 327138 314628
rect 282362 313216 282368 313268
rect 282420 313256 282426 313268
rect 325694 313256 325700 313268
rect 282420 313228 325700 313256
rect 282420 313216 282426 313228
rect 325694 313216 325700 313228
rect 325752 313216 325758 313268
rect 539962 311924 539968 311976
rect 540020 311964 540026 311976
rect 542078 311964 542084 311976
rect 540020 311936 542084 311964
rect 540020 311924 540026 311936
rect 542078 311924 542084 311936
rect 542136 311924 542142 311976
rect 545206 311896 545212 311908
rect 543752 311868 545212 311896
rect 543090 311788 543096 311840
rect 543148 311828 543154 311840
rect 543752 311828 543780 311868
rect 545206 311856 545212 311868
rect 545264 311856 545270 311908
rect 573358 311896 573364 311908
rect 569972 311868 573364 311896
rect 543148 311800 543780 311828
rect 543148 311788 543154 311800
rect 567930 311788 567936 311840
rect 567988 311828 567994 311840
rect 569972 311828 570000 311868
rect 573358 311856 573364 311868
rect 573416 311856 573422 311908
rect 567988 311800 570000 311828
rect 567988 311788 567994 311800
rect 535454 311108 535460 311160
rect 535512 311148 535518 311160
rect 542998 311148 543004 311160
rect 535512 311120 543004 311148
rect 535512 311108 535518 311120
rect 542998 311108 543004 311120
rect 543056 311108 543062 311160
rect 545114 310972 545120 311024
rect 545172 311012 545178 311024
rect 549898 311012 549904 311024
rect 545172 310984 549904 311012
rect 545172 310972 545178 310984
rect 549898 310972 549904 310984
rect 549956 310972 549962 311024
rect 281902 310428 281908 310480
rect 281960 310468 281966 310480
rect 323578 310468 323584 310480
rect 281960 310440 323584 310468
rect 281960 310428 281966 310440
rect 323578 310428 323584 310440
rect 323636 310428 323642 310480
rect 563054 309952 563060 310004
rect 563112 309992 563118 310004
rect 567930 309992 567936 310004
rect 563112 309964 567936 309992
rect 563112 309952 563118 309964
rect 567930 309952 567936 309964
rect 567988 309952 567994 310004
rect 519538 309748 519544 309800
rect 519596 309788 519602 309800
rect 539962 309788 539968 309800
rect 519596 309760 539968 309788
rect 519596 309748 519602 309760
rect 539962 309748 539968 309760
rect 540020 309748 540026 309800
rect 535454 309176 535460 309188
rect 532712 309148 535460 309176
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 17310 309108 17316 309120
rect 3384 309080 17316 309108
rect 3384 309068 3390 309080
rect 17310 309068 17316 309080
rect 17368 309068 17374 309120
rect 532326 309068 532332 309120
rect 532384 309108 532390 309120
rect 532712 309108 532740 309148
rect 535454 309136 535460 309148
rect 535512 309136 535518 309188
rect 569954 309136 569960 309188
rect 570012 309176 570018 309188
rect 572714 309176 572720 309188
rect 570012 309148 572720 309176
rect 570012 309136 570018 309148
rect 572714 309136 572720 309148
rect 572772 309136 572778 309188
rect 532384 309080 532740 309108
rect 532384 309068 532390 309080
rect 539686 308660 539692 308712
rect 539744 308700 539750 308712
rect 545114 308700 545120 308712
rect 539744 308672 545120 308700
rect 539744 308660 539750 308672
rect 545114 308660 545120 308672
rect 545172 308660 545178 308712
rect 565078 308388 565084 308440
rect 565136 308428 565142 308440
rect 569954 308428 569960 308440
rect 565136 308400 569960 308428
rect 565136 308388 565142 308400
rect 569954 308388 569960 308400
rect 570012 308388 570018 308440
rect 563054 307816 563060 307828
rect 561692 307788 563060 307816
rect 282822 307708 282828 307760
rect 282880 307748 282886 307760
rect 302878 307748 302884 307760
rect 282880 307720 302884 307748
rect 282880 307708 282886 307720
rect 302878 307708 302884 307720
rect 302936 307708 302942 307760
rect 557534 307708 557540 307760
rect 557592 307748 557598 307760
rect 561692 307748 561720 307788
rect 563054 307776 563060 307788
rect 563112 307776 563118 307828
rect 557592 307720 561720 307748
rect 557592 307708 557598 307720
rect 522482 307096 522488 307148
rect 522540 307136 522546 307148
rect 523494 307136 523500 307148
rect 522540 307108 523500 307136
rect 522540 307096 522546 307108
rect 523494 307096 523500 307108
rect 523552 307096 523558 307148
rect 56502 306348 56508 306400
rect 56560 306388 56566 306400
rect 57514 306388 57520 306400
rect 56560 306360 57520 306388
rect 56560 306348 56566 306360
rect 57514 306348 57520 306360
rect 57572 306348 57578 306400
rect 57606 306348 57612 306400
rect 57664 306388 57670 306400
rect 57974 306388 57980 306400
rect 57664 306360 57980 306388
rect 57664 306348 57670 306360
rect 57974 306348 57980 306360
rect 58032 306348 58038 306400
rect 282086 306280 282092 306332
rect 282144 306320 282150 306332
rect 321554 306320 321560 306332
rect 282144 306292 321560 306320
rect 282144 306280 282150 306292
rect 321554 306280 321560 306292
rect 321612 306280 321618 306332
rect 517514 305600 517520 305652
rect 517572 305640 517578 305652
rect 522482 305640 522488 305652
rect 517572 305612 522488 305640
rect 517572 305600 517578 305612
rect 522482 305600 522488 305612
rect 522540 305600 522546 305652
rect 516134 304988 516140 305040
rect 516192 305028 516198 305040
rect 519538 305028 519544 305040
rect 516192 305000 519544 305028
rect 516192 304988 516198 305000
rect 519538 304988 519544 305000
rect 519596 304988 519602 305040
rect 540974 304988 540980 305040
rect 541032 305028 541038 305040
rect 543090 305028 543096 305040
rect 541032 305000 543096 305028
rect 541032 304988 541038 305000
rect 543090 304988 543096 305000
rect 543148 304988 543154 305040
rect 546494 304988 546500 305040
rect 546552 305028 546558 305040
rect 548518 305028 548524 305040
rect 546552 305000 548524 305028
rect 546552 304988 546558 305000
rect 548518 304988 548524 305000
rect 548576 304988 548582 305040
rect 59262 304444 59268 304496
rect 59320 304484 59326 304496
rect 59446 304484 59452 304496
rect 59320 304456 59452 304484
rect 59320 304444 59326 304456
rect 59446 304444 59452 304456
rect 59504 304444 59510 304496
rect 58710 304308 58716 304360
rect 58768 304348 58774 304360
rect 59538 304348 59544 304360
rect 58768 304320 59544 304348
rect 58768 304308 58774 304320
rect 59538 304308 59544 304320
rect 59596 304308 59602 304360
rect 58802 303424 58808 303476
rect 58860 303464 58866 303476
rect 60642 303464 60648 303476
rect 58860 303436 60648 303464
rect 58860 303424 58866 303436
rect 60642 303424 60648 303436
rect 60700 303424 60706 303476
rect 553394 302744 553400 302796
rect 553452 302784 553458 302796
rect 557534 302784 557540 302796
rect 553452 302756 557540 302784
rect 553452 302744 553458 302756
rect 557534 302744 557540 302756
rect 557592 302744 557598 302796
rect 559098 302336 559104 302388
rect 559156 302376 559162 302388
rect 560938 302376 560944 302388
rect 559156 302348 560944 302376
rect 559156 302336 559162 302348
rect 560938 302336 560944 302348
rect 560996 302336 561002 302388
rect 536834 300976 536840 301028
rect 536892 301016 536898 301028
rect 539686 301016 539692 301028
rect 536892 300988 539692 301016
rect 536892 300976 536898 300988
rect 539686 300976 539692 300988
rect 539744 300976 539750 301028
rect 514754 300840 514760 300892
rect 514812 300880 514818 300892
rect 517514 300880 517520 300892
rect 514812 300852 517520 300880
rect 514812 300840 514818 300852
rect 517514 300840 517520 300852
rect 517572 300840 517578 300892
rect 57882 300772 57888 300824
rect 57940 300812 57946 300824
rect 580258 300812 580264 300824
rect 57940 300784 580264 300812
rect 57940 300772 57946 300784
rect 580258 300772 580264 300784
rect 580316 300772 580322 300824
rect 56686 300704 56692 300756
rect 56744 300744 56750 300756
rect 580350 300744 580356 300756
rect 56744 300716 580356 300744
rect 56744 300704 56750 300716
rect 580350 300704 580356 300716
rect 580408 300704 580414 300756
rect 59446 300636 59452 300688
rect 59504 300676 59510 300688
rect 565078 300676 565084 300688
rect 59504 300648 565084 300676
rect 59504 300636 59510 300648
rect 565078 300636 565084 300648
rect 565136 300636 565142 300688
rect 59998 300568 60004 300620
rect 60056 300608 60062 300620
rect 559098 300608 559104 300620
rect 60056 300580 559104 300608
rect 60056 300568 60062 300580
rect 559098 300568 559104 300580
rect 559156 300568 559162 300620
rect 60642 300500 60648 300552
rect 60700 300540 60706 300552
rect 553394 300540 553400 300552
rect 60700 300512 553400 300540
rect 60700 300500 60706 300512
rect 553394 300500 553400 300512
rect 553452 300500 553458 300552
rect 58618 300432 58624 300484
rect 58676 300472 58682 300484
rect 546494 300472 546500 300484
rect 58676 300444 546500 300472
rect 58676 300432 58682 300444
rect 546494 300432 546500 300444
rect 546552 300432 546558 300484
rect 58434 300364 58440 300416
rect 58492 300404 58498 300416
rect 540882 300404 540888 300416
rect 58492 300376 540888 300404
rect 58492 300364 58498 300376
rect 540882 300364 540888 300376
rect 540940 300364 540946 300416
rect 59538 300296 59544 300348
rect 59596 300336 59602 300348
rect 536834 300336 536840 300348
rect 59596 300308 536840 300336
rect 59596 300296 59602 300308
rect 536834 300296 536840 300308
rect 536892 300296 536898 300348
rect 58986 300228 58992 300280
rect 59044 300268 59050 300280
rect 532326 300268 532332 300280
rect 59044 300240 532332 300268
rect 59044 300228 59050 300240
rect 532326 300228 532332 300240
rect 532384 300228 532390 300280
rect 58894 300160 58900 300212
rect 58952 300200 58958 300212
rect 516134 300200 516140 300212
rect 58952 300172 516140 300200
rect 58952 300160 58958 300172
rect 516134 300160 516140 300172
rect 516192 300160 516198 300212
rect 58526 300092 58532 300144
rect 58584 300132 58590 300144
rect 514754 300132 514760 300144
rect 58584 300104 514760 300132
rect 58584 300092 58590 300104
rect 514754 300092 514760 300104
rect 514812 300092 514818 300144
rect 56778 299412 56784 299464
rect 56836 299452 56842 299464
rect 579798 299452 579804 299464
rect 56836 299424 579804 299452
rect 56836 299412 56842 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 39298 298052 39304 298104
rect 39356 298092 39362 298104
rect 68646 298092 68652 298104
rect 39356 298064 68652 298092
rect 39356 298052 39362 298064
rect 68646 298052 68652 298064
rect 68704 298052 68710 298104
rect 82722 298052 82728 298104
rect 82780 298092 82786 298104
rect 193214 298092 193220 298104
rect 82780 298064 193220 298092
rect 82780 298052 82786 298064
rect 193214 298052 193220 298064
rect 193272 298052 193278 298104
rect 32398 297984 32404 298036
rect 32456 298024 32462 298036
rect 78398 298024 78404 298036
rect 32456 297996 78404 298024
rect 32456 297984 32462 297996
rect 78398 297984 78404 297996
rect 78456 297984 78462 298036
rect 86862 297984 86868 298036
rect 86920 298024 86926 298036
rect 201034 298024 201040 298036
rect 86920 297996 201040 298024
rect 86920 297984 86926 297996
rect 201034 297984 201040 297996
rect 201092 297984 201098 298036
rect 4062 297916 4068 297968
rect 4120 297956 4126 297968
rect 64782 297956 64788 297968
rect 4120 297928 64788 297956
rect 4120 297916 4126 297928
rect 64782 297916 64788 297928
rect 64840 297916 64846 297968
rect 89622 297916 89628 297968
rect 89680 297956 89686 297968
rect 204898 297956 204904 297968
rect 89680 297928 204904 297956
rect 89680 297916 89686 297928
rect 204898 297916 204904 297928
rect 204956 297916 204962 297968
rect 10962 297848 10968 297900
rect 11020 297888 11026 297900
rect 76466 297888 76472 297900
rect 11020 297860 76472 297888
rect 11020 297848 11026 297860
rect 76466 297848 76472 297860
rect 76524 297848 76530 297900
rect 96522 297848 96528 297900
rect 96580 297888 96586 297900
rect 216582 297888 216588 297900
rect 96580 297860 216588 297888
rect 96580 297848 96586 297860
rect 216582 297848 216588 297860
rect 216640 297848 216646 297900
rect 16482 297780 16488 297832
rect 16540 297820 16546 297832
rect 86218 297820 86224 297832
rect 16540 297792 86224 297820
rect 16540 297780 16546 297792
rect 86218 297780 86224 297792
rect 86276 297780 86282 297832
rect 93762 297780 93768 297832
rect 93820 297820 93826 297832
rect 212718 297820 212724 297832
rect 93820 297792 212724 297820
rect 93820 297780 93826 297792
rect 212718 297780 212724 297792
rect 212776 297780 212782 297832
rect 42702 297712 42708 297764
rect 42760 297752 42766 297764
rect 128998 297752 129004 297764
rect 42760 297724 129004 297752
rect 42760 297712 42766 297724
rect 128998 297712 129004 297724
rect 129056 297712 129062 297764
rect 134518 297712 134524 297764
rect 134576 297752 134582 297764
rect 255498 297752 255504 297764
rect 134576 297724 255504 297752
rect 134576 297712 134582 297724
rect 255498 297712 255504 297724
rect 255556 297712 255562 297764
rect 15102 297644 15108 297696
rect 15160 297684 15166 297696
rect 84194 297684 84200 297696
rect 15160 297656 84200 297684
rect 15160 297644 15166 297656
rect 84194 297644 84200 297656
rect 84252 297644 84258 297696
rect 100662 297644 100668 297696
rect 100720 297684 100726 297696
rect 224402 297684 224408 297696
rect 100720 297656 224408 297684
rect 100720 297644 100726 297656
rect 224402 297644 224408 297656
rect 224460 297644 224466 297696
rect 20622 297576 20628 297628
rect 20680 297616 20686 297628
rect 92014 297616 92020 297628
rect 20680 297588 92020 297616
rect 20680 297576 20686 297588
rect 92014 297576 92020 297588
rect 92072 297576 92078 297628
rect 103422 297576 103428 297628
rect 103480 297616 103486 297628
rect 228266 297616 228272 297628
rect 103480 297588 228272 297616
rect 103480 297576 103486 297588
rect 228266 297576 228272 297588
rect 228324 297576 228330 297628
rect 21910 297508 21916 297560
rect 21968 297548 21974 297560
rect 93946 297548 93952 297560
rect 21968 297520 93952 297548
rect 21968 297508 21974 297520
rect 93946 297508 93952 297520
rect 94004 297508 94010 297560
rect 107562 297508 107568 297560
rect 107620 297548 107626 297560
rect 234154 297548 234160 297560
rect 107620 297520 234160 297548
rect 107620 297508 107626 297520
rect 234154 297508 234160 297520
rect 234212 297508 234218 297560
rect 24762 297440 24768 297492
rect 24820 297480 24826 297492
rect 99834 297480 99840 297492
rect 24820 297452 99840 297480
rect 24820 297440 24826 297452
rect 99834 297440 99840 297452
rect 99892 297440 99898 297492
rect 107470 297440 107476 297492
rect 107528 297480 107534 297492
rect 236086 297480 236092 297492
rect 107528 297452 236092 297480
rect 107528 297440 107534 297452
rect 236086 297440 236092 297452
rect 236144 297440 236150 297492
rect 26142 297372 26148 297424
rect 26200 297412 26206 297424
rect 101766 297412 101772 297424
rect 26200 297384 101772 297412
rect 26200 297372 26206 297384
rect 101766 297372 101772 297384
rect 101824 297372 101830 297424
rect 114462 297372 114468 297424
rect 114520 297412 114526 297424
rect 245838 297412 245844 297424
rect 114520 297384 245844 297412
rect 114520 297372 114526 297384
rect 245838 297372 245844 297384
rect 245896 297372 245902 297424
rect 51810 297304 51816 297356
rect 51868 297344 51874 297356
rect 70578 297344 70584 297356
rect 51868 297316 70584 297344
rect 51868 297304 51874 297316
rect 70578 297304 70584 297316
rect 70636 297304 70642 297356
rect 79962 297304 79968 297356
rect 80020 297344 80026 297356
rect 189350 297344 189356 297356
rect 80020 297316 189356 297344
rect 80020 297304 80026 297316
rect 189350 297304 189356 297316
rect 189408 297304 189414 297356
rect 74442 297236 74448 297288
rect 74500 297276 74506 297288
rect 181530 297276 181536 297288
rect 74500 297248 181536 297276
rect 74500 297236 74506 297248
rect 181530 297236 181536 297248
rect 181588 297236 181594 297288
rect 72970 297168 72976 297220
rect 73028 297208 73034 297220
rect 177666 297208 177672 297220
rect 73028 297180 177672 297208
rect 73028 297168 73034 297180
rect 177666 297168 177672 297180
rect 177724 297168 177730 297220
rect 67542 297100 67548 297152
rect 67600 297140 67606 297152
rect 169846 297140 169852 297152
rect 67600 297112 169852 297140
rect 67600 297100 67606 297112
rect 169846 297100 169852 297112
rect 169904 297100 169910 297152
rect 64782 297032 64788 297084
rect 64840 297072 64846 297084
rect 165982 297072 165988 297084
rect 64840 297044 165988 297072
rect 64840 297032 64846 297044
rect 165982 297032 165988 297044
rect 166040 297032 166046 297084
rect 62022 296964 62028 297016
rect 62080 297004 62086 297016
rect 160186 297004 160192 297016
rect 62080 296976 160192 297004
rect 62080 296964 62086 296976
rect 160186 296964 160192 296976
rect 160244 296964 160250 297016
rect 50982 296896 50988 296948
rect 51040 296936 51046 296948
rect 142614 296936 142620 296948
rect 51040 296908 142620 296936
rect 51040 296896 51046 296908
rect 142614 296896 142620 296908
rect 142672 296896 142678 296948
rect 48130 296828 48136 296880
rect 48188 296868 48194 296880
rect 136818 296868 136824 296880
rect 48188 296840 136824 296868
rect 48188 296828 48194 296840
rect 136818 296828 136824 296840
rect 136876 296828 136882 296880
rect 39942 296760 39948 296812
rect 40000 296800 40006 296812
rect 124766 296800 124772 296812
rect 40000 296772 124772 296800
rect 40000 296760 40006 296772
rect 124766 296760 124772 296772
rect 124824 296760 124830 296812
rect 124858 296760 124864 296812
rect 124916 296800 124922 296812
rect 146570 296800 146576 296812
rect 124916 296772 146576 296800
rect 124916 296760 124922 296772
rect 146570 296760 146576 296772
rect 146628 296760 146634 296812
rect 42058 296692 42064 296744
rect 42116 296732 42122 296744
rect 107286 296732 107292 296744
rect 42116 296704 107292 296732
rect 42116 296692 42122 296704
rect 107286 296692 107292 296704
rect 107344 296692 107350 296744
rect 56686 296624 56692 296676
rect 56744 296664 56750 296676
rect 57330 296664 57336 296676
rect 56744 296636 57336 296664
rect 56744 296624 56750 296636
rect 57330 296624 57336 296636
rect 57388 296624 57394 296676
rect 57514 296624 57520 296676
rect 57572 296664 57578 296676
rect 57882 296664 57888 296676
rect 57572 296636 57888 296664
rect 57572 296624 57578 296636
rect 57882 296624 57888 296636
rect 57940 296624 57946 296676
rect 2958 295264 2964 295316
rect 3016 295304 3022 295316
rect 57238 295304 57244 295316
rect 3016 295276 57244 295304
rect 3016 295264 3022 295276
rect 57238 295264 57244 295276
rect 57296 295264 57302 295316
rect 61010 292544 61016 292596
rect 61068 292544 61074 292596
rect 61028 292516 61056 292544
rect 61102 292516 61108 292528
rect 61028 292488 61108 292516
rect 61102 292476 61108 292488
rect 61160 292476 61166 292528
rect 61010 288396 61016 288448
rect 61068 288436 61074 288448
rect 61102 288436 61108 288448
rect 61068 288408 61108 288436
rect 61068 288396 61074 288408
rect 61102 288396 61108 288408
rect 61160 288396 61166 288448
rect 56778 287104 56784 287156
rect 56836 287144 56842 287156
rect 57606 287144 57612 287156
rect 56836 287116 57612 287144
rect 56836 287104 56842 287116
rect 57606 287104 57612 287116
rect 57664 287104 57670 287156
rect 56686 287036 56692 287088
rect 56744 287076 56750 287088
rect 57330 287076 57336 287088
rect 56744 287048 57336 287076
rect 56744 287036 56750 287048
rect 57330 287036 57336 287048
rect 57388 287036 57394 287088
rect 57514 287036 57520 287088
rect 57572 287076 57578 287088
rect 57882 287076 57888 287088
rect 57572 287048 57888 287076
rect 57572 287036 57578 287048
rect 57882 287036 57888 287048
rect 57940 287036 57946 287088
rect 67542 280372 67548 280424
rect 67600 280372 67606 280424
rect 67560 280288 67588 280372
rect 67542 280236 67548 280288
rect 67600 280236 67606 280288
rect 3326 280100 3332 280152
rect 3384 280140 3390 280152
rect 37918 280140 37924 280152
rect 3384 280112 37924 280140
rect 3384 280100 3390 280112
rect 37918 280100 37924 280112
rect 37976 280100 37982 280152
rect 57238 277312 57244 277364
rect 57296 277352 57302 277364
rect 57514 277352 57520 277364
rect 57296 277324 57520 277352
rect 57296 277312 57302 277324
rect 57514 277312 57520 277324
rect 57572 277312 57578 277364
rect 57606 277312 57612 277364
rect 57664 277352 57670 277364
rect 57882 277352 57888 277364
rect 57664 277324 57888 277352
rect 57664 277312 57670 277324
rect 57882 277312 57888 277324
rect 57940 277312 57946 277364
rect 56870 275952 56876 276004
rect 56928 275992 56934 276004
rect 580166 275992 580172 276004
rect 56928 275964 580172 275992
rect 56928 275952 56934 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 60734 273232 60740 273284
rect 60792 273272 60798 273284
rect 61102 273272 61108 273284
rect 60792 273244 61108 273272
rect 60792 273232 60798 273244
rect 61102 273232 61108 273244
rect 61160 273232 61166 273284
rect 56778 268404 56784 268456
rect 56836 268444 56842 268456
rect 57330 268444 57336 268456
rect 56836 268416 57336 268444
rect 56836 268404 56842 268416
rect 57330 268404 57336 268416
rect 57388 268404 57394 268456
rect 57606 268404 57612 268456
rect 57664 268444 57670 268456
rect 57882 268444 57888 268456
rect 57664 268416 57888 268444
rect 57664 268404 57670 268416
rect 57882 268404 57888 268416
rect 57940 268404 57946 268456
rect 3142 266296 3148 266348
rect 3200 266336 3206 266348
rect 20070 266336 20076 266348
rect 3200 266308 20076 266336
rect 3200 266296 3206 266308
rect 20070 266296 20076 266308
rect 20128 266296 20134 266348
rect 56962 264868 56968 264920
rect 57020 264908 57026 264920
rect 580166 264908 580172 264920
rect 57020 264880 580172 264908
rect 57020 264868 57026 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 57238 263576 57244 263628
rect 57296 263616 57302 263628
rect 57514 263616 57520 263628
rect 57296 263588 57520 263616
rect 57296 263576 57302 263588
rect 57514 263576 57520 263588
rect 57572 263576 57578 263628
rect 60918 263508 60924 263560
rect 60976 263548 60982 263560
rect 61102 263548 61108 263560
rect 60976 263520 61108 263548
rect 60976 263508 60982 263520
rect 61102 263508 61108 263520
rect 61160 263508 61166 263560
rect 60826 260788 60832 260840
rect 60884 260828 60890 260840
rect 61102 260828 61108 260840
rect 60884 260800 61108 260828
rect 60884 260788 60890 260800
rect 61102 260788 61108 260800
rect 61160 260788 61166 260840
rect 57054 252492 57060 252544
rect 57112 252532 57118 252544
rect 579798 252532 579804 252544
rect 57112 252504 579804 252532
rect 57112 252492 57118 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 60826 251200 60832 251252
rect 60884 251240 60890 251252
rect 61010 251240 61016 251252
rect 60884 251212 61016 251240
rect 60884 251200 60890 251212
rect 61010 251200 61016 251212
rect 61068 251200 61074 251252
rect 3234 237328 3240 237380
rect 3292 237368 3298 237380
rect 39390 237368 39396 237380
rect 3292 237340 39396 237368
rect 3292 237328 3298 237340
rect 39390 237328 39396 237340
rect 39448 237328 39454 237380
rect 67358 231820 67364 231872
rect 67416 231820 67422 231872
rect 67376 231736 67404 231820
rect 67358 231684 67364 231736
rect 67416 231684 67422 231736
rect 67266 230392 67272 230444
rect 67324 230432 67330 230444
rect 67358 230432 67364 230444
rect 67324 230404 67364 230432
rect 67324 230392 67330 230404
rect 67358 230392 67364 230404
rect 67416 230392 67422 230444
rect 57146 229032 57152 229084
rect 57204 229072 57210 229084
rect 580166 229072 580172 229084
rect 57204 229044 580172 229072
rect 57204 229032 57210 229044
rect 580166 229032 580172 229044
rect 580224 229032 580230 229084
rect 60734 224952 60740 225004
rect 60792 224952 60798 225004
rect 60752 224856 60780 224952
rect 60918 224856 60924 224868
rect 60752 224828 60924 224856
rect 60918 224816 60924 224828
rect 60976 224816 60982 224868
rect 3326 223524 3332 223576
rect 3384 223564 3390 223576
rect 28258 223564 28264 223576
rect 3384 223536 28264 223564
rect 3384 223524 3390 223536
rect 28258 223524 28264 223536
rect 28316 223524 28322 223576
rect 67266 220804 67272 220856
rect 67324 220844 67330 220856
rect 67542 220844 67548 220856
rect 67324 220816 67548 220844
rect 67324 220804 67330 220816
rect 67542 220804 67548 220816
rect 67600 220804 67606 220856
rect 57330 217948 57336 218000
rect 57388 217988 57394 218000
rect 580166 217988 580172 218000
rect 57388 217960 580172 217988
rect 57388 217948 57394 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 60734 215296 60740 215348
rect 60792 215336 60798 215348
rect 60918 215336 60924 215348
rect 60792 215308 60924 215336
rect 60792 215296 60798 215308
rect 60918 215296 60924 215308
rect 60976 215296 60982 215348
rect 67542 212548 67548 212560
rect 67468 212520 67548 212548
rect 67468 212492 67496 212520
rect 67542 212508 67548 212520
rect 67600 212508 67606 212560
rect 67450 212440 67456 212492
rect 67508 212440 67514 212492
rect 67450 211080 67456 211132
rect 67508 211120 67514 211132
rect 67542 211120 67548 211132
rect 67508 211092 67548 211120
rect 67508 211080 67514 211092
rect 67542 211080 67548 211092
rect 67600 211080 67606 211132
rect 57422 205572 57428 205624
rect 57480 205612 57486 205624
rect 579798 205612 579804 205624
rect 57480 205584 579804 205612
rect 57480 205572 57486 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 60642 205504 60648 205556
rect 60700 205544 60706 205556
rect 60918 205544 60924 205556
rect 60700 205516 60924 205544
rect 60700 205504 60706 205516
rect 60918 205504 60924 205516
rect 60976 205504 60982 205556
rect 67542 202852 67548 202904
rect 67600 202852 67606 202904
rect 67450 202784 67456 202836
rect 67508 202824 67514 202836
rect 67560 202824 67588 202852
rect 67508 202796 67588 202824
rect 67508 202784 67514 202796
rect 60918 195984 60924 196036
rect 60976 195984 60982 196036
rect 60936 195956 60964 195984
rect 61010 195956 61016 195968
rect 60936 195928 61016 195956
rect 61010 195916 61016 195928
rect 61068 195916 61074 195968
rect 3510 194488 3516 194540
rect 3568 194528 3574 194540
rect 50338 194528 50344 194540
rect 3568 194500 50344 194528
rect 3568 194488 3574 194500
rect 50338 194488 50344 194500
rect 50396 194488 50402 194540
rect 57514 182112 57520 182164
rect 57572 182152 57578 182164
rect 580166 182152 580172 182164
rect 57572 182124 580172 182152
rect 57572 182112 57578 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 60918 181500 60924 181552
rect 60976 181540 60982 181552
rect 61102 181540 61108 181552
rect 60976 181512 61108 181540
rect 60976 181500 60982 181512
rect 61102 181500 61108 181512
rect 61160 181500 61166 181552
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 33778 180792 33784 180804
rect 3292 180764 33784 180792
rect 3292 180752 3298 180764
rect 33778 180752 33784 180764
rect 33836 180752 33842 180804
rect 57606 171028 57612 171080
rect 57664 171068 57670 171080
rect 580166 171068 580172 171080
rect 57664 171040 580172 171068
rect 57664 171028 57670 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 60918 166948 60924 167000
rect 60976 166988 60982 167000
rect 61102 166988 61108 167000
rect 60976 166960 61108 166988
rect 60976 166948 60982 166960
rect 61102 166948 61108 166960
rect 61160 166948 61166 167000
rect 59354 158652 59360 158704
rect 59412 158692 59418 158704
rect 579798 158692 579804 158704
rect 59412 158664 579804 158692
rect 59412 158652 59418 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 61194 157468 61200 157480
rect 61028 157440 61200 157468
rect 61028 157276 61056 157440
rect 61194 157428 61200 157440
rect 61252 157428 61258 157480
rect 61010 157224 61016 157276
rect 61068 157224 61074 157276
rect 61010 153144 61016 153196
rect 61068 153184 61074 153196
rect 61194 153184 61200 153196
rect 61068 153156 61200 153184
rect 61068 153144 61074 153156
rect 61194 153144 61200 153156
rect 61252 153144 61258 153196
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 51718 151756 51724 151768
rect 3200 151728 51724 151756
rect 3200 151716 3206 151728
rect 51718 151716 51724 151728
rect 51776 151716 51782 151768
rect 60918 137980 60924 138032
rect 60976 137980 60982 138032
rect 60936 137952 60964 137980
rect 61010 137952 61016 137964
rect 60936 137924 61016 137952
rect 61010 137912 61016 137924
rect 61068 137912 61074 137964
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 35158 136592 35164 136604
rect 3292 136564 35164 136592
rect 3292 136552 3298 136564
rect 35158 136552 35164 136564
rect 35216 136552 35222 136604
rect 57698 135192 57704 135244
rect 57756 135232 57762 135244
rect 580166 135232 580172 135244
rect 57756 135204 580172 135232
rect 57756 135192 57762 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 57790 124108 57796 124160
rect 57848 124148 57854 124160
rect 580166 124148 580172 124160
rect 57848 124120 580172 124148
rect 57848 124108 57854 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 2774 122272 2780 122324
rect 2832 122312 2838 122324
rect 4982 122312 4988 122324
rect 2832 122284 4988 122312
rect 2832 122272 2838 122284
rect 4982 122272 4988 122284
rect 5040 122272 5046 122324
rect 60918 118668 60924 118720
rect 60976 118668 60982 118720
rect 60936 118640 60964 118668
rect 61010 118640 61016 118652
rect 60936 118612 61016 118640
rect 61010 118600 61016 118612
rect 61068 118600 61074 118652
rect 67450 115880 67456 115932
rect 67508 115920 67514 115932
rect 67542 115920 67548 115932
rect 67508 115892 67548 115920
rect 67508 115880 67514 115892
rect 67542 115880 67548 115892
rect 67600 115880 67606 115932
rect 67266 114452 67272 114504
rect 67324 114492 67330 114504
rect 67450 114492 67456 114504
rect 67324 114464 67456 114492
rect 67324 114452 67330 114464
rect 67450 114452 67456 114464
rect 67508 114452 67514 114504
rect 59078 111732 59084 111784
rect 59136 111772 59142 111784
rect 579798 111772 579804 111784
rect 59136 111744 579804 111772
rect 59136 111732 59142 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 17218 108984 17224 108996
rect 3292 108956 17224 108984
rect 3292 108944 3298 108956
rect 17218 108944 17224 108956
rect 17276 108944 17282 108996
rect 67266 104864 67272 104916
rect 67324 104904 67330 104916
rect 67542 104904 67548 104916
rect 67324 104876 67548 104904
rect 67324 104864 67330 104876
rect 67542 104864 67548 104876
rect 67600 104864 67606 104916
rect 60734 99356 60740 99408
rect 60792 99356 60798 99408
rect 60752 99260 60780 99356
rect 61102 99260 61108 99272
rect 60752 99232 61108 99260
rect 61102 99220 61108 99232
rect 61160 99220 61166 99272
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 43438 93820 43444 93832
rect 3476 93792 43444 93820
rect 3476 93780 3482 93792
rect 43438 93780 43444 93792
rect 43496 93780 43502 93832
rect 56594 88272 56600 88324
rect 56652 88312 56658 88324
rect 580166 88312 580172 88324
rect 56652 88284 580172 88312
rect 56652 88272 56658 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 60734 86912 60740 86964
rect 60792 86952 60798 86964
rect 61010 86952 61016 86964
rect 60792 86924 61016 86952
rect 60792 86912 60798 86924
rect 61010 86912 61016 86924
rect 61068 86912 61074 86964
rect 2774 79772 2780 79824
rect 2832 79812 2838 79824
rect 4890 79812 4896 79824
rect 2832 79784 4896 79812
rect 2832 79772 2838 79784
rect 4890 79772 4896 79784
rect 4948 79772 4954 79824
rect 60734 77256 60740 77308
rect 60792 77296 60798 77308
rect 60918 77296 60924 77308
rect 60792 77268 60924 77296
rect 60792 77256 60798 77268
rect 60918 77256 60924 77268
rect 60976 77256 60982 77308
rect 89530 76100 89536 76152
rect 89588 76140 89594 76152
rect 89806 76140 89812 76152
rect 89588 76112 89812 76140
rect 89588 76100 89594 76112
rect 89806 76100 89812 76112
rect 89864 76100 89870 76152
rect 147582 76100 147588 76152
rect 147640 76140 147646 76152
rect 154482 76140 154488 76152
rect 147640 76112 154488 76140
rect 147640 76100 147646 76112
rect 154482 76100 154488 76112
rect 154540 76100 154546 76152
rect 115934 75964 115940 76016
rect 115992 76004 115998 76016
rect 118878 76004 118884 76016
rect 115992 75976 118884 76004
rect 115992 75964 115998 75976
rect 118878 75964 118884 75976
rect 118936 75964 118942 76016
rect 60642 75828 60648 75880
rect 60700 75868 60706 75880
rect 60918 75868 60924 75880
rect 60700 75840 60924 75868
rect 60700 75828 60706 75840
rect 60918 75828 60924 75840
rect 60976 75828 60982 75880
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 53098 64852 53104 64864
rect 3384 64824 53104 64852
rect 3384 64812 3390 64824
rect 53098 64812 53104 64824
rect 53156 64812 53162 64864
rect 59170 64812 59176 64864
rect 59228 64852 59234 64864
rect 579798 64852 579804 64864
rect 59228 64824 579804 64852
rect 59228 64812 59234 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 60918 60664 60924 60716
rect 60976 60704 60982 60716
rect 61102 60704 61108 60716
rect 60976 60676 61108 60704
rect 60976 60664 60982 60676
rect 61102 60664 61108 60676
rect 61160 60664 61166 60716
rect 60826 57876 60832 57928
rect 60884 57916 60890 57928
rect 61102 57916 61108 57928
rect 60884 57888 61108 57916
rect 60884 57876 60890 57888
rect 61102 57876 61108 57888
rect 61160 57876 61166 57928
rect 67450 57876 67456 57928
rect 67508 57916 67514 57928
rect 67542 57916 67548 57928
rect 67508 57888 67548 57916
rect 67508 57876 67514 57888
rect 67542 57876 67548 57888
rect 67600 57876 67606 57928
rect 67266 56516 67272 56568
rect 67324 56556 67330 56568
rect 67450 56556 67456 56568
rect 67324 56528 67456 56556
rect 67324 56516 67330 56528
rect 67450 56516 67456 56528
rect 67508 56516 67514 56568
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 46198 51048 46204 51060
rect 3476 51020 46204 51048
rect 3476 51008 3482 51020
rect 46198 51008 46204 51020
rect 46256 51008 46262 51060
rect 60826 48288 60832 48340
rect 60884 48328 60890 48340
rect 61010 48328 61016 48340
rect 60884 48300 61016 48328
rect 60884 48288 60890 48300
rect 61010 48288 61016 48300
rect 61068 48288 61074 48340
rect 67266 46928 67272 46980
rect 67324 46968 67330 46980
rect 67542 46968 67548 46980
rect 67324 46940 67548 46968
rect 67324 46928 67330 46940
rect 67542 46928 67548 46940
rect 67600 46928 67606 46980
rect 147582 40196 147588 40248
rect 147640 40236 147646 40248
rect 154482 40236 154488 40248
rect 147640 40208 154488 40236
rect 147640 40196 147646 40208
rect 154482 40196 154488 40208
rect 154540 40196 154546 40248
rect 89530 40128 89536 40180
rect 89588 40168 89594 40180
rect 91738 40168 91744 40180
rect 89588 40140 91744 40168
rect 89588 40128 89594 40140
rect 91738 40128 91744 40140
rect 91796 40128 91802 40180
rect 115934 40060 115940 40112
rect 115992 40100 115998 40112
rect 118878 40100 118884 40112
rect 115992 40072 118884 40100
rect 115992 40060 115998 40072
rect 118878 40060 118884 40072
rect 118936 40060 118942 40112
rect 67450 37272 67456 37324
rect 67508 37312 67514 37324
rect 67542 37312 67548 37324
rect 67508 37284 67548 37312
rect 67508 37272 67514 37284
rect 67542 37272 67548 37284
rect 67600 37272 67606 37324
rect 2774 35844 2780 35896
rect 2832 35884 2838 35896
rect 4798 35884 4804 35896
rect 2832 35856 4804 35884
rect 2832 35844 2838 35856
rect 4798 35844 4804 35856
rect 4856 35844 4862 35896
rect 60918 31832 60924 31884
rect 60976 31832 60982 31884
rect 60936 31748 60964 31832
rect 60918 31696 60924 31748
rect 60976 31696 60982 31748
rect 86862 29248 86868 29300
rect 86920 29248 86926 29300
rect 86880 29164 86908 29248
rect 147582 29180 147588 29232
rect 147640 29220 147646 29232
rect 154482 29220 154488 29232
rect 147640 29192 154488 29220
rect 147640 29180 147646 29192
rect 154482 29180 154488 29192
rect 154540 29180 154546 29232
rect 86862 29112 86868 29164
rect 86920 29112 86926 29164
rect 115934 29044 115940 29096
rect 115992 29084 115998 29096
rect 120810 29084 120816 29096
rect 115992 29056 120816 29084
rect 115992 29044 115998 29056
rect 120810 29044 120816 29056
rect 120868 29044 120874 29096
rect 67542 27616 67548 27668
rect 67600 27656 67606 27668
rect 67726 27656 67732 27668
rect 67600 27628 67732 27656
rect 67600 27616 67606 27628
rect 67726 27616 67732 27628
rect 67784 27616 67790 27668
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 19978 22080 19984 22092
rect 2924 22052 19984 22080
rect 2924 22040 2930 22052
rect 19978 22040 19984 22052
rect 20036 22040 20042 22092
rect 67542 19252 67548 19304
rect 67600 19252 67606 19304
rect 66990 19184 66996 19236
rect 67048 19224 67054 19236
rect 67560 19224 67588 19252
rect 67048 19196 67588 19224
rect 67048 19184 67054 19196
rect 59262 17892 59268 17944
rect 59320 17932 59326 17944
rect 579798 17932 579804 17944
rect 59320 17904 579804 17932
rect 59320 17892 59326 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 60734 12452 60740 12504
rect 60792 12452 60798 12504
rect 60752 12356 60780 12452
rect 60826 12356 60832 12368
rect 60752 12328 60832 12356
rect 60826 12316 60832 12328
rect 60884 12316 60890 12368
rect 59170 9596 59176 9648
rect 59228 9636 59234 9648
rect 60826 9636 60832 9648
rect 59228 9608 60832 9636
rect 59228 9596 59234 9608
rect 60826 9596 60832 9608
rect 60884 9596 60890 9648
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 48958 8276 48964 8288
rect 3476 8248 48964 8276
rect 3476 8236 3482 8248
rect 48958 8236 48964 8248
rect 49016 8236 49022 8288
rect 59998 6400 60004 6452
rect 60056 6440 60062 6452
rect 157334 6440 157340 6452
rect 60056 6412 157340 6440
rect 60056 6400 60062 6412
rect 157334 6400 157340 6412
rect 157392 6400 157398 6452
rect 108758 6332 108764 6384
rect 108816 6372 108822 6384
rect 237374 6372 237380 6384
rect 108816 6344 237380 6372
rect 108816 6332 108822 6344
rect 237374 6332 237380 6344
rect 237432 6332 237438 6384
rect 112346 6264 112352 6316
rect 112404 6304 112410 6316
rect 242894 6304 242900 6316
rect 112404 6276 242900 6304
rect 112404 6264 112410 6276
rect 242894 6264 242900 6276
rect 242952 6264 242958 6316
rect 115934 6196 115940 6248
rect 115992 6236 115998 6248
rect 248414 6236 248420 6248
rect 115992 6208 248420 6236
rect 115992 6196 115998 6208
rect 248414 6196 248420 6208
rect 248472 6196 248478 6248
rect 123018 6128 123024 6180
rect 123076 6168 123082 6180
rect 260834 6168 260840 6180
rect 123076 6140 260840 6168
rect 123076 6128 123082 6140
rect 260834 6128 260840 6140
rect 260892 6128 260898 6180
rect 93854 5516 93860 5568
rect 93912 5556 93918 5568
rect 99466 5556 99472 5568
rect 93912 5528 99472 5556
rect 93912 5516 93918 5528
rect 99466 5516 99472 5528
rect 99524 5516 99530 5568
rect 108942 5516 108948 5568
rect 109000 5556 109006 5568
rect 109034 5556 109040 5568
rect 109000 5528 109040 5556
rect 109000 5516 109006 5528
rect 109034 5516 109040 5528
rect 109092 5516 109098 5568
rect 7650 5448 7656 5500
rect 7708 5488 7714 5500
rect 71774 5488 71780 5500
rect 7708 5460 71780 5488
rect 7708 5448 7714 5460
rect 71774 5448 71780 5460
rect 71832 5448 71838 5500
rect 71866 5448 71872 5500
rect 71924 5488 71930 5500
rect 71924 5460 80192 5488
rect 71924 5448 71930 5460
rect 12434 5380 12440 5432
rect 12492 5420 12498 5432
rect 80054 5420 80060 5432
rect 12492 5392 80060 5420
rect 12492 5380 12498 5392
rect 80054 5380 80060 5392
rect 80112 5380 80118 5432
rect 80164 5420 80192 5460
rect 80238 5448 80244 5500
rect 80296 5488 80302 5500
rect 190454 5488 190460 5500
rect 80296 5460 190460 5488
rect 80296 5448 80302 5460
rect 190454 5448 190460 5460
rect 190512 5448 190518 5500
rect 83734 5420 83740 5432
rect 80164 5392 83740 5420
rect 83734 5380 83740 5392
rect 83792 5380 83798 5432
rect 83826 5380 83832 5432
rect 83884 5420 83890 5432
rect 195974 5420 195980 5432
rect 83884 5392 195980 5420
rect 83884 5380 83890 5392
rect 195974 5380 195980 5392
rect 196032 5380 196038 5432
rect 17218 5312 17224 5364
rect 17276 5352 17282 5364
rect 86954 5352 86960 5364
rect 17276 5324 86960 5352
rect 17276 5312 17282 5324
rect 86954 5312 86960 5324
rect 87012 5312 87018 5364
rect 87322 5312 87328 5364
rect 87380 5352 87386 5364
rect 202874 5352 202880 5364
rect 87380 5324 202880 5352
rect 87380 5312 87386 5324
rect 202874 5312 202880 5324
rect 202932 5312 202938 5364
rect 65518 5244 65524 5296
rect 65576 5284 65582 5296
rect 71866 5284 71872 5296
rect 65576 5256 71872 5284
rect 65576 5244 65582 5256
rect 71866 5244 71872 5256
rect 71924 5244 71930 5296
rect 84102 5244 84108 5296
rect 84160 5284 84166 5296
rect 93854 5284 93860 5296
rect 84160 5256 93860 5284
rect 84160 5244 84166 5256
rect 93854 5244 93860 5256
rect 93912 5244 93918 5296
rect 108942 5284 108948 5296
rect 99392 5256 108948 5284
rect 22002 5176 22008 5228
rect 22060 5216 22066 5228
rect 95234 5216 95240 5228
rect 22060 5188 95240 5216
rect 22060 5176 22066 5188
rect 95234 5176 95240 5188
rect 95292 5176 95298 5228
rect 98086 5176 98092 5228
rect 98144 5216 98150 5228
rect 99392 5216 99420 5256
rect 108942 5244 108948 5256
rect 109000 5244 109006 5296
rect 109034 5244 109040 5296
rect 109092 5284 109098 5296
rect 219434 5284 219440 5296
rect 109092 5256 219440 5284
rect 109092 5244 109098 5256
rect 219434 5244 219440 5256
rect 219492 5244 219498 5296
rect 98144 5188 99420 5216
rect 98144 5176 98150 5188
rect 99466 5176 99472 5228
rect 99524 5216 99530 5228
rect 99524 5188 104112 5216
rect 99524 5176 99530 5188
rect 26694 5108 26700 5160
rect 26752 5148 26758 5160
rect 103514 5148 103520 5160
rect 26752 5120 103520 5148
rect 26752 5108 26758 5120
rect 103514 5108 103520 5120
rect 103572 5108 103578 5160
rect 104084 5148 104112 5188
rect 105170 5176 105176 5228
rect 105228 5216 105234 5228
rect 231854 5216 231860 5228
rect 105228 5188 231860 5216
rect 105228 5176 105234 5188
rect 231854 5176 231860 5188
rect 231912 5176 231918 5228
rect 124858 5148 124864 5160
rect 104084 5120 124864 5148
rect 124858 5108 124864 5120
rect 124916 5108 124922 5160
rect 127802 5108 127808 5160
rect 127860 5148 127866 5160
rect 137370 5148 137376 5160
rect 127860 5120 137376 5148
rect 127860 5108 127866 5120
rect 137370 5108 137376 5120
rect 137428 5108 137434 5160
rect 137646 5108 137652 5160
rect 137704 5148 137710 5160
rect 266354 5148 266360 5160
rect 137704 5120 266360 5148
rect 137704 5108 137710 5120
rect 266354 5108 266360 5120
rect 266412 5108 266418 5160
rect 30282 5040 30288 5092
rect 30340 5080 30346 5092
rect 109126 5080 109132 5092
rect 30340 5052 109132 5080
rect 30340 5040 30346 5052
rect 109126 5040 109132 5052
rect 109184 5040 109190 5092
rect 119430 5040 119436 5092
rect 119488 5080 119494 5092
rect 134518 5080 134524 5092
rect 119488 5052 134524 5080
rect 119488 5040 119494 5052
rect 134518 5040 134524 5052
rect 134576 5040 134582 5092
rect 134610 5040 134616 5092
rect 134668 5080 134674 5092
rect 137186 5080 137192 5092
rect 134668 5052 137192 5080
rect 134668 5040 134674 5052
rect 137186 5040 137192 5052
rect 137244 5040 137250 5092
rect 271874 5080 271880 5092
rect 137296 5052 271880 5080
rect 33870 4972 33876 5024
rect 33928 5012 33934 5024
rect 114554 5012 114560 5024
rect 33928 4984 114560 5012
rect 33928 4972 33934 4984
rect 114554 4972 114560 4984
rect 114612 4972 114618 5024
rect 130194 4972 130200 5024
rect 130252 5012 130258 5024
rect 137296 5012 137324 5052
rect 271874 5040 271880 5052
rect 271932 5040 271938 5092
rect 130252 4984 137324 5012
rect 130252 4972 130258 4984
rect 137462 4972 137468 5024
rect 137520 5012 137526 5024
rect 269114 5012 269120 5024
rect 137520 4984 269120 5012
rect 137520 4972 137526 4984
rect 269114 4972 269120 4984
rect 269172 4972 269178 5024
rect 37366 4904 37372 4956
rect 37424 4944 37430 4956
rect 120074 4944 120080 4956
rect 37424 4916 120080 4944
rect 37424 4904 37430 4916
rect 120074 4904 120080 4916
rect 120132 4904 120138 4956
rect 126606 4904 126612 4956
rect 126664 4944 126670 4956
rect 126664 4916 127480 4944
rect 126664 4904 126670 4916
rect 40954 4836 40960 4888
rect 41012 4876 41018 4888
rect 126974 4876 126980 4888
rect 41012 4848 126980 4876
rect 41012 4836 41018 4848
rect 126974 4836 126980 4848
rect 127032 4836 127038 4888
rect 127452 4876 127480 4916
rect 128998 4904 129004 4956
rect 129056 4944 129062 4956
rect 270494 4944 270500 4956
rect 129056 4916 270500 4944
rect 129056 4904 129062 4916
rect 270494 4904 270500 4916
rect 270552 4904 270558 4956
rect 137462 4876 137468 4888
rect 127452 4848 137468 4876
rect 137462 4836 137468 4848
rect 137520 4836 137526 4888
rect 137554 4836 137560 4888
rect 137612 4876 137618 4888
rect 276014 4876 276020 4888
rect 137612 4848 276020 4876
rect 137612 4836 137618 4848
rect 276014 4836 276020 4848
rect 276072 4836 276078 4888
rect 44542 4768 44548 4820
rect 44600 4808 44606 4820
rect 132494 4808 132500 4820
rect 44600 4780 132500 4808
rect 44600 4768 44606 4780
rect 132494 4768 132500 4780
rect 132552 4768 132558 4820
rect 132586 4768 132592 4820
rect 132644 4808 132650 4820
rect 134610 4808 134616 4820
rect 132644 4780 134616 4808
rect 132644 4768 132650 4780
rect 134610 4768 134616 4780
rect 134668 4768 134674 4820
rect 134886 4768 134892 4820
rect 134944 4808 134950 4820
rect 278774 4808 278780 4820
rect 134944 4780 278780 4808
rect 134944 4768 134950 4780
rect 278774 4768 278780 4780
rect 278832 4768 278838 4820
rect 52822 4700 52828 4752
rect 52880 4740 52886 4752
rect 65518 4740 65524 4752
rect 52880 4712 65524 4740
rect 52880 4700 52886 4712
rect 65518 4700 65524 4712
rect 65576 4700 65582 4752
rect 76650 4700 76656 4752
rect 76708 4740 76714 4752
rect 184934 4740 184940 4752
rect 76708 4712 184940 4740
rect 76708 4700 76714 4712
rect 184934 4700 184940 4712
rect 184992 4700 184998 4752
rect 73062 4632 73068 4684
rect 73120 4672 73126 4684
rect 179414 4672 179420 4684
rect 73120 4644 179420 4672
rect 73120 4632 73126 4644
rect 179414 4632 179420 4644
rect 179472 4632 179478 4684
rect 69474 4564 69480 4616
rect 69532 4604 69538 4616
rect 172514 4604 172520 4616
rect 69532 4576 172520 4604
rect 69532 4564 69538 4576
rect 172514 4564 172520 4576
rect 172572 4564 172578 4616
rect 65978 4496 65984 4548
rect 66036 4536 66042 4548
rect 166994 4536 167000 4548
rect 66036 4508 167000 4536
rect 66036 4496 66042 4508
rect 166994 4496 167000 4508
rect 167052 4496 167058 4548
rect 62390 4428 62396 4480
rect 62448 4468 62454 4480
rect 161474 4468 161480 4480
rect 62448 4440 161480 4468
rect 62448 4428 62454 4440
rect 161474 4428 161480 4440
rect 161532 4428 161538 4480
rect 58802 4360 58808 4412
rect 58860 4400 58866 4412
rect 155954 4400 155960 4412
rect 58860 4372 155960 4400
rect 58860 4360 58866 4372
rect 155954 4360 155960 4372
rect 156012 4360 156018 4412
rect 55214 4292 55220 4344
rect 55272 4332 55278 4344
rect 150434 4332 150440 4344
rect 55272 4304 150440 4332
rect 55272 4292 55278 4304
rect 150434 4292 150440 4304
rect 150492 4292 150498 4344
rect 51626 4224 51632 4276
rect 51684 4264 51690 4276
rect 143534 4264 143540 4276
rect 51684 4236 143540 4264
rect 51684 4224 51690 4236
rect 143534 4224 143540 4236
rect 143592 4224 143598 4276
rect 48222 4156 48228 4208
rect 48280 4196 48286 4208
rect 138014 4196 138020 4208
rect 48280 4168 138020 4196
rect 48280 4156 48286 4168
rect 138014 4156 138020 4168
rect 138072 4156 138078 4208
rect 3970 4088 3976 4140
rect 4028 4128 4034 4140
rect 61102 4128 61108 4140
rect 4028 4100 61108 4128
rect 4028 4088 4034 4100
rect 61102 4088 61108 4100
rect 61160 4088 61166 4140
rect 61194 4088 61200 4140
rect 61252 4128 61258 4140
rect 62022 4128 62028 4140
rect 61252 4100 62028 4128
rect 61252 4088 61258 4100
rect 62022 4088 62028 4100
rect 62080 4088 62086 4140
rect 68278 4088 68284 4140
rect 68336 4128 68342 4140
rect 73338 4128 73344 4140
rect 68336 4100 73344 4128
rect 68336 4088 68342 4100
rect 73338 4088 73344 4100
rect 73396 4088 73402 4140
rect 81434 4128 81440 4140
rect 74644 4100 81440 4128
rect 8846 4020 8852 4072
rect 8904 4060 8910 4072
rect 74534 4060 74540 4072
rect 8904 4032 74540 4060
rect 8904 4020 8910 4032
rect 74534 4020 74540 4032
rect 74592 4020 74598 4072
rect 13630 3952 13636 4004
rect 13688 3992 13694 4004
rect 74644 3992 74672 4100
rect 81434 4088 81440 4100
rect 81492 4088 81498 4140
rect 81544 4100 82952 4128
rect 77846 4020 77852 4072
rect 77904 4060 77910 4072
rect 81544 4060 81572 4100
rect 77904 4032 81572 4060
rect 77904 4020 77910 4032
rect 82630 4020 82636 4072
rect 82688 4060 82694 4072
rect 82924 4060 82952 4100
rect 82998 4088 83004 4140
rect 83056 4128 83062 4140
rect 183554 4128 183560 4140
rect 83056 4100 183560 4128
rect 83056 4088 83062 4100
rect 183554 4088 183560 4100
rect 183612 4088 183618 4140
rect 186314 4060 186320 4072
rect 82688 4032 82860 4060
rect 82924 4032 186320 4060
rect 82688 4020 82694 4032
rect 13688 3964 74672 3992
rect 13688 3952 13694 3964
rect 75454 3952 75460 4004
rect 75512 3992 75518 4004
rect 78950 3992 78956 4004
rect 75512 3964 78956 3992
rect 75512 3952 75518 3964
rect 78950 3952 78956 3964
rect 79008 3952 79014 4004
rect 79042 3952 79048 4004
rect 79100 3992 79106 4004
rect 79962 3992 79968 4004
rect 79100 3964 79968 3992
rect 79100 3952 79106 3964
rect 79962 3952 79968 3964
rect 80020 3952 80026 4004
rect 81434 3952 81440 4004
rect 81492 3992 81498 4004
rect 82722 3992 82728 4004
rect 81492 3964 82728 3992
rect 81492 3952 81498 3964
rect 82722 3952 82728 3964
rect 82780 3952 82786 4004
rect 82832 3992 82860 4032
rect 186314 4020 186320 4032
rect 186372 4020 186378 4072
rect 194594 3992 194600 4004
rect 82832 3964 194600 3992
rect 194594 3952 194600 3964
rect 194652 3952 194658 4004
rect 18322 3884 18328 3936
rect 18380 3924 18386 3936
rect 86034 3924 86040 3936
rect 18380 3896 86040 3924
rect 18380 3884 18386 3896
rect 86034 3884 86040 3896
rect 86092 3884 86098 3936
rect 86126 3884 86132 3936
rect 86184 3924 86190 3936
rect 86862 3924 86868 3936
rect 86184 3896 86868 3924
rect 86184 3884 86190 3896
rect 86862 3884 86868 3896
rect 86920 3884 86926 3936
rect 88518 3884 88524 3936
rect 88576 3924 88582 3936
rect 89622 3924 89628 3936
rect 88576 3896 89628 3924
rect 88576 3884 88582 3896
rect 89622 3884 89628 3896
rect 89680 3884 89686 3936
rect 89714 3884 89720 3936
rect 89772 3924 89778 3936
rect 93210 3924 93216 3936
rect 89772 3896 93216 3924
rect 89772 3884 89778 3896
rect 93210 3884 93216 3896
rect 93268 3884 93274 3936
rect 93302 3884 93308 3936
rect 93360 3924 93366 3936
rect 93762 3924 93768 3936
rect 93360 3896 93768 3924
rect 93360 3884 93366 3896
rect 93762 3884 93768 3896
rect 93820 3884 93826 3936
rect 93854 3884 93860 3936
rect 93912 3924 93918 3936
rect 205634 3924 205640 3936
rect 93912 3896 205640 3924
rect 93912 3884 93918 3896
rect 205634 3884 205640 3896
rect 205692 3884 205698 3936
rect 24302 3816 24308 3868
rect 24360 3856 24366 3868
rect 24762 3856 24768 3868
rect 24360 3828 24768 3856
rect 24360 3816 24366 3828
rect 24762 3816 24768 3828
rect 24820 3816 24826 3868
rect 25498 3816 25504 3868
rect 25556 3856 25562 3868
rect 26142 3856 26148 3868
rect 25556 3828 26148 3856
rect 25556 3816 25562 3828
rect 26142 3816 26148 3828
rect 26200 3816 26206 3868
rect 95510 3856 95516 3868
rect 26252 3828 95516 3856
rect 23106 3748 23112 3800
rect 23164 3788 23170 3800
rect 26252 3788 26280 3828
rect 95510 3816 95516 3828
rect 95568 3816 95574 3868
rect 95620 3828 96660 3856
rect 23164 3760 26280 3788
rect 23164 3748 23170 3760
rect 27890 3748 27896 3800
rect 27948 3788 27954 3800
rect 95620 3788 95648 3828
rect 27948 3760 95648 3788
rect 27948 3748 27954 3760
rect 95694 3748 95700 3800
rect 95752 3788 95758 3800
rect 96522 3788 96528 3800
rect 95752 3760 96528 3788
rect 95752 3748 95758 3760
rect 96522 3748 96528 3760
rect 96580 3748 96586 3800
rect 96632 3788 96660 3828
rect 96890 3816 96896 3868
rect 96948 3856 96954 3868
rect 218054 3856 218060 3868
rect 96948 3828 218060 3856
rect 96948 3816 96954 3828
rect 218054 3816 218060 3828
rect 218112 3816 218118 3868
rect 102686 3788 102692 3800
rect 96632 3760 102692 3788
rect 102686 3748 102692 3760
rect 102744 3748 102750 3800
rect 102778 3748 102784 3800
rect 102836 3788 102842 3800
rect 103422 3788 103428 3800
rect 102836 3760 103428 3788
rect 102836 3748 102842 3760
rect 103422 3748 103428 3760
rect 103480 3748 103486 3800
rect 106366 3748 106372 3800
rect 106424 3788 106430 3800
rect 107562 3788 107568 3800
rect 106424 3760 107568 3788
rect 106424 3748 106430 3760
rect 107562 3748 107568 3760
rect 107620 3748 107626 3800
rect 107654 3748 107660 3800
rect 107712 3788 107718 3800
rect 113174 3788 113180 3800
rect 107712 3760 113180 3788
rect 107712 3748 107718 3760
rect 113174 3748 113180 3760
rect 113232 3748 113238 3800
rect 113542 3748 113548 3800
rect 113600 3788 113606 3800
rect 114462 3788 114468 3800
rect 113600 3760 114468 3788
rect 113600 3748 113606 3760
rect 114462 3748 114468 3760
rect 114520 3748 114526 3800
rect 114738 3748 114744 3800
rect 114796 3788 114802 3800
rect 115842 3788 115848 3800
rect 114796 3760 115848 3788
rect 114796 3748 114802 3760
rect 115842 3748 115848 3760
rect 115900 3748 115906 3800
rect 238754 3788 238760 3800
rect 115952 3760 238760 3788
rect 31478 3680 31484 3732
rect 31536 3720 31542 3732
rect 110414 3720 110420 3732
rect 31536 3692 110420 3720
rect 31536 3680 31542 3692
rect 110414 3680 110420 3692
rect 110472 3680 110478 3732
rect 34974 3612 34980 3664
rect 35032 3652 35038 3664
rect 109862 3652 109868 3664
rect 35032 3624 109868 3652
rect 35032 3612 35038 3624
rect 109862 3612 109868 3624
rect 109920 3612 109926 3664
rect 109954 3612 109960 3664
rect 110012 3652 110018 3664
rect 115952 3652 115980 3760
rect 238754 3748 238760 3760
rect 238812 3748 238818 3800
rect 241514 3720 241520 3732
rect 110012 3624 115980 3652
rect 116136 3692 241520 3720
rect 110012 3612 110018 3624
rect 32674 3544 32680 3596
rect 32732 3584 32738 3596
rect 107654 3584 107660 3596
rect 32732 3556 107660 3584
rect 32732 3544 32738 3556
rect 107654 3544 107660 3556
rect 107712 3544 107718 3596
rect 111150 3544 111156 3596
rect 111208 3584 111214 3596
rect 116136 3584 116164 3692
rect 241514 3680 241520 3692
rect 241572 3680 241578 3732
rect 117130 3612 117136 3664
rect 117188 3652 117194 3664
rect 117188 3624 120580 3652
rect 117188 3612 117194 3624
rect 111208 3556 116164 3584
rect 111208 3544 111214 3556
rect 118234 3544 118240 3596
rect 118292 3584 118298 3596
rect 120552 3584 120580 3624
rect 120626 3612 120632 3664
rect 120684 3652 120690 3664
rect 121362 3652 121368 3664
rect 120684 3624 121368 3652
rect 120684 3612 120690 3624
rect 121362 3612 121368 3624
rect 121420 3612 121426 3664
rect 121822 3612 121828 3664
rect 121880 3652 121886 3664
rect 122742 3652 122748 3664
rect 121880 3624 122748 3652
rect 121880 3612 121886 3624
rect 122742 3612 122748 3624
rect 122800 3612 122806 3664
rect 122834 3612 122840 3664
rect 122892 3652 122898 3664
rect 252554 3652 252560 3664
rect 122892 3624 252560 3652
rect 122892 3612 122898 3624
rect 252554 3612 252560 3624
rect 252612 3612 252618 3664
rect 251174 3584 251180 3596
rect 118292 3556 120488 3584
rect 120552 3556 122788 3584
rect 118292 3544 118298 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 4062 3516 4068 3528
rect 2924 3488 4068 3516
rect 2924 3476 2930 3488
rect 4062 3476 4068 3488
rect 4120 3476 4126 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16482 3516 16488 3528
rect 16080 3488 16488 3516
rect 16080 3476 16086 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 19518 3476 19524 3528
rect 19576 3516 19582 3528
rect 20622 3516 20628 3528
rect 19576 3488 20628 3516
rect 19576 3476 19582 3488
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 21910 3516 21916 3528
rect 20772 3488 21916 3516
rect 20772 3476 20778 3488
rect 21910 3476 21916 3488
rect 21968 3476 21974 3528
rect 42150 3476 42156 3528
rect 42208 3516 42214 3528
rect 42702 3516 42708 3528
rect 42208 3488 42708 3516
rect 42208 3476 42214 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 45370 3476 45376 3528
rect 45428 3516 45434 3528
rect 74626 3516 74632 3528
rect 45428 3488 74632 3516
rect 45428 3476 45434 3488
rect 74626 3476 74632 3488
rect 74684 3476 74690 3528
rect 84010 3476 84016 3528
rect 84068 3516 84074 3528
rect 93946 3516 93952 3528
rect 84068 3488 93952 3516
rect 84068 3476 84074 3488
rect 93946 3476 93952 3488
rect 94004 3476 94010 3528
rect 99466 3476 99472 3528
rect 99524 3516 99530 3528
rect 118786 3516 118792 3528
rect 99524 3488 118792 3516
rect 99524 3476 99530 3488
rect 118786 3476 118792 3488
rect 118844 3476 118850 3528
rect 120460 3516 120488 3556
rect 122650 3516 122656 3528
rect 120460 3488 122656 3516
rect 122650 3476 122656 3488
rect 122708 3476 122714 3528
rect 122760 3516 122788 3556
rect 123036 3556 251180 3584
rect 123036 3516 123064 3556
rect 251174 3544 251180 3556
rect 251232 3544 251238 3596
rect 122760 3488 123064 3516
rect 124214 3476 124220 3528
rect 124272 3516 124278 3528
rect 262214 3516 262220 3528
rect 124272 3488 262220 3516
rect 124272 3476 124278 3488
rect 262214 3476 262220 3488
rect 262272 3476 262278 3528
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 32398 3448 32404 3460
rect 11296 3420 32404 3448
rect 11296 3408 11302 3420
rect 32398 3408 32404 3420
rect 32456 3408 32462 3460
rect 45462 3408 45468 3460
rect 45520 3448 45526 3460
rect 46842 3448 46848 3460
rect 45520 3420 46848 3448
rect 45520 3408 45526 3420
rect 46842 3408 46848 3420
rect 46900 3408 46906 3460
rect 46934 3408 46940 3460
rect 46992 3448 46998 3460
rect 48130 3448 48136 3460
rect 46992 3420 48136 3448
rect 46992 3408 46998 3420
rect 48130 3408 48136 3420
rect 48188 3408 48194 3460
rect 50522 3408 50528 3460
rect 50580 3448 50586 3460
rect 50982 3448 50988 3460
rect 50580 3420 50988 3448
rect 50580 3408 50586 3420
rect 50982 3408 50988 3420
rect 51040 3408 51046 3460
rect 61102 3408 61108 3460
rect 61160 3448 61166 3460
rect 66254 3448 66260 3460
rect 61160 3420 66260 3448
rect 61160 3408 61166 3420
rect 66254 3408 66260 3420
rect 66312 3408 66318 3460
rect 71866 3408 71872 3460
rect 71924 3448 71930 3460
rect 72970 3448 72976 3460
rect 71924 3420 72976 3448
rect 71924 3408 71930 3420
rect 72970 3408 72976 3420
rect 73028 3408 73034 3460
rect 84102 3408 84108 3460
rect 84160 3448 84166 3460
rect 93854 3448 93860 3460
rect 84160 3420 93860 3448
rect 84160 3408 84166 3420
rect 93854 3408 93860 3420
rect 93912 3408 93918 3460
rect 99374 3408 99380 3460
rect 99432 3448 99438 3460
rect 122926 3448 122932 3460
rect 99432 3420 122932 3448
rect 99432 3408 99438 3420
rect 122926 3408 122932 3420
rect 122984 3408 122990 3460
rect 125410 3408 125416 3460
rect 125468 3448 125474 3460
rect 264974 3448 264980 3460
rect 125468 3420 264980 3448
rect 125468 3408 125474 3420
rect 264974 3408 264980 3420
rect 265032 3408 265038 3460
rect 566 3340 572 3392
rect 624 3380 630 3392
rect 59170 3380 59176 3392
rect 624 3352 59176 3380
rect 624 3340 630 3352
rect 59170 3340 59176 3352
rect 59228 3340 59234 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64138 3380 64144 3392
rect 63644 3352 64144 3380
rect 63644 3340 63650 3352
rect 64138 3340 64144 3352
rect 64196 3340 64202 3392
rect 73246 3340 73252 3392
rect 73304 3380 73310 3392
rect 175274 3380 175280 3392
rect 73304 3352 175280 3380
rect 73304 3340 73310 3352
rect 175274 3340 175280 3352
rect 175332 3340 175338 3392
rect 1670 3272 1676 3324
rect 1728 3312 1734 3324
rect 62206 3312 62212 3324
rect 1728 3284 62212 3312
rect 1728 3272 1734 3284
rect 62206 3272 62212 3284
rect 62264 3272 62270 3324
rect 68646 3312 68652 3324
rect 64064 3284 68652 3312
rect 6454 3204 6460 3256
rect 6512 3244 6518 3256
rect 6914 3244 6920 3256
rect 6512 3216 6920 3244
rect 6512 3204 6518 3216
rect 6914 3204 6920 3216
rect 6972 3204 6978 3256
rect 21358 3204 21364 3256
rect 21416 3244 21422 3256
rect 35894 3244 35900 3256
rect 21416 3216 35900 3244
rect 21416 3204 21422 3216
rect 35894 3204 35900 3216
rect 35952 3204 35958 3256
rect 36170 3204 36176 3256
rect 36228 3244 36234 3256
rect 45370 3244 45376 3256
rect 36228 3216 45376 3244
rect 36228 3204 36234 3216
rect 45370 3204 45376 3216
rect 45428 3204 45434 3256
rect 46842 3204 46848 3256
rect 46900 3244 46906 3256
rect 64064 3244 64092 3284
rect 68646 3272 68652 3284
rect 68704 3272 68710 3324
rect 73338 3272 73344 3324
rect 73396 3312 73402 3324
rect 171134 3312 171140 3324
rect 73396 3284 171140 3312
rect 73396 3272 73402 3284
rect 171134 3272 171140 3284
rect 171192 3272 171198 3324
rect 46900 3216 64092 3244
rect 46900 3204 46906 3216
rect 64138 3204 64144 3256
rect 64196 3244 64202 3256
rect 162854 3244 162860 3256
rect 64196 3216 162860 3244
rect 64196 3204 64202 3216
rect 162854 3204 162860 3216
rect 162912 3204 162918 3256
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 5316 3148 24348 3176
rect 5316 3136 5322 3148
rect 6914 3068 6920 3120
rect 6972 3108 6978 3120
rect 21358 3108 21364 3120
rect 6972 3080 21364 3108
rect 6972 3068 6978 3080
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 24320 3108 24348 3148
rect 26804 3148 36124 3176
rect 26804 3108 26832 3148
rect 24320 3080 26832 3108
rect 29086 3068 29092 3120
rect 29144 3108 29150 3120
rect 36096 3108 36124 3148
rect 57606 3136 57612 3188
rect 57664 3176 57670 3188
rect 153194 3176 153200 3188
rect 57664 3148 153200 3176
rect 57664 3136 57670 3148
rect 153194 3136 153200 3148
rect 153252 3136 153258 3188
rect 39298 3108 39304 3120
rect 29144 3080 35940 3108
rect 36096 3080 39304 3108
rect 29144 3068 29150 3080
rect 35912 2972 35940 3080
rect 39298 3068 39304 3080
rect 39356 3068 39362 3120
rect 56410 3068 56416 3120
rect 56468 3108 56474 3120
rect 151814 3108 151820 3120
rect 56468 3080 151820 3108
rect 56468 3068 56474 3080
rect 151814 3068 151820 3080
rect 151872 3068 151878 3120
rect 35986 3000 35992 3052
rect 36044 3040 36050 3052
rect 51810 3040 51816 3052
rect 36044 3012 51816 3040
rect 36044 3000 36050 3012
rect 51810 3000 51816 3012
rect 51868 3000 51874 3052
rect 54018 3000 54024 3052
rect 54076 3040 54082 3052
rect 147674 3040 147680 3052
rect 54076 3012 147680 3040
rect 54076 3000 54082 3012
rect 147674 3000 147680 3012
rect 147732 3000 147738 3052
rect 42058 2972 42064 2984
rect 35912 2944 42064 2972
rect 42058 2932 42064 2944
rect 42116 2932 42122 2984
rect 49326 2932 49332 2984
rect 49384 2972 49390 2984
rect 139394 2972 139400 2984
rect 49384 2944 139400 2972
rect 49384 2932 49390 2944
rect 139394 2932 139400 2944
rect 139452 2932 139458 2984
rect 38562 2864 38568 2916
rect 38620 2904 38626 2916
rect 45462 2904 45468 2916
rect 38620 2876 45468 2904
rect 38620 2864 38626 2876
rect 45462 2864 45468 2876
rect 45520 2864 45526 2916
rect 45738 2864 45744 2916
rect 45796 2904 45802 2916
rect 133966 2904 133972 2916
rect 45796 2876 133972 2904
rect 45796 2864 45802 2876
rect 133966 2864 133972 2876
rect 134024 2864 134030 2916
rect 43346 2796 43352 2848
rect 43404 2836 43410 2848
rect 129826 2836 129832 2848
rect 43404 2808 124168 2836
rect 43404 2796 43410 2808
rect 124140 2768 124168 2808
rect 127820 2808 129832 2836
rect 127820 2768 127848 2808
rect 129826 2796 129832 2808
rect 129884 2796 129890 2848
rect 124140 2740 127848 2768
rect 70670 1096 70676 1148
rect 70728 1136 70734 1148
rect 73246 1136 73252 1148
rect 70728 1108 73252 1136
rect 70728 1096 70734 1108
rect 73246 1096 73252 1108
rect 73304 1096 73310 1148
<< via1 >>
rect 58808 700952 58860 701004
rect 202788 700952 202840 701004
rect 58716 700884 58768 700936
rect 218980 700884 219032 700936
rect 58992 700816 59044 700868
rect 267648 700816 267700 700868
rect 58900 700748 58952 700800
rect 283840 700748 283892 700800
rect 59084 700680 59136 700732
rect 332508 700680 332560 700732
rect 57704 700612 57756 700664
rect 348792 700612 348844 700664
rect 59176 700544 59228 700596
rect 397460 700544 397512 700596
rect 57796 700476 57848 700528
rect 413652 700476 413704 700528
rect 57888 700408 57940 700460
rect 478512 700408 478564 700460
rect 59268 700340 59320 700392
rect 527180 700340 527232 700392
rect 59360 700272 59412 700324
rect 543464 700272 543516 700324
rect 58532 700204 58584 700256
rect 136640 700204 136692 700256
rect 137284 700204 137336 700256
rect 235172 700204 235224 700256
rect 57612 700136 57664 700188
rect 154120 700136 154172 700188
rect 57520 700068 57572 700120
rect 89168 700068 89220 700120
rect 136640 700068 136692 700120
rect 137836 700068 137888 700120
rect 58440 700000 58492 700052
rect 72976 700000 73028 700052
rect 40500 699932 40552 699984
rect 42064 699932 42116 699984
rect 8116 699660 8168 699712
rect 10324 699660 10376 699712
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 104992 698232 105044 698284
rect 105544 698232 105596 698284
rect 364432 698232 364484 698284
rect 365076 698232 365128 698284
rect 560300 697280 560352 697332
rect 565176 697280 565228 697332
rect 166908 697144 166960 697196
rect 172428 697144 172480 697196
rect 540980 697144 541032 697196
rect 548616 697144 548668 697196
rect 70308 697076 70360 697128
rect 77208 697076 77260 697128
rect 89628 697076 89680 697128
rect 96528 697076 96580 697128
rect 108948 697076 109000 697128
rect 115848 697076 115900 697128
rect 128268 697076 128320 697128
rect 135168 697076 135220 697128
rect 147588 697076 147640 697128
rect 154488 697076 154540 697128
rect 186228 697076 186280 697128
rect 193128 697076 193180 697128
rect 205548 697076 205600 697128
rect 212448 697076 212500 697128
rect 224868 697076 224920 697128
rect 231768 697076 231820 697128
rect 244188 697076 244240 697128
rect 251088 697076 251140 697128
rect 263508 697076 263560 697128
rect 270408 697076 270460 697128
rect 282828 697076 282880 697128
rect 289728 697076 289780 697128
rect 302148 697076 302200 697128
rect 309048 697076 309100 697128
rect 321468 697076 321520 697128
rect 328368 697076 328420 697128
rect 169760 695444 169812 695496
rect 170036 695444 170088 695496
rect 429200 692792 429252 692844
rect 429936 692792 429988 692844
rect 494060 692792 494112 692844
rect 494888 692792 494940 692844
rect 173900 686264 173952 686316
rect 178776 686264 178828 686316
rect 367100 686264 367152 686316
rect 371976 686264 372028 686316
rect 560300 686264 560352 686316
rect 565176 686264 565228 686316
rect 154580 686128 154632 686180
rect 162216 686128 162268 686180
rect 289820 686128 289872 686180
rect 294512 686128 294564 686180
rect 347780 686128 347832 686180
rect 355416 686128 355468 686180
rect 540980 686128 541032 686180
rect 548616 686128 548668 686180
rect 169760 685856 169812 685908
rect 169944 685856 169996 685908
rect 299572 685856 299624 685908
rect 300124 685856 300176 685908
rect 559012 684496 559064 684548
rect 559656 684496 559708 684548
rect 299572 684428 299624 684480
rect 299664 684428 299716 684480
rect 2780 681708 2832 681760
rect 5080 681708 5132 681760
rect 299664 678988 299716 679040
rect 299572 678920 299624 678972
rect 429200 676132 429252 676184
rect 429292 676132 429344 676184
rect 559012 674840 559064 674892
rect 559380 674840 559432 674892
rect 173900 673888 173952 673940
rect 178776 673888 178828 673940
rect 367100 673888 367152 673940
rect 371976 673888 372028 673940
rect 560300 673888 560352 673940
rect 565176 673888 565228 673940
rect 154580 673752 154632 673804
rect 162216 673752 162268 673804
rect 289820 673752 289872 673804
rect 292672 673752 292724 673804
rect 347780 673752 347832 673804
rect 355416 673752 355468 673804
rect 540980 673752 541032 673804
rect 548616 673752 548668 673804
rect 104900 673480 104952 673532
rect 105084 673480 105136 673532
rect 494060 673480 494112 673532
rect 494244 673480 494296 673532
rect 364432 669400 364484 669452
rect 364432 669264 364484 669316
rect 3424 667904 3476 667956
rect 21364 667904 21416 667956
rect 299572 666544 299624 666596
rect 299756 666544 299808 666596
rect 429292 666544 429344 666596
rect 429384 666544 429436 666596
rect 559104 661716 559156 661768
rect 559380 661716 559432 661768
rect 170036 659676 170088 659728
rect 299756 659676 299808 659728
rect 429384 659676 429436 659728
rect 169944 659608 169996 659660
rect 299572 659608 299624 659660
rect 429292 659608 429344 659660
rect 559104 656888 559156 656940
rect 559196 656888 559248 656940
rect 169760 655460 169812 655512
rect 169944 655460 169996 655512
rect 104900 654100 104952 654152
rect 105084 654100 105136 654152
rect 364340 654100 364392 654152
rect 364524 654100 364576 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 507860 653352 507912 653404
rect 513380 653352 513432 653404
rect 513380 652808 513432 652860
rect 518900 652808 518952 652860
rect 3056 652740 3108 652792
rect 13084 652740 13136 652792
rect 129280 652740 129332 652792
rect 133604 652740 133656 652792
rect 139584 652740 139636 652792
rect 259184 652740 259236 652792
rect 263784 652740 263836 652792
rect 269120 652740 269172 652792
rect 378508 652740 378560 652792
rect 383476 652740 383528 652792
rect 389364 652740 389416 652792
rect 507860 652740 507912 652792
rect 57428 650836 57480 650888
rect 104900 650836 104952 650888
rect 59544 650768 59596 650820
rect 364340 650768 364392 650820
rect 58348 650700 58400 650752
rect 462320 650700 462372 650752
rect 59452 650632 59504 650684
rect 494060 650632 494112 650684
rect 139400 650360 139452 650412
rect 266360 650360 266412 650412
rect 282000 650360 282052 650412
rect 389180 650360 389232 650412
rect 516416 650360 516468 650412
rect 58624 650292 58676 650344
rect 580172 650292 580224 650344
rect 266360 650020 266412 650072
rect 281540 650020 281592 650072
rect 282000 650020 282052 650072
rect 299572 649952 299624 650004
rect 299756 649952 299808 650004
rect 429292 649952 429344 650004
rect 429476 649952 429528 650004
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 142068 645872 142120 645924
rect 187700 645872 187752 645924
rect 291936 645872 291988 645924
rect 307392 645872 307444 645924
rect 399484 645872 399536 645924
rect 437480 645872 437532 645924
rect 140688 644444 140740 644496
rect 187700 644444 187752 644496
rect 290556 644444 290608 644496
rect 307116 644444 307168 644496
rect 398104 644444 398156 644496
rect 437480 644444 437532 644496
rect 137928 643084 137980 643136
rect 187700 643084 187752 643136
rect 287704 643084 287756 643136
rect 307116 643084 307168 643136
rect 395344 643084 395396 643136
rect 437480 643084 437532 643136
rect 299480 642336 299532 642388
rect 299756 642336 299808 642388
rect 160744 641724 160796 641776
rect 187700 641724 187752 641776
rect 286324 641724 286376 641776
rect 307668 641724 307720 641776
rect 393964 641724 394016 641776
rect 437480 641724 437532 641776
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 159364 640296 159416 640348
rect 187700 640296 187752 640348
rect 284944 640296 284996 640348
rect 307668 640296 307720 640348
rect 392584 640296 392636 640348
rect 437480 640296 437532 640348
rect 283564 638936 283616 638988
rect 306656 638936 306708 638988
rect 391204 638936 391256 638988
rect 437480 638936 437532 638988
rect 299480 637644 299532 637696
rect 294604 637576 294656 637628
rect 299572 637576 299624 637628
rect 299664 637576 299716 637628
rect 388444 637576 388496 637628
rect 437480 637576 437532 637628
rect 429200 637508 429252 637560
rect 429384 637508 429436 637560
rect 169668 636216 169720 636268
rect 169944 636216 169996 636268
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 169668 627920 169720 627972
rect 170036 627920 170088 627972
rect 299848 627920 299900 627972
rect 300032 627920 300084 627972
rect 429200 627920 429252 627972
rect 429568 627920 429620 627972
rect 3884 623772 3936 623824
rect 5172 623772 5224 623824
rect 299848 621052 299900 621104
rect 429568 621052 429620 621104
rect 299756 620916 299808 620968
rect 429476 620916 429528 620968
rect 169852 618264 169904 618316
rect 170036 618264 170088 618316
rect 169944 611396 169996 611448
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 170036 611192 170088 611244
rect 3424 609968 3476 610020
rect 31024 609968 31076 610020
rect 299572 608540 299624 608592
rect 299664 608540 299716 608592
rect 429292 608540 429344 608592
rect 429384 608540 429436 608592
rect 559012 608540 559064 608592
rect 559104 608540 559156 608592
rect 299572 601672 299624 601724
rect 299848 601672 299900 601724
rect 429292 601672 429344 601724
rect 429568 601672 429620 601724
rect 559012 601672 559064 601724
rect 559288 601672 559340 601724
rect 169852 598952 169904 599004
rect 170036 598952 170088 599004
rect 299664 598884 299716 598936
rect 299848 598884 299900 598936
rect 429384 598884 429436 598936
rect 429568 598884 429620 598936
rect 559104 598884 559156 598936
rect 559288 598884 559340 598936
rect 3240 594804 3292 594856
rect 14464 594804 14516 594856
rect 169944 592084 169996 592136
rect 170036 591880 170088 591932
rect 299664 589296 299716 589348
rect 299940 589296 299992 589348
rect 429384 589296 429436 589348
rect 429660 589296 429712 589348
rect 559104 589296 559156 589348
rect 559380 589296 559432 589348
rect 299940 582428 299992 582480
rect 429660 582428 429712 582480
rect 559380 582428 559432 582480
rect 299848 582292 299900 582344
rect 429568 582292 429620 582344
rect 559288 582292 559340 582344
rect 270040 580252 270092 580304
rect 281632 580252 281684 580304
rect 177948 579640 178000 579692
rect 187700 579640 187752 579692
rect 285036 579640 285088 579692
rect 306932 579640 306984 579692
rect 402244 579640 402296 579692
rect 437480 579640 437532 579692
rect 170128 578212 170180 578264
rect 170312 578212 170364 578264
rect 282184 578212 282236 578264
rect 306380 578212 306432 578264
rect 170128 572704 170180 572756
rect 170128 572568 170180 572620
rect 3976 567196 4028 567248
rect 5264 567196 5316 567248
rect 170128 563116 170180 563168
rect 170036 562980 170088 563032
rect 281724 561620 281776 561672
rect 282184 561620 282236 561672
rect 59636 560872 59688 560924
rect 188988 560872 189040 560924
rect 281724 560872 281776 560924
rect 306288 560872 306340 560924
rect 438124 560872 438176 560924
rect 559012 560260 559064 560312
rect 559104 560260 559156 560312
rect 79324 558832 79376 558884
rect 81440 558832 81492 558884
rect 81532 558832 81584 558884
rect 86868 558832 86920 558884
rect 80704 558764 80756 558816
rect 90088 558832 90140 558884
rect 91008 558832 91060 558884
rect 335452 558832 335504 558884
rect 344284 558832 344336 558884
rect 355324 558832 355376 558884
rect 483020 558832 483072 558884
rect 87880 558764 87932 558816
rect 96620 558764 96672 558816
rect 223580 558764 223632 558816
rect 231952 558764 232004 558816
rect 343732 558764 343784 558816
rect 351920 558764 351972 558816
rect 458824 558764 458876 558816
rect 468024 558764 468076 558816
rect 477132 558764 477184 558816
rect 485780 558764 485832 558816
rect 79508 558696 79560 558748
rect 88984 558696 89036 558748
rect 77392 558628 77444 558680
rect 81532 558628 81584 558680
rect 81624 558628 81676 558680
rect 91376 558628 91428 558680
rect 100300 558696 100352 558748
rect 216772 558696 216824 558748
rect 225788 558696 225840 558748
rect 226340 558696 226392 558748
rect 227168 558696 227220 558748
rect 236000 558696 236052 558748
rect 344284 558696 344336 558748
rect 353300 558696 353352 558748
rect 460664 558696 460716 558748
rect 468576 558696 468628 558748
rect 475568 558696 475620 558748
rect 484400 558696 484452 558748
rect 95332 558628 95384 558680
rect 105360 558628 105412 558680
rect 106096 558628 106148 558680
rect 215300 558628 215352 558680
rect 224408 558628 224460 558680
rect 233240 558628 233292 558680
rect 338948 558628 339000 558680
rect 348332 558628 348384 558680
rect 357440 558628 357492 558680
rect 75736 558560 75788 558612
rect 84292 558560 84344 558612
rect 93584 558560 93636 558612
rect 108580 558560 108632 558612
rect 211344 558560 211396 558612
rect 212540 558560 212592 558612
rect 213184 558560 213236 558612
rect 222292 558560 222344 558612
rect 231860 558560 231912 558612
rect 336648 558560 336700 558612
rect 346308 558560 346360 558612
rect 346952 558560 347004 558612
rect 356060 558560 356112 558612
rect 356796 558560 356848 558612
rect 484492 558628 484544 558680
rect 453488 558560 453540 558612
rect 462964 558560 463016 558612
rect 463608 558560 463660 558612
rect 464344 558560 464396 558612
rect 473544 558560 473596 558612
rect 483020 558560 483072 558612
rect 72424 558492 72476 558544
rect 81624 558492 81676 558544
rect 86868 558492 86920 558544
rect 95332 558492 95384 558544
rect 96620 558492 96672 558544
rect 106280 558492 106332 558544
rect 107476 558492 107528 558544
rect 107844 558492 107896 558544
rect 209780 558492 209832 558544
rect 211160 558492 211212 558544
rect 211896 558492 211948 558544
rect 221096 558492 221148 558544
rect 230480 558492 230532 558544
rect 337384 558492 337436 558544
rect 460388 558492 460440 558544
rect 460848 558492 460900 558544
rect 470048 558492 470100 558544
rect 479432 558492 479484 558544
rect 488540 558492 488592 558544
rect 76012 558424 76064 558476
rect 85396 558424 85448 558476
rect 94596 558424 94648 558476
rect 103980 558424 104032 558476
rect 104716 558424 104768 558476
rect 166908 558424 166960 558476
rect 201500 558424 201552 558476
rect 331312 558424 331364 558476
rect 331772 558424 331824 558476
rect 340972 558424 341024 558476
rect 350540 558424 350592 558476
rect 453304 558424 453356 558476
rect 461768 558424 461820 558476
rect 471244 558424 471296 558476
rect 480444 558424 480496 558476
rect 73712 558356 73764 558408
rect 82912 558356 82964 558408
rect 92480 558356 92532 558408
rect 100760 558356 100812 558408
rect 165528 558356 165580 558408
rect 200212 558356 200264 558408
rect 218060 558356 218112 558408
rect 218888 558356 218940 558408
rect 227720 558356 227772 558408
rect 227812 558356 227864 558408
rect 229468 558356 229520 558408
rect 238760 558356 238812 558408
rect 332692 558356 332744 558408
rect 342536 558356 342588 558408
rect 347964 558356 348016 558408
rect 358176 558356 358228 558408
rect 455420 558356 455472 558408
rect 463608 558356 463660 558408
rect 472256 558356 472308 558408
rect 481640 558356 481692 558408
rect 75828 558288 75880 558340
rect 80060 558288 80112 558340
rect 88984 558288 89036 558340
rect 98276 558288 98328 558340
rect 107844 558288 107896 558340
rect 162768 558288 162820 558340
rect 198740 558288 198792 558340
rect 213920 558288 213972 558340
rect 223580 558288 223632 558340
rect 225788 558288 225840 558340
rect 234620 558288 234672 558340
rect 339868 558288 339920 558340
rect 349528 558288 349580 558340
rect 357716 558288 357768 558340
rect 359464 558288 359516 558340
rect 456800 558288 456852 558340
rect 465172 558288 465224 558340
rect 474832 558288 474884 558340
rect 477592 558288 477644 558340
rect 478328 558288 478380 558340
rect 487160 558288 487212 558340
rect 78496 558220 78548 558272
rect 87880 558220 87932 558272
rect 91008 558220 91060 558272
rect 99564 558220 99616 558272
rect 108580 558220 108632 558272
rect 161388 558220 161440 558272
rect 197360 558220 197412 558272
rect 216680 558220 216732 558272
rect 217600 558220 217652 558272
rect 226340 558220 226392 558272
rect 227720 558220 227772 558272
rect 237380 558220 237432 558272
rect 291844 558220 291896 558272
rect 329840 558220 329892 558272
rect 334072 558220 334124 558272
rect 343732 558220 343784 558272
rect 346308 558220 346360 558272
rect 354680 558220 354732 558272
rect 359556 558220 359608 558272
rect 458180 558220 458232 558272
rect 467104 558220 467156 558272
rect 488540 558220 488592 558272
rect 64328 558152 64380 558204
rect 193772 558152 193824 558204
rect 313740 558152 313792 558204
rect 443092 558152 443144 558204
rect 443644 558152 443696 558204
rect 459560 558152 459612 558204
rect 465724 558152 465776 558204
rect 487160 558152 487212 558204
rect 128268 558084 128320 558136
rect 195980 558084 196032 558136
rect 204904 558084 204956 558136
rect 213920 558084 213972 558136
rect 290464 558084 290516 558136
rect 331220 558084 331272 558136
rect 349804 558084 349856 558136
rect 452660 558084 452712 558136
rect 454684 558084 454736 558136
rect 464252 558084 464304 558136
rect 464344 558084 464396 558136
rect 485780 558084 485832 558136
rect 80704 558016 80756 558068
rect 82820 558016 82872 558068
rect 100760 558016 100812 558068
rect 101864 558016 101916 558068
rect 198740 558016 198792 558068
rect 206284 558016 206336 558068
rect 215300 558016 215352 558068
rect 322204 558016 322256 558068
rect 328460 558016 328512 558068
rect 329104 558016 329156 558068
rect 337384 558016 337436 558068
rect 352564 558016 352616 558068
rect 476120 558016 476172 558068
rect 100300 557948 100352 558000
rect 197360 557948 197412 558000
rect 209228 557948 209280 558000
rect 216680 557948 216732 558000
rect 327724 557948 327776 558000
rect 336648 557948 336700 558000
rect 352656 557948 352708 558000
rect 477500 557948 477552 558000
rect 71688 557880 71740 557932
rect 78680 557880 78732 557932
rect 202144 557880 202196 557932
rect 211160 557880 211212 557932
rect 322296 557880 322348 557932
rect 331312 557880 331364 557932
rect 352748 557880 352800 557932
rect 478880 557880 478932 557932
rect 70308 557812 70360 557864
rect 77300 557812 77352 557864
rect 93584 557812 93636 557864
rect 102692 557812 102744 557864
rect 201500 557812 201552 557864
rect 203524 557812 203576 557864
rect 212540 557812 212592 557864
rect 302884 557812 302936 557864
rect 322940 557812 322992 557864
rect 323676 557812 323728 557864
rect 332692 557812 332744 557864
rect 353944 557812 353996 557864
rect 480536 557812 480588 557864
rect 66168 557744 66220 557796
rect 74540 557744 74592 557796
rect 106096 557744 106148 557796
rect 205640 557744 205692 557796
rect 287796 557744 287848 557796
rect 317420 557744 317472 557796
rect 324964 557744 325016 557796
rect 334072 557744 334124 557796
rect 356704 557744 356756 557796
rect 483020 557744 483072 557796
rect 67456 557676 67508 557728
rect 75920 557676 75972 557728
rect 107476 557676 107528 557728
rect 207020 557676 207072 557728
rect 207664 557676 207716 557728
rect 216772 557676 216824 557728
rect 286416 557676 286468 557728
rect 320180 557676 320232 557728
rect 326344 557676 326396 557728
rect 335452 557676 335504 557728
rect 354036 557676 354088 557728
rect 481640 557676 481692 557728
rect 63408 557608 63460 557660
rect 73160 557608 73212 557660
rect 104716 557608 104768 557660
rect 202880 557608 202932 557660
rect 209044 557608 209096 557660
rect 218060 557608 218112 557660
rect 329288 557608 329340 557660
rect 338948 557608 339000 557660
rect 358084 557608 358136 557660
rect 454040 557608 454092 557660
rect 456064 557608 456116 557660
rect 465172 557608 465224 557660
rect 468576 557608 468628 557660
rect 477592 557608 477644 557660
rect 62028 557540 62080 557592
rect 71780 557540 71832 557592
rect 74448 557540 74500 557592
rect 78680 557540 78732 557592
rect 210424 557540 210476 557592
rect 220084 557540 220136 557592
rect 227812 557540 227864 557592
rect 330484 557540 330536 557592
rect 339868 557540 339920 557592
rect 450544 557540 450596 557592
rect 451372 557540 451424 557592
rect 457444 557540 457496 557592
rect 466552 557540 466604 557592
rect 474648 557540 474700 557592
rect 474832 557540 474884 557592
rect 483020 557540 483072 557592
rect 58256 556180 58308 556232
rect 579620 556180 579672 556232
rect 169852 553392 169904 553444
rect 170036 553392 170088 553444
rect 57336 545096 57388 545148
rect 580172 545096 580224 545148
rect 56784 543668 56836 543720
rect 146024 543668 146076 543720
rect 206928 543668 206980 543720
rect 220728 543668 220780 543720
rect 229008 543668 229060 543720
rect 260196 543668 260248 543720
rect 56876 543600 56928 543652
rect 148140 543600 148192 543652
rect 205548 543600 205600 543652
rect 218704 543600 218756 543652
rect 227628 543600 227680 543652
rect 258080 543600 258132 543652
rect 61016 543532 61068 543584
rect 62028 543532 62080 543584
rect 56968 543464 57020 543516
rect 150164 543532 150216 543584
rect 164700 543532 164752 543584
rect 165528 543532 165580 543584
rect 177212 543532 177264 543584
rect 177948 543532 178000 543584
rect 208308 543532 208360 543584
rect 222844 543532 222896 543584
rect 231768 543532 231820 543584
rect 264336 543532 264388 543584
rect 57060 543396 57112 543448
rect 152280 543464 152332 543516
rect 160560 543464 160612 543516
rect 161388 543464 161440 543516
rect 193772 543464 193824 543516
rect 209044 543464 209096 543516
rect 209688 543464 209740 543516
rect 224868 543464 224920 543516
rect 230388 543464 230440 543516
rect 262220 543464 262272 543516
rect 57152 543328 57204 543380
rect 154396 543396 154448 543448
rect 195888 543396 195940 543448
rect 210424 543396 210476 543448
rect 210976 543396 211028 543448
rect 226984 543396 227036 543448
rect 233056 543396 233108 543448
rect 266452 543396 266504 543448
rect 57244 543260 57296 543312
rect 156420 543328 156472 543380
rect 189632 543328 189684 543380
rect 207664 543328 207716 543380
rect 212448 543328 212500 543380
rect 231124 543328 231176 543380
rect 233148 543328 233200 543380
rect 268476 543328 268528 543380
rect 65156 543260 65208 543312
rect 66168 543260 66220 543312
rect 73436 543260 73488 543312
rect 74448 543260 74500 543312
rect 77576 543260 77628 543312
rect 79324 543260 79376 543312
rect 79692 543260 79744 543312
rect 80704 543260 80756 543312
rect 80796 543260 80848 543312
rect 168840 543260 168892 543312
rect 191748 543260 191800 543312
rect 209228 543260 209280 543312
rect 211068 543260 211120 543312
rect 229100 543260 229152 543312
rect 234528 543260 234580 543312
rect 270592 543260 270644 543312
rect 70124 543192 70176 543244
rect 170956 543192 171008 543244
rect 187516 543192 187568 543244
rect 206284 543192 206336 543244
rect 213828 543192 213880 543244
rect 233240 543192 233292 543244
rect 235908 543192 235960 543244
rect 272616 543192 272668 543244
rect 70216 543124 70268 543176
rect 173072 543124 173124 543176
rect 185492 543124 185544 543176
rect 204904 543124 204956 543176
rect 216588 543124 216640 543176
rect 237380 543124 237432 543176
rect 238668 543124 238720 543176
rect 276756 543124 276808 543176
rect 71596 543056 71648 543108
rect 175096 543056 175148 543108
rect 183376 543056 183428 543108
rect 203524 543056 203576 543108
rect 215208 543056 215260 543108
rect 235264 543056 235316 543108
rect 237288 543056 237340 543108
rect 274732 543056 274784 543108
rect 56692 542988 56744 543040
rect 179236 542988 179288 543040
rect 181352 542988 181404 543040
rect 202144 542988 202196 543040
rect 202788 542988 202840 543040
rect 214564 542988 214616 543040
rect 217968 542988 218020 543040
rect 239404 542988 239456 543040
rect 240048 542988 240100 543040
rect 278872 542988 278924 543040
rect 67548 542920 67600 542972
rect 144000 542920 144052 542972
rect 204168 542920 204220 542972
rect 216588 542920 216640 542972
rect 226248 542920 226300 542972
rect 256056 542920 256108 542972
rect 68928 542852 68980 542904
rect 80796 542852 80848 542904
rect 91008 542852 91060 542904
rect 92112 542852 92164 542904
rect 92388 542852 92440 542904
rect 94136 542852 94188 542904
rect 100668 542852 100720 542904
rect 108672 542852 108724 542904
rect 108948 542852 109000 542904
rect 123208 542852 123260 542904
rect 127348 542852 127400 542904
rect 128268 542852 128320 542904
rect 129464 542852 129516 542904
rect 188436 542852 188488 542904
rect 226156 542852 226208 542904
rect 253940 542852 253992 542904
rect 93676 542784 93728 542836
rect 96252 542784 96304 542836
rect 99288 542784 99340 542836
rect 106648 542784 106700 542836
rect 110328 542784 110380 542836
rect 125324 542784 125376 542836
rect 131488 542784 131540 542836
rect 188344 542784 188396 542836
rect 223488 542784 223540 542836
rect 249800 542784 249852 542836
rect 93768 542716 93820 542768
rect 98368 542716 98420 542768
rect 107568 542716 107620 542768
rect 121184 542716 121236 542768
rect 139860 542716 139912 542768
rect 140688 542716 140740 542768
rect 140780 542716 140832 542768
rect 159364 542716 159416 542768
rect 224684 542716 224736 542768
rect 251916 542716 251968 542768
rect 69296 542648 69348 542700
rect 70308 542648 70360 542700
rect 96528 542648 96580 542700
rect 102508 542648 102560 542700
rect 83832 542580 83884 542632
rect 85672 542580 85724 542632
rect 97908 542580 97960 542632
rect 104532 542648 104584 542700
rect 106188 542648 106240 542700
rect 119068 542648 119120 542700
rect 135720 542648 135772 542700
rect 160744 542648 160796 542700
rect 220544 542648 220596 542700
rect 245660 542648 245712 542700
rect 103428 542580 103480 542632
rect 114928 542580 114980 542632
rect 222108 542580 222160 542632
rect 247776 542580 247828 542632
rect 81716 542512 81768 542564
rect 84200 542512 84252 542564
rect 104808 542512 104860 542564
rect 117044 542512 117096 542564
rect 133604 542512 133656 542564
rect 140780 542512 140832 542564
rect 217876 542512 217928 542564
rect 241520 542512 241572 542564
rect 95148 542444 95200 542496
rect 100392 542444 100444 542496
rect 101956 542444 102008 542496
rect 112812 542444 112864 542496
rect 219348 542444 219400 542496
rect 243544 542444 243596 542496
rect 102048 542376 102100 542428
rect 110788 542376 110840 542428
rect 211160 540948 211212 541000
rect 211436 540948 211488 541000
rect 56784 540268 56836 540320
rect 137284 540268 137336 540320
rect 56692 540200 56744 540252
rect 170036 540200 170088 540252
rect 56876 539180 56928 539232
rect 299756 539180 299808 539232
rect 59728 539112 59780 539164
rect 429476 539112 429528 539164
rect 59636 539044 59688 539096
rect 559196 539044 559248 539096
rect 57980 538976 58032 539028
rect 580356 538976 580408 539028
rect 58072 538908 58124 538960
rect 580632 538908 580684 538960
rect 57060 538840 57112 538892
rect 580540 538840 580592 538892
rect 2964 538364 3016 538416
rect 5356 538364 5408 538416
rect 60740 538364 60792 538416
rect 541624 538364 541676 538416
rect 60004 538296 60056 538348
rect 563704 538296 563756 538348
rect 19984 538228 20036 538280
rect 57244 538228 57296 538280
rect 58164 538228 58216 538280
rect 579804 538228 579856 538280
rect 57152 537888 57204 537940
rect 580264 537888 580316 537940
rect 48964 536800 49016 536852
rect 57244 536800 57296 536852
rect 60096 536800 60148 536852
rect 60740 536800 60792 536852
rect 282828 536732 282880 536784
rect 467104 536732 467156 536784
rect 282828 535372 282880 535424
rect 465724 535372 465776 535424
rect 4804 534080 4856 534132
rect 57244 534080 57296 534132
rect 282828 532652 282880 532704
rect 464344 532652 464396 532704
rect 53104 531360 53156 531412
rect 57244 531360 57296 531412
rect 282828 531224 282880 531276
rect 356796 531224 356848 531276
rect 541624 530544 541676 530596
rect 556160 530544 556212 530596
rect 563704 530000 563756 530052
rect 46204 529932 46256 529984
rect 57244 529932 57296 529984
rect 569224 529864 569276 529916
rect 556160 529184 556212 529236
rect 568488 529184 568540 529236
rect 282828 528504 282880 528556
rect 356704 528504 356756 528556
rect 4896 527144 4948 527196
rect 57244 527144 57296 527196
rect 17224 525784 17276 525836
rect 57244 525784 57296 525836
rect 568488 525784 568540 525836
rect 282828 525716 282880 525768
rect 355324 525716 355376 525768
rect 571984 525716 572036 525768
rect 282828 524356 282880 524408
rect 354036 524356 354088 524408
rect 43444 522996 43496 523048
rect 57244 522996 57296 523048
rect 4988 521636 5040 521688
rect 57244 521636 57296 521688
rect 282828 521568 282880 521620
rect 353944 521568 353996 521620
rect 569224 521568 569276 521620
rect 570972 521568 571024 521620
rect 282828 520208 282880 520260
rect 352748 520208 352800 520260
rect 51724 518916 51776 518968
rect 57244 518916 57296 518968
rect 35164 517488 35216 517540
rect 57244 517488 57296 517540
rect 570972 517488 571024 517540
rect 281908 517420 281960 517472
rect 352656 517420 352708 517472
rect 573364 517420 573416 517472
rect 3424 514768 3476 514820
rect 57244 514768 57296 514820
rect 282828 514700 282880 514752
rect 352564 514700 352616 514752
rect 50344 513340 50396 513392
rect 57244 513340 57296 513392
rect 282092 513272 282144 513324
rect 476212 513272 476264 513324
rect 571984 513272 572036 513324
rect 574744 513272 574796 513324
rect 33784 510620 33836 510672
rect 57244 510620 57296 510672
rect 282828 510552 282880 510604
rect 474740 510552 474792 510604
rect 2780 509532 2832 509584
rect 5448 509532 5500 509584
rect 3516 509260 3568 509312
rect 57244 509260 57296 509312
rect 282276 509192 282328 509244
rect 473360 509192 473412 509244
rect 574744 507764 574796 507816
rect 577964 507764 578016 507816
rect 39396 506472 39448 506524
rect 57244 506472 57296 506524
rect 281908 506404 281960 506456
rect 471980 506404 472032 506456
rect 577964 506268 578016 506320
rect 580264 506268 580316 506320
rect 28264 505112 28316 505164
rect 57244 505112 57296 505164
rect 282828 503616 282880 503668
rect 470600 503616 470652 503668
rect 3608 502324 3660 502376
rect 57244 502324 57296 502376
rect 282092 502256 282144 502308
rect 469220 502256 469272 502308
rect 37924 500964 37976 501016
rect 57244 500964 57296 501016
rect 573364 499536 573416 499588
rect 282828 499468 282880 499520
rect 467932 499468 467984 499520
rect 576768 499468 576820 499520
rect 20076 498176 20128 498228
rect 57244 498176 57296 498228
rect 282276 498108 282328 498160
rect 467840 498108 467892 498160
rect 281908 495388 281960 495440
rect 466460 495388 466512 495440
rect 32404 494028 32456 494080
rect 57244 494028 57296 494080
rect 282460 493960 282512 494012
rect 465080 493960 465132 494012
rect 576860 493824 576912 493876
rect 578884 493824 578936 493876
rect 17316 491308 17368 491360
rect 57244 491308 57296 491360
rect 282092 491240 282144 491292
rect 463700 491240 463752 491292
rect 56968 491172 57020 491224
rect 57244 491172 57296 491224
rect 282828 488452 282880 488504
rect 462320 488452 462372 488504
rect 3700 487160 3752 487212
rect 56600 487160 56652 487212
rect 282828 487092 282880 487144
rect 461032 487092 461084 487144
rect 15844 485800 15896 485852
rect 56600 485800 56652 485852
rect 282828 484304 282880 484356
rect 460940 484304 460992 484356
rect 3792 483012 3844 483064
rect 56600 483012 56652 483064
rect 282460 482944 282512 482996
rect 443644 482944 443696 482996
rect 4068 481652 4120 481704
rect 56600 481652 56652 481704
rect 3240 480632 3292 480684
rect 5540 480632 5592 480684
rect 282092 480156 282144 480208
rect 359556 480156 359608 480208
rect 3976 478864 4028 478916
rect 56600 478864 56652 478916
rect 282828 477436 282880 477488
rect 359464 477436 359516 477488
rect 3332 476008 3384 476060
rect 56600 476008 56652 476060
rect 282552 476008 282604 476060
rect 358176 476008 358228 476060
rect 5540 474648 5592 474700
rect 56600 474648 56652 474700
rect 282092 473288 282144 473340
rect 358084 473288 358136 473340
rect 5448 471928 5500 471980
rect 56600 471928 56652 471980
rect 282460 471928 282512 471980
rect 349804 471928 349856 471980
rect 3884 470500 3936 470552
rect 56508 470500 56560 470552
rect 282092 469140 282144 469192
rect 452752 469140 452804 469192
rect 5356 467780 5408 467832
rect 56508 467780 56560 467832
rect 5264 466352 5316 466404
rect 56508 466352 56560 466404
rect 282828 466352 282880 466404
rect 330484 466352 330536 466404
rect 282276 464992 282328 465044
rect 329288 464992 329340 465044
rect 31024 463632 31076 463684
rect 56508 463632 56560 463684
rect 14464 462272 14516 462324
rect 56508 462272 56560 462324
rect 282828 462272 282880 462324
rect 329104 462272 329156 462324
rect 576860 462000 576912 462052
rect 579988 462000 580040 462052
rect 282460 460844 282512 460896
rect 327724 460844 327776 460896
rect 571800 459552 571852 459604
rect 576860 459552 576912 459604
rect 5172 459484 5224 459536
rect 56600 459484 56652 459536
rect 282092 458124 282144 458176
rect 326344 458124 326396 458176
rect 21364 456696 21416 456748
rect 56600 456696 56652 456748
rect 566464 456016 566516 456068
rect 571800 456016 571852 456068
rect 13084 455336 13136 455388
rect 56600 455336 56652 455388
rect 282828 455336 282880 455388
rect 324964 455336 325016 455388
rect 282828 453976 282880 454028
rect 323676 453976 323728 454028
rect 5080 452480 5132 452532
rect 56600 452480 56652 452532
rect 3332 452344 3384 452396
rect 56508 452344 56560 452396
rect 24768 451188 24820 451240
rect 56600 451188 56652 451240
rect 282828 451188 282880 451240
rect 322296 451188 322348 451240
rect 282460 449828 282512 449880
rect 460388 449828 460440 449880
rect 56600 448604 56652 448656
rect 57520 448604 57572 448656
rect 10324 448468 10376 448520
rect 57520 448468 57572 448520
rect 42064 447040 42116 447092
rect 57520 447040 57572 447092
rect 282828 447040 282880 447092
rect 460204 447040 460256 447092
rect 563244 445680 563296 445732
rect 566464 445748 566516 445800
rect 282828 444320 282880 444372
rect 458824 444320 458876 444372
rect 282828 442892 282880 442944
rect 457444 442892 457496 442944
rect 562416 442144 562468 442196
rect 563244 442144 563296 442196
rect 578608 440240 578660 440292
rect 580264 440240 580316 440292
rect 282828 440172 282880 440224
rect 456064 440172 456116 440224
rect 560944 438880 560996 438932
rect 562416 438880 562468 438932
rect 576124 438880 576176 438932
rect 578608 438880 578660 438932
rect 282460 438812 282512 438864
rect 454684 438812 454736 438864
rect 577964 437588 578016 437640
rect 579620 437588 579672 437640
rect 282828 436024 282880 436076
rect 453488 436024 453540 436076
rect 575848 435480 575900 435532
rect 577964 435480 578016 435532
rect 57612 433984 57664 434036
rect 60096 433984 60148 434036
rect 282828 433236 282880 433288
rect 453304 433236 453356 433288
rect 574744 432488 574796 432540
rect 575848 432488 575900 432540
rect 282828 431876 282880 431928
rect 291936 431876 291988 431928
rect 58716 429156 58768 429208
rect 60004 429156 60056 429208
rect 282828 429088 282880 429140
rect 290556 429088 290608 429140
rect 570604 426776 570656 426828
rect 576124 426776 576176 426828
rect 282828 426572 282880 426624
rect 287704 426572 287756 426624
rect 282460 425008 282512 425060
rect 286324 425008 286376 425060
rect 570788 422696 570840 422748
rect 574744 422696 574796 422748
rect 282092 422220 282144 422272
rect 284944 422220 284996 422272
rect 281724 420792 281776 420844
rect 283564 420792 283616 420844
rect 567844 419500 567896 419552
rect 570788 419500 570840 419552
rect 558184 418140 558236 418192
rect 560944 418140 560996 418192
rect 282828 418072 282880 418124
rect 294604 418072 294656 418124
rect 282828 416712 282880 416764
rect 316040 416712 316092 416764
rect 57704 413924 57756 413976
rect 58716 413924 58768 413976
rect 281908 413924 281960 413976
rect 399484 413924 399536 413976
rect 282828 411204 282880 411256
rect 398104 411204 398156 411256
rect 282092 409776 282144 409828
rect 395344 409776 395396 409828
rect 282828 407056 282880 407108
rect 393964 407056 394016 407108
rect 578976 405696 579028 405748
rect 580264 405696 580316 405748
rect 282828 405628 282880 405680
rect 392584 405628 392636 405680
rect 577596 403520 577648 403572
rect 578976 403520 579028 403572
rect 281908 402908 281960 402960
rect 391204 402908 391256 402960
rect 577504 400188 577556 400240
rect 580908 400188 580960 400240
rect 282828 400120 282880 400172
rect 388444 400120 388496 400172
rect 556804 399644 556856 399696
rect 558184 399644 558236 399696
rect 282092 398760 282144 398812
rect 445760 398760 445812 398812
rect 282092 395836 282144 395888
rect 285036 395836 285088 395888
rect 282276 394612 282328 394664
rect 402244 394612 402296 394664
rect 569224 394612 569276 394664
rect 570604 394612 570656 394664
rect 566556 391960 566608 392012
rect 567844 391960 567896 392012
rect 577872 391960 577924 392012
rect 579620 391960 579672 392012
rect 281908 391892 281960 391944
rect 320272 391892 320324 391944
rect 574100 390600 574152 390652
rect 577596 390600 577648 390652
rect 282460 389784 282512 389836
rect 286416 389784 286468 389836
rect 282092 387744 282144 387796
rect 318800 387744 318852 387796
rect 555424 387744 555476 387796
rect 556804 387744 556856 387796
rect 571984 387132 572036 387184
rect 574100 387132 574152 387184
rect 576216 385024 576268 385076
rect 577872 385024 577924 385076
rect 282828 384616 282880 384668
rect 287796 384616 287848 384668
rect 282828 383596 282880 383648
rect 450544 383596 450596 383648
rect 567384 382236 567436 382288
rect 571984 382236 572036 382288
rect 574100 382236 574152 382288
rect 576216 382236 576268 382288
rect 282828 380808 282880 380860
rect 449164 380808 449216 380860
rect 282460 379448 282512 379500
rect 447784 379448 447836 379500
rect 566648 377680 566700 377732
rect 567384 377680 567436 377732
rect 282092 376660 282144 376712
rect 446404 376660 446456 376712
rect 570972 376320 571024 376372
rect 574100 376320 574152 376372
rect 282828 373940 282880 373992
rect 358820 373940 358872 373992
rect 282552 372512 282604 372564
rect 357440 372512 357492 372564
rect 566464 371696 566516 371748
rect 569224 371696 569276 371748
rect 568764 371560 568816 371612
rect 570972 371560 571024 371612
rect 565268 369860 565320 369912
rect 566648 369860 566700 369912
rect 282828 369792 282880 369844
rect 356060 369792 356112 369844
rect 564072 369792 564124 369844
rect 568764 369860 568816 369912
rect 282460 368432 282512 368484
rect 354772 368432 354824 368484
rect 563704 368432 563756 368484
rect 566556 368432 566608 368484
rect 563796 368024 563848 368076
rect 565268 368024 565320 368076
rect 560944 367072 560996 367124
rect 564072 367072 564124 367124
rect 577596 367072 577648 367124
rect 579528 367072 579580 367124
rect 2964 367004 3016 367056
rect 15844 367004 15896 367056
rect 282092 365644 282144 365696
rect 353300 365644 353352 365696
rect 282828 362856 282880 362908
rect 352012 362856 352064 362908
rect 282552 361496 282604 361548
rect 352196 361496 352248 361548
rect 553308 360816 553360 360868
rect 563796 360816 563848 360868
rect 282828 358708 282880 358760
rect 350540 358708 350592 358760
rect 282460 357348 282512 357400
rect 349160 357348 349212 357400
rect 562416 357008 562468 357060
rect 563704 357008 563756 357060
rect 551284 356600 551336 356652
rect 553308 356600 553360 356652
rect 576860 356056 576912 356108
rect 579528 356056 579580 356108
rect 574744 354696 574796 354748
rect 577504 354696 577556 354748
rect 282092 354628 282144 354680
rect 347780 354628 347832 354680
rect 571984 353404 572036 353456
rect 576860 353404 576912 353456
rect 549260 351908 549312 351960
rect 551284 351908 551336 351960
rect 554044 351908 554096 351960
rect 555424 351908 555476 351960
rect 282828 351840 282880 351892
rect 346400 351840 346452 351892
rect 561036 350548 561088 350600
rect 562416 350548 562468 350600
rect 282552 350480 282604 350532
rect 345020 350480 345072 350532
rect 564440 349800 564492 349852
rect 571984 349800 572036 349852
rect 559564 348372 559616 348424
rect 560944 348372 560996 348424
rect 282828 347692 282880 347744
rect 343732 347692 343784 347744
rect 561680 347420 561732 347472
rect 564440 347420 564492 347472
rect 573364 347420 573416 347472
rect 574744 347420 574796 347472
rect 282460 346332 282512 346384
rect 343640 346332 343692 346384
rect 548524 345856 548576 345908
rect 549260 345856 549312 345908
rect 574100 345040 574152 345092
rect 577596 345040 577648 345092
rect 559656 343612 559708 343664
rect 561036 343612 561088 343664
rect 282828 343544 282880 343596
rect 342260 343544 342312 343596
rect 558460 343544 558512 343596
rect 561680 343612 561732 343664
rect 552664 342252 552716 342304
rect 554044 342252 554096 342304
rect 553400 340892 553452 340944
rect 558460 340892 558512 340944
rect 571432 340892 571484 340944
rect 574100 340892 574152 340944
rect 282828 340824 282880 340876
rect 340880 340824 340932 340876
rect 578884 340144 578936 340196
rect 580172 340144 580224 340196
rect 57060 339396 57112 339448
rect 58716 339396 58768 339448
rect 282828 339396 282880 339448
rect 339500 339396 339552 339448
rect 563428 338648 563480 338700
rect 566464 338648 566516 338700
rect 551376 338104 551428 338156
rect 553400 338104 553452 338156
rect 3332 338036 3384 338088
rect 56968 338036 57020 338088
rect 57704 336676 57756 336728
rect 58624 336676 58676 336728
rect 282828 336676 282880 336728
rect 338120 336676 338172 336728
rect 561772 336608 561824 336660
rect 563428 336608 563480 336660
rect 570972 336336 571024 336388
rect 571432 336336 571484 336388
rect 282368 335248 282420 335300
rect 336832 335248 336884 335300
rect 551284 333956 551336 334008
rect 552664 333956 552716 334008
rect 558828 333956 558880 334008
rect 561772 333956 561824 334008
rect 282828 332528 282880 332580
rect 336740 332528 336792 332580
rect 57152 331576 57204 331628
rect 58808 331576 58860 331628
rect 556804 331440 556856 331492
rect 558828 331440 558880 331492
rect 567844 331304 567896 331356
rect 570972 331304 571024 331356
rect 546500 331168 546552 331220
rect 548524 331168 548576 331220
rect 57336 330488 57388 330540
rect 57704 330488 57756 330540
rect 565084 330080 565136 330132
rect 567844 330080 567896 330132
rect 282828 329740 282880 329792
rect 335360 329740 335412 329792
rect 57428 328380 57480 328432
rect 58900 328380 58952 328432
rect 282828 328380 282880 328432
rect 333980 328380 334032 328432
rect 576860 328380 576912 328432
rect 578884 328380 578936 328432
rect 549352 328108 549404 328160
rect 551376 328108 551428 328160
rect 549260 327700 549312 327752
rect 559656 327700 559708 327752
rect 57704 327020 57756 327072
rect 58992 327020 59044 327072
rect 282828 325592 282880 325644
rect 332600 325592 332652 325644
rect 543740 325592 543792 325644
rect 546500 325660 546552 325712
rect 552664 325320 552716 325372
rect 559564 325320 559616 325372
rect 545120 324300 545172 324352
rect 549352 324300 549404 324352
rect 553400 324300 553452 324352
rect 556804 324300 556856 324352
rect 3056 324232 3108 324284
rect 32404 324232 32456 324284
rect 282368 324232 282420 324284
rect 290464 324232 290516 324284
rect 535460 323552 535512 323604
rect 543740 323552 543792 323604
rect 57796 322940 57848 322992
rect 59084 322940 59136 322992
rect 549168 322940 549220 322992
rect 552664 322940 552716 322992
rect 57612 322056 57664 322108
rect 59268 322056 59320 322108
rect 532884 321580 532936 321632
rect 535460 321580 535512 321632
rect 282828 321512 282880 321564
rect 329932 321512 329984 321564
rect 544108 321444 544160 321496
rect 549260 321580 549312 321632
rect 548524 320696 548576 320748
rect 551284 320696 551336 320748
rect 543004 320152 543056 320204
rect 545120 320152 545172 320204
rect 56600 320084 56652 320136
rect 58532 320084 58584 320136
rect 546500 319744 546552 319796
rect 549168 319744 549220 319796
rect 549904 319472 549956 319524
rect 553400 319472 553452 319524
rect 529572 319200 529624 319252
rect 532884 319200 532936 319252
rect 574836 318792 574888 318844
rect 576768 318792 576820 318844
rect 282828 318724 282880 318776
rect 291844 318724 291896 318776
rect 57796 317840 57848 317892
rect 57520 317364 57572 317416
rect 58440 317364 58492 317416
rect 282828 317364 282880 317416
rect 322204 317364 322256 317416
rect 57520 317228 57572 317280
rect 572720 317024 572772 317076
rect 574836 317024 574888 317076
rect 542084 316956 542136 317008
rect 544108 316956 544160 317008
rect 545212 316616 545264 316668
rect 546500 316616 546552 316668
rect 56600 315936 56652 315988
rect 57520 315936 57572 315988
rect 523500 315936 523552 315988
rect 529572 316004 529624 316056
rect 57704 315800 57756 315852
rect 57980 315800 58032 315852
rect 59084 314644 59136 314696
rect 60004 314644 60056 314696
rect 560944 314644 560996 314696
rect 565084 314644 565136 314696
rect 282828 314576 282880 314628
rect 327080 314576 327132 314628
rect 282368 313216 282420 313268
rect 325700 313216 325752 313268
rect 539968 311924 540020 311976
rect 542084 311924 542136 311976
rect 543096 311788 543148 311840
rect 545212 311856 545264 311908
rect 567936 311788 567988 311840
rect 573364 311856 573416 311908
rect 535460 311108 535512 311160
rect 543004 311108 543056 311160
rect 545120 310972 545172 311024
rect 549904 310972 549956 311024
rect 281908 310428 281960 310480
rect 323584 310428 323636 310480
rect 563060 309952 563112 310004
rect 567936 309952 567988 310004
rect 519544 309748 519596 309800
rect 539968 309748 540020 309800
rect 3332 309068 3384 309120
rect 17316 309068 17368 309120
rect 532332 309068 532384 309120
rect 535460 309136 535512 309188
rect 569960 309136 570012 309188
rect 572720 309136 572772 309188
rect 539692 308660 539744 308712
rect 545120 308660 545172 308712
rect 565084 308388 565136 308440
rect 569960 308388 570012 308440
rect 282828 307708 282880 307760
rect 302884 307708 302936 307760
rect 557540 307708 557592 307760
rect 563060 307776 563112 307828
rect 522488 307096 522540 307148
rect 523500 307096 523552 307148
rect 56508 306348 56560 306400
rect 57520 306348 57572 306400
rect 57612 306348 57664 306400
rect 57980 306348 58032 306400
rect 282092 306280 282144 306332
rect 321560 306280 321612 306332
rect 517520 305600 517572 305652
rect 522488 305600 522540 305652
rect 516140 304988 516192 305040
rect 519544 304988 519596 305040
rect 540980 304988 541032 305040
rect 543096 304988 543148 305040
rect 546500 304988 546552 305040
rect 548524 304988 548576 305040
rect 59268 304444 59320 304496
rect 59452 304444 59504 304496
rect 58716 304308 58768 304360
rect 59544 304308 59596 304360
rect 58808 303424 58860 303476
rect 60648 303424 60700 303476
rect 553400 302744 553452 302796
rect 557540 302744 557592 302796
rect 559104 302336 559156 302388
rect 560944 302336 560996 302388
rect 536840 300976 536892 301028
rect 539692 300976 539744 301028
rect 514760 300840 514812 300892
rect 517520 300840 517572 300892
rect 57888 300772 57940 300824
rect 580264 300772 580316 300824
rect 56692 300704 56744 300756
rect 580356 300704 580408 300756
rect 59452 300636 59504 300688
rect 565084 300636 565136 300688
rect 60004 300568 60056 300620
rect 559104 300568 559156 300620
rect 60648 300500 60700 300552
rect 553400 300500 553452 300552
rect 58624 300432 58676 300484
rect 546500 300432 546552 300484
rect 58440 300364 58492 300416
rect 540888 300364 540940 300416
rect 59544 300296 59596 300348
rect 536840 300296 536892 300348
rect 58992 300228 59044 300280
rect 532332 300228 532384 300280
rect 58900 300160 58952 300212
rect 516140 300160 516192 300212
rect 58532 300092 58584 300144
rect 514760 300092 514812 300144
rect 56784 299412 56836 299464
rect 579804 299412 579856 299464
rect 39304 298052 39356 298104
rect 68652 298052 68704 298104
rect 82728 298052 82780 298104
rect 193220 298052 193272 298104
rect 32404 297984 32456 298036
rect 78404 297984 78456 298036
rect 86868 297984 86920 298036
rect 201040 297984 201092 298036
rect 4068 297916 4120 297968
rect 64788 297916 64840 297968
rect 89628 297916 89680 297968
rect 204904 297916 204956 297968
rect 10968 297848 11020 297900
rect 76472 297848 76524 297900
rect 96528 297848 96580 297900
rect 216588 297848 216640 297900
rect 16488 297780 16540 297832
rect 86224 297780 86276 297832
rect 93768 297780 93820 297832
rect 212724 297780 212776 297832
rect 42708 297712 42760 297764
rect 129004 297712 129056 297764
rect 134524 297712 134576 297764
rect 255504 297712 255556 297764
rect 15108 297644 15160 297696
rect 84200 297644 84252 297696
rect 100668 297644 100720 297696
rect 224408 297644 224460 297696
rect 20628 297576 20680 297628
rect 92020 297576 92072 297628
rect 103428 297576 103480 297628
rect 228272 297576 228324 297628
rect 21916 297508 21968 297560
rect 93952 297508 94004 297560
rect 107568 297508 107620 297560
rect 234160 297508 234212 297560
rect 24768 297440 24820 297492
rect 99840 297440 99892 297492
rect 107476 297440 107528 297492
rect 236092 297440 236144 297492
rect 26148 297372 26200 297424
rect 101772 297372 101824 297424
rect 114468 297372 114520 297424
rect 245844 297372 245896 297424
rect 51816 297304 51868 297356
rect 70584 297304 70636 297356
rect 79968 297304 80020 297356
rect 189356 297304 189408 297356
rect 74448 297236 74500 297288
rect 181536 297236 181588 297288
rect 72976 297168 73028 297220
rect 177672 297168 177724 297220
rect 67548 297100 67600 297152
rect 169852 297100 169904 297152
rect 64788 297032 64840 297084
rect 165988 297032 166040 297084
rect 62028 296964 62080 297016
rect 160192 296964 160244 297016
rect 50988 296896 51040 296948
rect 142620 296896 142672 296948
rect 48136 296828 48188 296880
rect 136824 296828 136876 296880
rect 39948 296760 40000 296812
rect 124772 296760 124824 296812
rect 124864 296760 124916 296812
rect 146576 296760 146628 296812
rect 42064 296692 42116 296744
rect 107292 296692 107344 296744
rect 56692 296624 56744 296676
rect 57336 296624 57388 296676
rect 57520 296624 57572 296676
rect 57888 296624 57940 296676
rect 2964 295264 3016 295316
rect 57244 295264 57296 295316
rect 61016 292544 61068 292596
rect 61108 292476 61160 292528
rect 61016 288396 61068 288448
rect 61108 288396 61160 288448
rect 56784 287104 56836 287156
rect 57612 287104 57664 287156
rect 56692 287036 56744 287088
rect 57336 287036 57388 287088
rect 57520 287036 57572 287088
rect 57888 287036 57940 287088
rect 67548 280372 67600 280424
rect 67548 280236 67600 280288
rect 3332 280100 3384 280152
rect 37924 280100 37976 280152
rect 57244 277312 57296 277364
rect 57520 277312 57572 277364
rect 57612 277312 57664 277364
rect 57888 277312 57940 277364
rect 56876 275952 56928 276004
rect 580172 275952 580224 276004
rect 60740 273232 60792 273284
rect 61108 273232 61160 273284
rect 56784 268404 56836 268456
rect 57336 268404 57388 268456
rect 57612 268404 57664 268456
rect 57888 268404 57940 268456
rect 3148 266296 3200 266348
rect 20076 266296 20128 266348
rect 56968 264868 57020 264920
rect 580172 264868 580224 264920
rect 57244 263576 57296 263628
rect 57520 263576 57572 263628
rect 60924 263508 60976 263560
rect 61108 263508 61160 263560
rect 60832 260788 60884 260840
rect 61108 260788 61160 260840
rect 57060 252492 57112 252544
rect 579804 252492 579856 252544
rect 60832 251200 60884 251252
rect 61016 251200 61068 251252
rect 3240 237328 3292 237380
rect 39396 237328 39448 237380
rect 67364 231820 67416 231872
rect 67364 231684 67416 231736
rect 67272 230392 67324 230444
rect 67364 230392 67416 230444
rect 57152 229032 57204 229084
rect 580172 229032 580224 229084
rect 60740 224952 60792 225004
rect 60924 224816 60976 224868
rect 3332 223524 3384 223576
rect 28264 223524 28316 223576
rect 67272 220804 67324 220856
rect 67548 220804 67600 220856
rect 57336 217948 57388 218000
rect 580172 217948 580224 218000
rect 60740 215296 60792 215348
rect 60924 215296 60976 215348
rect 67548 212508 67600 212560
rect 67456 212440 67508 212492
rect 67456 211080 67508 211132
rect 67548 211080 67600 211132
rect 57428 205572 57480 205624
rect 579804 205572 579856 205624
rect 60648 205504 60700 205556
rect 60924 205504 60976 205556
rect 67548 202852 67600 202904
rect 67456 202784 67508 202836
rect 60924 195984 60976 196036
rect 61016 195916 61068 195968
rect 3516 194488 3568 194540
rect 50344 194488 50396 194540
rect 57520 182112 57572 182164
rect 580172 182112 580224 182164
rect 60924 181500 60976 181552
rect 61108 181500 61160 181552
rect 3240 180752 3292 180804
rect 33784 180752 33836 180804
rect 57612 171028 57664 171080
rect 580172 171028 580224 171080
rect 60924 166948 60976 167000
rect 61108 166948 61160 167000
rect 59360 158652 59412 158704
rect 579804 158652 579856 158704
rect 61200 157428 61252 157480
rect 61016 157224 61068 157276
rect 61016 153144 61068 153196
rect 61200 153144 61252 153196
rect 3148 151716 3200 151768
rect 51724 151716 51776 151768
rect 60924 137980 60976 138032
rect 61016 137912 61068 137964
rect 3240 136552 3292 136604
rect 35164 136552 35216 136604
rect 57704 135192 57756 135244
rect 580172 135192 580224 135244
rect 57796 124108 57848 124160
rect 580172 124108 580224 124160
rect 2780 122272 2832 122324
rect 4988 122272 5040 122324
rect 60924 118668 60976 118720
rect 61016 118600 61068 118652
rect 67456 115880 67508 115932
rect 67548 115880 67600 115932
rect 67272 114452 67324 114504
rect 67456 114452 67508 114504
rect 59084 111732 59136 111784
rect 579804 111732 579856 111784
rect 3240 108944 3292 108996
rect 17224 108944 17276 108996
rect 67272 104864 67324 104916
rect 67548 104864 67600 104916
rect 60740 99356 60792 99408
rect 61108 99220 61160 99272
rect 3424 93780 3476 93832
rect 43444 93780 43496 93832
rect 56600 88272 56652 88324
rect 580172 88272 580224 88324
rect 60740 86912 60792 86964
rect 61016 86912 61068 86964
rect 2780 79772 2832 79824
rect 4896 79772 4948 79824
rect 60740 77256 60792 77308
rect 60924 77256 60976 77308
rect 89536 76100 89588 76152
rect 89812 76100 89864 76152
rect 147588 76100 147640 76152
rect 154488 76100 154540 76152
rect 115940 75964 115992 76016
rect 118884 75964 118936 76016
rect 60648 75828 60700 75880
rect 60924 75828 60976 75880
rect 3332 64812 3384 64864
rect 53104 64812 53156 64864
rect 59176 64812 59228 64864
rect 579804 64812 579856 64864
rect 60924 60664 60976 60716
rect 61108 60664 61160 60716
rect 60832 57876 60884 57928
rect 61108 57876 61160 57928
rect 67456 57876 67508 57928
rect 67548 57876 67600 57928
rect 67272 56516 67324 56568
rect 67456 56516 67508 56568
rect 3424 51008 3476 51060
rect 46204 51008 46256 51060
rect 60832 48288 60884 48340
rect 61016 48288 61068 48340
rect 67272 46928 67324 46980
rect 67548 46928 67600 46980
rect 147588 40196 147640 40248
rect 154488 40196 154540 40248
rect 89536 40128 89588 40180
rect 91744 40128 91796 40180
rect 115940 40060 115992 40112
rect 118884 40060 118936 40112
rect 67456 37272 67508 37324
rect 67548 37272 67600 37324
rect 2780 35844 2832 35896
rect 4804 35844 4856 35896
rect 60924 31832 60976 31884
rect 60924 31696 60976 31748
rect 86868 29248 86920 29300
rect 147588 29180 147640 29232
rect 154488 29180 154540 29232
rect 86868 29112 86920 29164
rect 115940 29044 115992 29096
rect 120816 29044 120868 29096
rect 67548 27616 67600 27668
rect 67732 27616 67784 27668
rect 2872 22040 2924 22092
rect 19984 22040 20036 22092
rect 67548 19252 67600 19304
rect 66996 19184 67048 19236
rect 59268 17892 59320 17944
rect 579804 17892 579856 17944
rect 60740 12452 60792 12504
rect 60832 12316 60884 12368
rect 59176 9596 59228 9648
rect 60832 9596 60884 9648
rect 3424 8236 3476 8288
rect 48964 8236 49016 8288
rect 60004 6400 60056 6452
rect 157340 6400 157392 6452
rect 108764 6332 108816 6384
rect 237380 6332 237432 6384
rect 112352 6264 112404 6316
rect 242900 6264 242952 6316
rect 115940 6196 115992 6248
rect 248420 6196 248472 6248
rect 123024 6128 123076 6180
rect 260840 6128 260892 6180
rect 93860 5516 93912 5568
rect 99472 5516 99524 5568
rect 108948 5516 109000 5568
rect 109040 5516 109092 5568
rect 7656 5448 7708 5500
rect 71780 5448 71832 5500
rect 71872 5448 71924 5500
rect 12440 5380 12492 5432
rect 80060 5380 80112 5432
rect 80244 5448 80296 5500
rect 190460 5448 190512 5500
rect 83740 5380 83792 5432
rect 83832 5380 83884 5432
rect 195980 5380 196032 5432
rect 17224 5312 17276 5364
rect 86960 5312 87012 5364
rect 87328 5312 87380 5364
rect 202880 5312 202932 5364
rect 65524 5244 65576 5296
rect 71872 5244 71924 5296
rect 84108 5244 84160 5296
rect 93860 5244 93912 5296
rect 22008 5176 22060 5228
rect 95240 5176 95292 5228
rect 98092 5176 98144 5228
rect 108948 5244 109000 5296
rect 109040 5244 109092 5296
rect 219440 5244 219492 5296
rect 99472 5176 99524 5228
rect 26700 5108 26752 5160
rect 103520 5108 103572 5160
rect 105176 5176 105228 5228
rect 231860 5176 231912 5228
rect 124864 5108 124916 5160
rect 127808 5108 127860 5160
rect 137376 5108 137428 5160
rect 137652 5108 137704 5160
rect 266360 5108 266412 5160
rect 30288 5040 30340 5092
rect 109132 5040 109184 5092
rect 119436 5040 119488 5092
rect 134524 5040 134576 5092
rect 134616 5040 134668 5092
rect 137192 5040 137244 5092
rect 33876 4972 33928 5024
rect 114560 4972 114612 5024
rect 130200 4972 130252 5024
rect 271880 5040 271932 5092
rect 137468 4972 137520 5024
rect 269120 4972 269172 5024
rect 37372 4904 37424 4956
rect 120080 4904 120132 4956
rect 126612 4904 126664 4956
rect 40960 4836 41012 4888
rect 126980 4836 127032 4888
rect 129004 4904 129056 4956
rect 270500 4904 270552 4956
rect 137468 4836 137520 4888
rect 137560 4836 137612 4888
rect 276020 4836 276072 4888
rect 44548 4768 44600 4820
rect 132500 4768 132552 4820
rect 132592 4768 132644 4820
rect 134616 4768 134668 4820
rect 134892 4768 134944 4820
rect 278780 4768 278832 4820
rect 52828 4700 52880 4752
rect 65524 4700 65576 4752
rect 76656 4700 76708 4752
rect 184940 4700 184992 4752
rect 73068 4632 73120 4684
rect 179420 4632 179472 4684
rect 69480 4564 69532 4616
rect 172520 4564 172572 4616
rect 65984 4496 66036 4548
rect 167000 4496 167052 4548
rect 62396 4428 62448 4480
rect 161480 4428 161532 4480
rect 58808 4360 58860 4412
rect 155960 4360 156012 4412
rect 55220 4292 55272 4344
rect 150440 4292 150492 4344
rect 51632 4224 51684 4276
rect 143540 4224 143592 4276
rect 48228 4156 48280 4208
rect 138020 4156 138072 4208
rect 3976 4088 4028 4140
rect 61108 4088 61160 4140
rect 61200 4088 61252 4140
rect 62028 4088 62080 4140
rect 68284 4088 68336 4140
rect 73344 4088 73396 4140
rect 8852 4020 8904 4072
rect 74540 4020 74592 4072
rect 13636 3952 13688 4004
rect 81440 4088 81492 4140
rect 77852 4020 77904 4072
rect 82636 4020 82688 4072
rect 83004 4088 83056 4140
rect 183560 4088 183612 4140
rect 75460 3952 75512 4004
rect 78956 3952 79008 4004
rect 79048 3952 79100 4004
rect 79968 3952 80020 4004
rect 81440 3952 81492 4004
rect 82728 3952 82780 4004
rect 186320 4020 186372 4072
rect 194600 3952 194652 4004
rect 18328 3884 18380 3936
rect 86040 3884 86092 3936
rect 86132 3884 86184 3936
rect 86868 3884 86920 3936
rect 88524 3884 88576 3936
rect 89628 3884 89680 3936
rect 89720 3884 89772 3936
rect 93216 3884 93268 3936
rect 93308 3884 93360 3936
rect 93768 3884 93820 3936
rect 93860 3884 93912 3936
rect 205640 3884 205692 3936
rect 24308 3816 24360 3868
rect 24768 3816 24820 3868
rect 25504 3816 25556 3868
rect 26148 3816 26200 3868
rect 23112 3748 23164 3800
rect 95516 3816 95568 3868
rect 27896 3748 27948 3800
rect 95700 3748 95752 3800
rect 96528 3748 96580 3800
rect 96896 3816 96948 3868
rect 218060 3816 218112 3868
rect 102692 3748 102744 3800
rect 102784 3748 102836 3800
rect 103428 3748 103480 3800
rect 106372 3748 106424 3800
rect 107568 3748 107620 3800
rect 107660 3748 107712 3800
rect 113180 3748 113232 3800
rect 113548 3748 113600 3800
rect 114468 3748 114520 3800
rect 114744 3748 114796 3800
rect 115848 3748 115900 3800
rect 31484 3680 31536 3732
rect 110420 3680 110472 3732
rect 34980 3612 35032 3664
rect 109868 3612 109920 3664
rect 109960 3612 110012 3664
rect 238760 3748 238812 3800
rect 32680 3544 32732 3596
rect 107660 3544 107712 3596
rect 111156 3544 111208 3596
rect 241520 3680 241572 3732
rect 117136 3612 117188 3664
rect 118240 3544 118292 3596
rect 120632 3612 120684 3664
rect 121368 3612 121420 3664
rect 121828 3612 121880 3664
rect 122748 3612 122800 3664
rect 122840 3612 122892 3664
rect 252560 3612 252612 3664
rect 2872 3476 2924 3528
rect 4068 3476 4120 3528
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 16028 3476 16080 3528
rect 16488 3476 16540 3528
rect 19524 3476 19576 3528
rect 20628 3476 20680 3528
rect 20720 3476 20772 3528
rect 21916 3476 21968 3528
rect 42156 3476 42208 3528
rect 42708 3476 42760 3528
rect 45376 3476 45428 3528
rect 74632 3476 74684 3528
rect 84016 3476 84068 3528
rect 93952 3476 94004 3528
rect 99472 3476 99524 3528
rect 118792 3476 118844 3528
rect 122656 3476 122708 3528
rect 251180 3544 251232 3596
rect 124220 3476 124272 3528
rect 262220 3476 262272 3528
rect 11244 3408 11296 3460
rect 32404 3408 32456 3460
rect 45468 3408 45520 3460
rect 46848 3408 46900 3460
rect 46940 3408 46992 3460
rect 48136 3408 48188 3460
rect 50528 3408 50580 3460
rect 50988 3408 51040 3460
rect 61108 3408 61160 3460
rect 66260 3408 66312 3460
rect 71872 3408 71924 3460
rect 72976 3408 73028 3460
rect 84108 3408 84160 3460
rect 93860 3408 93912 3460
rect 99380 3408 99432 3460
rect 122932 3408 122984 3460
rect 125416 3408 125468 3460
rect 264980 3408 265032 3460
rect 572 3340 624 3392
rect 59176 3340 59228 3392
rect 63592 3340 63644 3392
rect 64144 3340 64196 3392
rect 73252 3340 73304 3392
rect 175280 3340 175332 3392
rect 1676 3272 1728 3324
rect 62212 3272 62264 3324
rect 6460 3204 6512 3256
rect 6920 3204 6972 3256
rect 21364 3204 21416 3256
rect 35900 3204 35952 3256
rect 36176 3204 36228 3256
rect 45376 3204 45428 3256
rect 46848 3204 46900 3256
rect 68652 3272 68704 3324
rect 73344 3272 73396 3324
rect 171140 3272 171192 3324
rect 64144 3204 64196 3256
rect 162860 3204 162912 3256
rect 5264 3136 5316 3188
rect 6920 3068 6972 3120
rect 21364 3068 21416 3120
rect 29092 3068 29144 3120
rect 57612 3136 57664 3188
rect 153200 3136 153252 3188
rect 39304 3068 39356 3120
rect 56416 3068 56468 3120
rect 151820 3068 151872 3120
rect 35992 3000 36044 3052
rect 51816 3000 51868 3052
rect 54024 3000 54076 3052
rect 147680 3000 147732 3052
rect 42064 2932 42116 2984
rect 49332 2932 49384 2984
rect 139400 2932 139452 2984
rect 38568 2864 38620 2916
rect 45468 2864 45520 2916
rect 45744 2864 45796 2916
rect 133972 2864 134024 2916
rect 43352 2796 43404 2848
rect 129832 2796 129884 2848
rect 70676 1096 70728 1148
rect 73252 1096 73304 1148
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 699718 8156 703520
rect 24320 699718 24348 703520
rect 40512 699990 40540 703520
rect 58808 701004 58860 701010
rect 58808 700946 58860 700952
rect 58716 700936 58768 700942
rect 58716 700878 58768 700884
rect 57704 700664 57756 700670
rect 57704 700606 57756 700612
rect 57612 700188 57664 700194
rect 57612 700130 57664 700136
rect 57520 700120 57572 700126
rect 57520 700062 57572 700068
rect 40500 699984 40552 699990
rect 40500 699926 40552 699932
rect 42064 699984 42116 699990
rect 42064 699926 42116 699932
rect 8116 699712 8168 699718
rect 8116 699654 8168 699660
rect 10324 699712 10376 699718
rect 10324 699654 10376 699660
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 2778 682272 2834 682281
rect 2778 682207 2834 682216
rect 2792 681766 2820 682207
rect 2780 681760 2832 681766
rect 2780 681702 2832 681708
rect 5080 681760 5132 681766
rect 5080 681702 5132 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3882 624880 3938 624889
rect 3882 624815 3938 624824
rect 3896 623830 3924 624815
rect 3884 623824 3936 623830
rect 3884 623766 3936 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 3974 567352 4030 567361
rect 3974 567287 4030 567296
rect 3988 567254 4016 567287
rect 3976 567248 4028 567254
rect 3976 567190 4028 567196
rect 3882 553072 3938 553081
rect 3882 553007 3938 553016
rect 2962 538656 3018 538665
rect 2962 538591 3018 538600
rect 2976 538422 3004 538591
rect 2964 538416 3016 538422
rect 2964 538358 3016 538364
rect 3424 514820 3476 514826
rect 3424 514762 3476 514768
rect 2778 509960 2834 509969
rect 2778 509895 2834 509904
rect 2792 509590 2820 509895
rect 2780 509584 2832 509590
rect 2780 509526 2832 509532
rect 3330 495544 3386 495553
rect 3330 495479 3386 495488
rect 3238 481128 3294 481137
rect 3238 481063 3294 481072
rect 3252 480690 3280 481063
rect 3240 480684 3292 480690
rect 3240 480626 3292 480632
rect 3344 476066 3372 495479
rect 3332 476060 3384 476066
rect 3332 476002 3384 476008
rect 3330 452432 3386 452441
rect 3330 452367 3332 452376
rect 3384 452367 3386 452376
rect 3332 452338 3384 452344
rect 2964 367056 3016 367062
rect 2964 366998 3016 367004
rect 2976 366217 3004 366998
rect 2962 366208 3018 366217
rect 2962 366143 3018 366152
rect 3332 338088 3384 338094
rect 3332 338030 3384 338036
rect 3344 337521 3372 338030
rect 3330 337512 3386 337521
rect 3330 337447 3386 337456
rect 3056 324284 3108 324290
rect 3056 324226 3108 324232
rect 3068 323105 3096 324226
rect 3054 323096 3110 323105
rect 3054 323031 3110 323040
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 2964 295316 3016 295322
rect 2964 295258 3016 295264
rect 2976 294409 3004 295258
rect 2962 294400 3018 294409
rect 2962 294335 3018 294344
rect 3332 280152 3384 280158
rect 3330 280120 3332 280129
rect 3384 280120 3386 280129
rect 3330 280055 3386 280064
rect 3148 266348 3200 266354
rect 3148 266290 3200 266296
rect 3160 265713 3188 266290
rect 3146 265704 3202 265713
rect 3146 265639 3202 265648
rect 3240 237380 3292 237386
rect 3240 237322 3292 237328
rect 3252 237017 3280 237322
rect 3238 237008 3294 237017
rect 3238 236943 3294 236952
rect 3332 223576 3384 223582
rect 3332 223518 3384 223524
rect 3344 222601 3372 223518
rect 3330 222592 3386 222601
rect 3330 222527 3386 222536
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3436 165073 3464 514762
rect 3516 509312 3568 509318
rect 3516 509254 3568 509260
rect 3528 208185 3556 509254
rect 3608 502376 3660 502382
rect 3608 502318 3660 502324
rect 3620 251297 3648 502318
rect 3700 487212 3752 487218
rect 3700 487154 3752 487160
rect 3712 380633 3740 487154
rect 3792 483064 3844 483070
rect 3792 483006 3844 483012
rect 3804 395049 3832 483006
rect 3896 470558 3924 553007
rect 4804 534132 4856 534138
rect 4804 534074 4856 534080
rect 4068 481704 4120 481710
rect 4068 481646 4120 481652
rect 3976 478916 4028 478922
rect 3976 478858 4028 478864
rect 3884 470552 3936 470558
rect 3884 470494 3936 470500
rect 3988 423745 4016 478858
rect 4080 438025 4108 481646
rect 4066 438016 4122 438025
rect 4066 437951 4122 437960
rect 3974 423736 4030 423745
rect 3974 423671 4030 423680
rect 3790 395040 3846 395049
rect 3790 394975 3846 394984
rect 3698 380624 3754 380633
rect 3698 380559 3754 380568
rect 4068 297968 4120 297974
rect 4068 297910 4120 297916
rect 3606 251288 3662 251297
rect 3606 251223 3662 251232
rect 3514 208176 3570 208185
rect 3514 208111 3570 208120
rect 3516 194540 3568 194546
rect 3516 194482 3568 194488
rect 3528 193905 3556 194482
rect 3514 193896 3570 193905
rect 3514 193831 3570 193840
rect 3422 165064 3478 165073
rect 3422 164999 3478 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 2780 122324 2832 122330
rect 2780 122266 2832 122272
rect 2792 122097 2820 122266
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 2780 79824 2832 79830
rect 2780 79766 2832 79772
rect 2792 78985 2820 79766
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 2780 35896 2832 35902
rect 2778 35864 2780 35873
rect 2832 35864 2834 35873
rect 2778 35799 2834 35808
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21457 2912 22034
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 572 3392 624 3398
rect 572 3334 624 3340
rect 584 480 612 3334
rect 1676 3324 1728 3330
rect 1676 3266 1728 3272
rect 1688 480 1716 3266
rect 2884 480 2912 3470
rect 3988 2122 4016 4082
rect 4080 3534 4108 297910
rect 4816 35902 4844 534074
rect 4896 527196 4948 527202
rect 4896 527138 4948 527144
rect 4908 79830 4936 527138
rect 4988 521688 5040 521694
rect 4988 521630 5040 521636
rect 5000 122330 5028 521630
rect 5092 452538 5120 681702
rect 5172 623824 5224 623830
rect 5172 623766 5224 623772
rect 5184 459542 5212 623766
rect 5264 567248 5316 567254
rect 5264 567190 5316 567196
rect 5276 466410 5304 567190
rect 5356 538416 5408 538422
rect 5356 538358 5408 538364
rect 5368 467838 5396 538358
rect 5448 509584 5500 509590
rect 5448 509526 5500 509532
rect 5460 471986 5488 509526
rect 5540 480684 5592 480690
rect 5540 480626 5592 480632
rect 5552 474706 5580 480626
rect 5540 474700 5592 474706
rect 5540 474642 5592 474648
rect 5448 471980 5500 471986
rect 5448 471922 5500 471928
rect 5356 467832 5408 467838
rect 5356 467774 5408 467780
rect 5264 466404 5316 466410
rect 5264 466346 5316 466352
rect 5172 459536 5224 459542
rect 5172 459478 5224 459484
rect 5080 452532 5132 452538
rect 5080 452474 5132 452480
rect 10336 448526 10364 699654
rect 21364 667956 21416 667962
rect 21364 667898 21416 667904
rect 13084 652792 13136 652798
rect 13084 652734 13136 652740
rect 13096 455394 13124 652734
rect 14464 594856 14516 594862
rect 14464 594798 14516 594804
rect 14476 462330 14504 594798
rect 19984 538280 20036 538286
rect 19984 538222 20036 538228
rect 17224 525836 17276 525842
rect 17224 525778 17276 525784
rect 15844 485852 15896 485858
rect 15844 485794 15896 485800
rect 14464 462324 14516 462330
rect 14464 462266 14516 462272
rect 13084 455388 13136 455394
rect 13084 455330 13136 455336
rect 10324 448520 10376 448526
rect 10324 448462 10376 448468
rect 15856 367062 15884 485794
rect 15844 367056 15896 367062
rect 15844 366998 15896 367004
rect 10968 297900 11020 297906
rect 10968 297842 11020 297848
rect 4988 122324 5040 122330
rect 4988 122266 5040 122272
rect 4896 79824 4948 79830
rect 4896 79766 4948 79772
rect 4804 35896 4856 35902
rect 4804 35838 4856 35844
rect 7656 5500 7708 5506
rect 7656 5442 7708 5448
rect 4068 3528 4120 3534
rect 4068 3470 4120 3476
rect 6460 3256 6512 3262
rect 6460 3198 6512 3204
rect 6920 3256 6972 3262
rect 6920 3198 6972 3204
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 3988 2094 4108 2122
rect 4080 480 4108 2094
rect 5276 480 5304 3130
rect 6472 480 6500 3198
rect 6932 3126 6960 3198
rect 6920 3120 6972 3126
rect 6920 3062 6972 3068
rect 7668 480 7696 5442
rect 8852 4072 8904 4078
rect 8852 4014 8904 4020
rect 8864 480 8892 4014
rect 10980 3534 11008 297842
rect 16488 297832 16540 297838
rect 16488 297774 16540 297780
rect 15108 297696 15160 297702
rect 15108 297638 15160 297644
rect 12440 5432 12492 5438
rect 12440 5374 12492 5380
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10060 480 10088 3470
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11256 480 11284 3402
rect 12452 480 12480 5374
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13648 480 13676 3946
rect 15120 3482 15148 297638
rect 16500 3534 16528 297774
rect 17236 109002 17264 525778
rect 17316 491360 17368 491366
rect 17316 491302 17368 491308
rect 17328 309126 17356 491302
rect 17316 309120 17368 309126
rect 17316 309062 17368 309068
rect 17224 108996 17276 109002
rect 17224 108938 17276 108944
rect 19996 22098 20024 538222
rect 20076 498228 20128 498234
rect 20076 498170 20128 498176
rect 20088 266354 20116 498170
rect 21376 456754 21404 667898
rect 21364 456748 21416 456754
rect 21364 456690 21416 456696
rect 24780 451246 24808 699654
rect 31024 610020 31076 610026
rect 31024 609962 31076 609968
rect 28264 505164 28316 505170
rect 28264 505106 28316 505112
rect 24768 451240 24820 451246
rect 24768 451182 24820 451188
rect 20628 297628 20680 297634
rect 20628 297570 20680 297576
rect 20076 266348 20128 266354
rect 20076 266290 20128 266296
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 17224 5364 17276 5370
rect 17224 5306 17276 5312
rect 14844 3454 15148 3482
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 14844 480 14872 3454
rect 16040 480 16068 3470
rect 17236 480 17264 5306
rect 18328 3936 18380 3942
rect 18328 3878 18380 3884
rect 18340 480 18368 3878
rect 20640 3534 20668 297570
rect 21916 297560 21968 297566
rect 21916 297502 21968 297508
rect 21928 3534 21956 297502
rect 24768 297492 24820 297498
rect 24768 297434 24820 297440
rect 22008 5228 22060 5234
rect 22008 5170 22060 5176
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 21916 3528 21968 3534
rect 21916 3470 21968 3476
rect 19536 480 19564 3470
rect 20732 480 20760 3470
rect 21364 3256 21416 3262
rect 21364 3198 21416 3204
rect 21376 3126 21404 3198
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 22020 2666 22048 5170
rect 24780 3874 24808 297434
rect 26148 297424 26200 297430
rect 26148 297366 26200 297372
rect 26160 3874 26188 297366
rect 28276 223582 28304 505106
rect 31036 463690 31064 609962
rect 35164 517540 35216 517546
rect 35164 517482 35216 517488
rect 33784 510672 33836 510678
rect 33784 510614 33836 510620
rect 32404 494080 32456 494086
rect 32404 494022 32456 494028
rect 31024 463684 31076 463690
rect 31024 463626 31076 463632
rect 32416 324290 32444 494022
rect 32404 324284 32456 324290
rect 32404 324226 32456 324232
rect 32404 298036 32456 298042
rect 32404 297978 32456 297984
rect 28264 223576 28316 223582
rect 28264 223518 28316 223524
rect 26700 5160 26752 5166
rect 26700 5102 26752 5108
rect 24308 3868 24360 3874
rect 24308 3810 24360 3816
rect 24768 3868 24820 3874
rect 24768 3810 24820 3816
rect 25504 3868 25556 3874
rect 25504 3810 25556 3816
rect 26148 3868 26200 3874
rect 26148 3810 26200 3816
rect 23112 3800 23164 3806
rect 23112 3742 23164 3748
rect 21928 2638 22048 2666
rect 21928 480 21956 2638
rect 23124 480 23152 3742
rect 24320 480 24348 3810
rect 25516 480 25544 3810
rect 26712 480 26740 5102
rect 30288 5092 30340 5098
rect 30288 5034 30340 5040
rect 27896 3800 27948 3806
rect 27896 3742 27948 3748
rect 27908 480 27936 3742
rect 29092 3120 29144 3126
rect 29092 3062 29144 3068
rect 29104 480 29132 3062
rect 30300 480 30328 5034
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31496 480 31524 3674
rect 32416 3466 32444 297978
rect 33796 180810 33824 510614
rect 33784 180804 33836 180810
rect 33784 180746 33836 180752
rect 35176 136610 35204 517482
rect 39396 506524 39448 506530
rect 39396 506466 39448 506472
rect 37924 501016 37976 501022
rect 37924 500958 37976 500964
rect 37936 280158 37964 500958
rect 39304 298104 39356 298110
rect 39304 298046 39356 298052
rect 37924 280152 37976 280158
rect 37924 280094 37976 280100
rect 35164 136604 35216 136610
rect 35164 136546 35216 136552
rect 33876 5024 33928 5030
rect 33876 4966 33928 4972
rect 32680 3596 32732 3602
rect 32680 3538 32732 3544
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 32692 480 32720 3538
rect 33888 480 33916 4966
rect 37372 4956 37424 4962
rect 37372 4898 37424 4904
rect 34980 3664 35032 3670
rect 34980 3606 35032 3612
rect 34992 480 35020 3606
rect 35900 3256 35952 3262
rect 36176 3256 36228 3262
rect 35952 3204 36032 3210
rect 35900 3198 36032 3204
rect 36176 3198 36228 3204
rect 35912 3182 36032 3198
rect 36004 3058 36032 3182
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 36188 480 36216 3198
rect 37384 480 37412 4898
rect 39316 3126 39344 298046
rect 39408 237386 39436 506466
rect 42076 447098 42104 699926
rect 57428 650888 57480 650894
rect 57428 650830 57480 650836
rect 56598 646096 56654 646105
rect 56598 646031 56654 646040
rect 56612 543017 56640 646031
rect 57242 645008 57298 645017
rect 57242 644943 57298 644952
rect 57150 643240 57206 643249
rect 57150 643175 57206 643184
rect 57058 642016 57114 642025
rect 57058 641951 57114 641960
rect 56966 640384 57022 640393
rect 56966 640319 57022 640328
rect 56874 639296 56930 639305
rect 56874 639231 56930 639240
rect 56782 637664 56838 637673
rect 56782 637599 56838 637608
rect 56690 579728 56746 579737
rect 56690 579663 56746 579672
rect 56704 543046 56732 579663
rect 56796 543726 56824 637599
rect 56784 543720 56836 543726
rect 56784 543662 56836 543668
rect 56888 543658 56916 639231
rect 56876 543652 56928 543658
rect 56876 543594 56928 543600
rect 56980 543522 57008 640319
rect 56968 543516 57020 543522
rect 56968 543458 57020 543464
rect 57072 543454 57100 641951
rect 57060 543448 57112 543454
rect 57060 543390 57112 543396
rect 57164 543386 57192 643175
rect 57152 543380 57204 543386
rect 57152 543322 57204 543328
rect 57256 543318 57284 644943
rect 57336 545148 57388 545154
rect 57336 545090 57388 545096
rect 57244 543312 57296 543318
rect 57244 543254 57296 543260
rect 56692 543040 56744 543046
rect 56598 543008 56654 543017
rect 56692 542982 56744 542988
rect 56598 542943 56654 542952
rect 56784 540320 56836 540326
rect 56784 540262 56836 540268
rect 56692 540252 56744 540258
rect 56692 540194 56744 540200
rect 48964 536852 49016 536858
rect 48964 536794 49016 536800
rect 46204 529984 46256 529990
rect 46204 529926 46256 529932
rect 43444 523048 43496 523054
rect 43444 522990 43496 522996
rect 42064 447092 42116 447098
rect 42064 447034 42116 447040
rect 42708 297764 42760 297770
rect 42708 297706 42760 297712
rect 39948 296812 40000 296818
rect 39948 296754 40000 296760
rect 39396 237380 39448 237386
rect 39396 237322 39448 237328
rect 39960 3346 39988 296754
rect 42064 296744 42116 296750
rect 42064 296686 42116 296692
rect 40960 4888 41012 4894
rect 40960 4830 41012 4836
rect 39776 3318 39988 3346
rect 39304 3120 39356 3126
rect 39304 3062 39356 3068
rect 38568 2916 38620 2922
rect 38568 2858 38620 2864
rect 38580 480 38608 2858
rect 39776 480 39804 3318
rect 40972 480 41000 4830
rect 42076 2990 42104 296686
rect 42720 3534 42748 297706
rect 43456 93838 43484 522990
rect 43444 93832 43496 93838
rect 43444 93774 43496 93780
rect 46216 51066 46244 529926
rect 48136 296880 48188 296886
rect 48136 296822 48188 296828
rect 46204 51060 46256 51066
rect 46204 51002 46256 51008
rect 44548 4820 44600 4826
rect 44548 4762 44600 4768
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 42064 2984 42116 2990
rect 42064 2926 42116 2932
rect 42168 480 42196 3470
rect 43352 2848 43404 2854
rect 43352 2790 43404 2796
rect 43364 480 43392 2790
rect 44560 480 44588 4762
rect 45376 3528 45428 3534
rect 45376 3470 45428 3476
rect 45388 3262 45416 3470
rect 48148 3466 48176 296822
rect 48976 8294 49004 536794
rect 53104 531412 53156 531418
rect 53104 531354 53156 531360
rect 51724 518968 51776 518974
rect 51724 518910 51776 518916
rect 50344 513392 50396 513398
rect 50344 513334 50396 513340
rect 50356 194546 50384 513334
rect 50988 296948 51040 296954
rect 50988 296890 51040 296896
rect 50344 194540 50396 194546
rect 50344 194482 50396 194488
rect 48964 8288 49016 8294
rect 48964 8230 49016 8236
rect 48228 4208 48280 4214
rect 48228 4150 48280 4156
rect 45468 3460 45520 3466
rect 45468 3402 45520 3408
rect 46848 3460 46900 3466
rect 46848 3402 46900 3408
rect 46940 3460 46992 3466
rect 46940 3402 46992 3408
rect 48136 3460 48188 3466
rect 48136 3402 48188 3408
rect 45376 3256 45428 3262
rect 45376 3198 45428 3204
rect 45480 2922 45508 3402
rect 46860 3262 46888 3402
rect 46848 3256 46900 3262
rect 46848 3198 46900 3204
rect 45468 2916 45520 2922
rect 45468 2858 45520 2864
rect 45744 2916 45796 2922
rect 45744 2858 45796 2864
rect 45756 480 45784 2858
rect 46952 480 46980 3402
rect 48240 2122 48268 4150
rect 51000 3466 51028 296890
rect 51736 151774 51764 518910
rect 51816 297356 51868 297362
rect 51816 297298 51868 297304
rect 51724 151768 51776 151774
rect 51724 151710 51776 151716
rect 51632 4276 51684 4282
rect 51632 4218 51684 4224
rect 50528 3460 50580 3466
rect 50528 3402 50580 3408
rect 50988 3460 51040 3466
rect 50988 3402 51040 3408
rect 49332 2984 49384 2990
rect 49332 2926 49384 2932
rect 48148 2094 48268 2122
rect 48148 480 48176 2094
rect 49344 480 49372 2926
rect 50540 480 50568 3402
rect 51644 480 51672 4218
rect 51828 3058 51856 297298
rect 53116 64870 53144 531354
rect 56598 488336 56654 488345
rect 56598 488271 56654 488280
rect 56612 487218 56640 488271
rect 56600 487212 56652 487218
rect 56600 487154 56652 487160
rect 56598 486296 56654 486305
rect 56598 486231 56654 486240
rect 56612 485858 56640 486231
rect 56600 485852 56652 485858
rect 56600 485794 56652 485800
rect 56598 484120 56654 484129
rect 56598 484055 56654 484064
rect 56612 483070 56640 484055
rect 56600 483064 56652 483070
rect 56600 483006 56652 483012
rect 56598 482080 56654 482089
rect 56598 482015 56654 482024
rect 56612 481710 56640 482015
rect 56600 481704 56652 481710
rect 56600 481646 56652 481652
rect 56598 480040 56654 480049
rect 56598 479975 56654 479984
rect 56612 478922 56640 479975
rect 56600 478916 56652 478922
rect 56600 478858 56652 478864
rect 56598 477864 56654 477873
rect 56598 477799 56654 477808
rect 56612 476218 56640 477799
rect 56520 476190 56640 476218
rect 56520 475674 56548 476190
rect 56600 476060 56652 476066
rect 56600 476002 56652 476008
rect 56612 475833 56640 476002
rect 56598 475824 56654 475833
rect 56598 475759 56654 475768
rect 56520 475646 56640 475674
rect 56612 474858 56640 475646
rect 56520 474830 56640 474858
rect 56520 473498 56548 474830
rect 56600 474700 56652 474706
rect 56600 474642 56652 474648
rect 56612 473657 56640 474642
rect 56598 473648 56654 473657
rect 56598 473583 56654 473592
rect 56520 473470 56640 473498
rect 56612 472138 56640 473470
rect 56520 472110 56640 472138
rect 56520 471458 56548 472110
rect 56600 471980 56652 471986
rect 56600 471922 56652 471928
rect 56612 471617 56640 471922
rect 56598 471608 56654 471617
rect 56598 471543 56654 471552
rect 56520 471430 56640 471458
rect 56508 470552 56560 470558
rect 56508 470494 56560 470500
rect 56520 469985 56548 470494
rect 56506 469976 56562 469985
rect 56506 469911 56562 469920
rect 56508 467832 56560 467838
rect 56506 467800 56508 467809
rect 56560 467800 56562 467809
rect 56506 467735 56562 467744
rect 56508 466404 56560 466410
rect 56508 466346 56560 466352
rect 56520 465769 56548 466346
rect 56506 465760 56562 465769
rect 56506 465695 56562 465704
rect 56508 463684 56560 463690
rect 56508 463626 56560 463632
rect 56520 463593 56548 463626
rect 56506 463584 56562 463593
rect 56506 463519 56562 463528
rect 56508 462324 56560 462330
rect 56508 462266 56560 462272
rect 56520 461553 56548 462266
rect 56506 461544 56562 461553
rect 56506 461479 56562 461488
rect 56612 459626 56640 471430
rect 56520 459598 56640 459626
rect 56520 458810 56548 459598
rect 56600 459536 56652 459542
rect 56600 459478 56652 459484
rect 56612 458969 56640 459478
rect 56598 458960 56654 458969
rect 56598 458895 56654 458904
rect 56520 458782 56640 458810
rect 56612 456906 56640 458782
rect 56520 456878 56640 456906
rect 56520 456634 56548 456878
rect 56598 456784 56654 456793
rect 56598 456719 56600 456728
rect 56652 456719 56654 456728
rect 56600 456690 56652 456696
rect 56520 456606 56640 456634
rect 56612 455546 56640 456606
rect 56520 455518 56640 455546
rect 56520 454594 56548 455518
rect 56600 455388 56652 455394
rect 56600 455330 56652 455336
rect 56612 454753 56640 455330
rect 56598 454744 56654 454753
rect 56598 454679 56654 454688
rect 56520 454566 56640 454594
rect 56612 452690 56640 454566
rect 56520 452662 56640 452690
rect 56520 452402 56548 452662
rect 56598 452568 56654 452577
rect 56598 452503 56600 452512
rect 56652 452503 56654 452512
rect 56600 452474 56652 452480
rect 56508 452396 56560 452402
rect 56508 452338 56560 452344
rect 56600 451240 56652 451246
rect 56600 451182 56652 451188
rect 56612 450537 56640 451182
rect 56598 450528 56654 450537
rect 56598 450463 56654 450472
rect 56600 448656 56652 448662
rect 56600 448598 56652 448604
rect 56612 444145 56640 448598
rect 56598 444136 56654 444145
rect 56598 444071 56654 444080
rect 56704 433673 56732 540194
rect 56690 433664 56746 433673
rect 56690 433599 56746 433608
rect 56796 427281 56824 540262
rect 56876 539232 56928 539238
rect 56876 539174 56928 539180
rect 56782 427272 56838 427281
rect 56782 427207 56838 427216
rect 56888 421025 56916 539174
rect 57242 538928 57298 538937
rect 57060 538892 57112 538898
rect 57242 538863 57298 538872
rect 57060 538834 57112 538840
rect 56966 496768 57022 496777
rect 56966 496703 57022 496712
rect 56980 491230 57008 496703
rect 56968 491224 57020 491230
rect 56968 491166 57020 491172
rect 56966 490512 57022 490521
rect 56966 490447 57022 490456
rect 56874 421016 56930 421025
rect 56874 420951 56930 420960
rect 56598 353696 56654 353705
rect 56598 353631 56654 353640
rect 56612 320142 56640 353631
rect 56690 343088 56746 343097
rect 56690 343023 56746 343032
rect 56600 320136 56652 320142
rect 56600 320078 56652 320084
rect 56600 315988 56652 315994
rect 56600 315930 56652 315936
rect 56612 309482 56640 315930
rect 56520 309454 56640 309482
rect 56520 306406 56548 309454
rect 56598 309360 56654 309369
rect 56598 309295 56654 309304
rect 56508 306400 56560 306406
rect 56508 306342 56560 306348
rect 56612 88330 56640 309295
rect 56704 300762 56732 343023
rect 56782 338872 56838 338881
rect 56782 338807 56838 338816
rect 56692 300756 56744 300762
rect 56692 300698 56744 300704
rect 56796 299470 56824 338807
rect 56980 338094 57008 490447
rect 57072 381041 57100 538834
rect 57256 538286 57284 538863
rect 57244 538280 57296 538286
rect 57244 538222 57296 538228
rect 57152 537940 57204 537946
rect 57152 537882 57204 537888
rect 57058 381032 57114 381041
rect 57058 380967 57114 380976
rect 57164 366217 57192 537882
rect 57242 536888 57298 536897
rect 57242 536823 57244 536832
rect 57296 536823 57298 536832
rect 57244 536794 57296 536800
rect 57242 534712 57298 534721
rect 57242 534647 57298 534656
rect 57256 534138 57284 534647
rect 57244 534132 57296 534138
rect 57244 534074 57296 534080
rect 57242 532672 57298 532681
rect 57242 532607 57298 532616
rect 57256 531418 57284 532607
rect 57244 531412 57296 531418
rect 57244 531354 57296 531360
rect 57242 530496 57298 530505
rect 57242 530431 57298 530440
rect 57256 529990 57284 530431
rect 57244 529984 57296 529990
rect 57244 529926 57296 529932
rect 57242 528456 57298 528465
rect 57242 528391 57298 528400
rect 57256 527202 57284 528391
rect 57244 527196 57296 527202
rect 57244 527138 57296 527144
rect 57242 526280 57298 526289
rect 57242 526215 57298 526224
rect 57256 525842 57284 526215
rect 57244 525836 57296 525842
rect 57244 525778 57296 525784
rect 57242 524240 57298 524249
rect 57242 524175 57298 524184
rect 57256 523054 57284 524175
rect 57244 523048 57296 523054
rect 57244 522990 57296 522996
rect 57242 522064 57298 522073
rect 57242 521999 57298 522008
rect 57256 521694 57284 521999
rect 57244 521688 57296 521694
rect 57244 521630 57296 521636
rect 57242 520024 57298 520033
rect 57242 519959 57298 519968
rect 57256 518974 57284 519959
rect 57244 518968 57296 518974
rect 57244 518910 57296 518916
rect 57242 517848 57298 517857
rect 57242 517783 57298 517792
rect 57256 517546 57284 517783
rect 57244 517540 57296 517546
rect 57244 517482 57296 517488
rect 57242 515808 57298 515817
rect 57242 515743 57298 515752
rect 57256 514826 57284 515743
rect 57244 514820 57296 514826
rect 57244 514762 57296 514768
rect 57242 513632 57298 513641
rect 57242 513567 57298 513576
rect 57256 513398 57284 513567
rect 57244 513392 57296 513398
rect 57244 513334 57296 513340
rect 57242 511592 57298 511601
rect 57242 511527 57298 511536
rect 57256 510678 57284 511527
rect 57244 510672 57296 510678
rect 57244 510614 57296 510620
rect 57242 509416 57298 509425
rect 57242 509351 57298 509360
rect 57256 509318 57284 509351
rect 57244 509312 57296 509318
rect 57244 509254 57296 509260
rect 57242 507376 57298 507385
rect 57242 507311 57298 507320
rect 57256 506530 57284 507311
rect 57244 506524 57296 506530
rect 57244 506466 57296 506472
rect 57242 505200 57298 505209
rect 57242 505135 57244 505144
rect 57296 505135 57298 505144
rect 57244 505106 57296 505112
rect 57242 503160 57298 503169
rect 57242 503095 57298 503104
rect 57256 502382 57284 503095
rect 57244 502376 57296 502382
rect 57244 502318 57296 502324
rect 57244 501016 57296 501022
rect 57242 500984 57244 500993
rect 57296 500984 57298 500993
rect 57242 500919 57298 500928
rect 57242 498944 57298 498953
rect 57242 498879 57298 498888
rect 57256 498234 57284 498879
rect 57244 498228 57296 498234
rect 57244 498170 57296 498176
rect 57242 494728 57298 494737
rect 57242 494663 57298 494672
rect 57256 494086 57284 494663
rect 57244 494080 57296 494086
rect 57244 494022 57296 494028
rect 57242 492552 57298 492561
rect 57242 492487 57298 492496
rect 57256 491366 57284 492487
rect 57244 491360 57296 491366
rect 57244 491302 57296 491308
rect 57244 491224 57296 491230
rect 57244 491166 57296 491172
rect 57150 366208 57206 366217
rect 57150 366143 57206 366152
rect 57058 361992 57114 362001
rect 57058 361927 57114 361936
rect 57072 339454 57100 361927
rect 57150 355736 57206 355745
rect 57150 355671 57206 355680
rect 57060 339448 57112 339454
rect 57060 339390 57112 339396
rect 56968 338088 57020 338094
rect 56968 338030 57020 338036
rect 56966 336832 57022 336841
rect 56966 336767 57022 336776
rect 56874 334656 56930 334665
rect 56874 334591 56930 334600
rect 56784 299464 56836 299470
rect 56784 299406 56836 299412
rect 56782 296712 56838 296721
rect 56692 296676 56744 296682
rect 56782 296647 56838 296656
rect 56692 296618 56744 296624
rect 56704 287094 56732 296618
rect 56796 287162 56824 296647
rect 56784 287156 56836 287162
rect 56784 287098 56836 287104
rect 56692 287088 56744 287094
rect 56692 287030 56744 287036
rect 56782 277400 56838 277409
rect 56782 277335 56838 277344
rect 56796 268462 56824 277335
rect 56888 276010 56916 334591
rect 56876 276004 56928 276010
rect 56876 275946 56928 275952
rect 56784 268456 56836 268462
rect 56784 268398 56836 268404
rect 56980 264926 57008 336767
rect 57058 332616 57114 332625
rect 57058 332551 57114 332560
rect 56968 264920 57020 264926
rect 56968 264862 57020 264868
rect 57072 252550 57100 332551
rect 57164 331634 57192 355671
rect 57152 331628 57204 331634
rect 57152 331570 57204 331576
rect 57150 328400 57206 328409
rect 57150 328335 57206 328344
rect 57060 252544 57112 252550
rect 57060 252486 57112 252492
rect 57164 229090 57192 328335
rect 57256 295322 57284 491166
rect 57348 374649 57376 545090
rect 57440 439929 57468 650830
rect 57532 448662 57560 700062
rect 57520 448656 57572 448662
rect 57520 448598 57572 448604
rect 57520 448520 57572 448526
rect 57520 448462 57572 448468
rect 57532 448361 57560 448462
rect 57518 448352 57574 448361
rect 57518 448287 57574 448296
rect 57520 447092 57572 447098
rect 57520 447034 57572 447040
rect 57532 446321 57560 447034
rect 57518 446312 57574 446321
rect 57518 446247 57574 446256
rect 57426 439920 57482 439929
rect 57426 439855 57482 439864
rect 57624 437889 57652 700130
rect 57610 437880 57666 437889
rect 57610 437815 57666 437824
rect 57612 434036 57664 434042
rect 57612 433978 57664 433984
rect 57334 374640 57390 374649
rect 57334 374575 57390 374584
rect 57624 368393 57652 433978
rect 57716 418985 57744 700606
rect 57796 700528 57848 700534
rect 57796 700470 57848 700476
rect 57702 418976 57758 418985
rect 57702 418911 57758 418920
rect 57704 413976 57756 413982
rect 57704 413918 57756 413924
rect 57610 368384 57666 368393
rect 57610 368319 57666 368328
rect 57716 364177 57744 413918
rect 57808 412593 57836 700470
rect 57888 700460 57940 700466
rect 57888 700402 57940 700408
rect 57794 412584 57850 412593
rect 57794 412519 57850 412528
rect 57900 406337 57928 700402
rect 58532 700256 58584 700262
rect 58532 700198 58584 700204
rect 58440 700052 58492 700058
rect 58440 699994 58492 700000
rect 58348 650752 58400 650758
rect 58348 650694 58400 650700
rect 58256 556232 58308 556238
rect 58256 556174 58308 556180
rect 57980 539028 58032 539034
rect 57980 538970 58032 538976
rect 57886 406328 57942 406337
rect 57886 406263 57942 406272
rect 57992 383081 58020 538970
rect 58072 538960 58124 538966
rect 58072 538902 58124 538908
rect 57978 383072 58034 383081
rect 57978 383007 58034 383016
rect 58084 376825 58112 538902
rect 58164 538280 58216 538286
rect 58164 538222 58216 538228
rect 58070 376816 58126 376825
rect 58070 376751 58126 376760
rect 58176 370433 58204 538222
rect 58268 372609 58296 556174
rect 58360 404161 58388 650694
rect 58452 442105 58480 699994
rect 58438 442096 58494 442105
rect 58438 442031 58494 442040
rect 58544 435713 58572 700198
rect 58624 650344 58676 650350
rect 58624 650286 58676 650292
rect 58530 435704 58586 435713
rect 58530 435639 58586 435648
rect 58346 404152 58402 404161
rect 58346 404087 58402 404096
rect 58636 385257 58664 650286
rect 58728 431497 58756 700878
rect 58714 431488 58770 431497
rect 58714 431423 58770 431432
rect 58820 429457 58848 700946
rect 58992 700868 59044 700874
rect 58992 700810 59044 700816
rect 58900 700800 58952 700806
rect 58900 700742 58952 700748
rect 58806 429448 58862 429457
rect 58806 429383 58862 429392
rect 58716 429208 58768 429214
rect 58716 429150 58768 429156
rect 58728 413982 58756 429150
rect 58912 425241 58940 700742
rect 58898 425232 58954 425241
rect 58898 425167 58954 425176
rect 59004 423065 59032 700810
rect 59084 700732 59136 700738
rect 59084 700674 59136 700680
rect 58990 423056 59046 423065
rect 58990 422991 59046 423000
rect 59096 416809 59124 700674
rect 59176 700596 59228 700602
rect 59176 700538 59228 700544
rect 59082 416800 59138 416809
rect 59082 416735 59138 416744
rect 58716 413976 58768 413982
rect 58716 413918 58768 413924
rect 59188 410553 59216 700538
rect 59268 700392 59320 700398
rect 59268 700334 59320 700340
rect 59174 410544 59230 410553
rect 59174 410479 59230 410488
rect 59280 397905 59308 700334
rect 59360 700324 59412 700330
rect 59360 700266 59412 700272
rect 59372 399945 59400 700266
rect 72988 700058 73016 703520
rect 89180 700126 89208 703520
rect 105464 703474 105492 703520
rect 105464 703446 105584 703474
rect 89168 700120 89220 700126
rect 89168 700062 89220 700068
rect 72976 700052 73028 700058
rect 72976 699994 73028 700000
rect 105556 698290 105584 703446
rect 136640 700256 136692 700262
rect 136640 700198 136692 700204
rect 137284 700256 137336 700262
rect 137284 700198 137336 700204
rect 136652 700126 136680 700198
rect 136640 700120 136692 700126
rect 136640 700062 136692 700068
rect 104992 698284 105044 698290
rect 104992 698226 105044 698232
rect 105544 698284 105596 698290
rect 105544 698226 105596 698232
rect 77206 697232 77262 697241
rect 77206 697167 77262 697176
rect 96526 697232 96582 697241
rect 96526 697167 96582 697176
rect 77220 697134 77248 697167
rect 96540 697134 96568 697167
rect 70308 697128 70360 697134
rect 70306 697096 70308 697105
rect 77208 697128 77260 697134
rect 70360 697096 70362 697105
rect 89628 697128 89680 697134
rect 77208 697070 77260 697076
rect 89626 697096 89628 697105
rect 96528 697128 96580 697134
rect 89680 697096 89682 697105
rect 70306 697031 70362 697040
rect 96528 697070 96580 697076
rect 89626 697031 89682 697040
rect 105004 688650 105032 698226
rect 115846 697232 115902 697241
rect 115846 697167 115902 697176
rect 135166 697232 135222 697241
rect 135166 697167 135222 697176
rect 115860 697134 115888 697167
rect 135180 697134 135208 697167
rect 108948 697128 109000 697134
rect 108946 697096 108948 697105
rect 115848 697128 115900 697134
rect 109000 697096 109002 697105
rect 128268 697128 128320 697134
rect 115848 697070 115900 697076
rect 128266 697096 128268 697105
rect 135168 697128 135220 697134
rect 128320 697096 128322 697105
rect 108946 697031 109002 697040
rect 135168 697070 135220 697076
rect 128266 697031 128322 697040
rect 104912 688622 105032 688650
rect 104912 683074 104940 688622
rect 104912 683046 105124 683074
rect 105096 673538 105124 683046
rect 104900 673532 104952 673538
rect 104900 673474 104952 673480
rect 105084 673532 105136 673538
rect 105084 673474 105136 673480
rect 104912 663762 104940 673474
rect 104912 663734 105124 663762
rect 105096 654158 105124 663734
rect 104900 654152 104952 654158
rect 104900 654094 104952 654100
rect 105084 654152 105136 654158
rect 105084 654094 105136 654100
rect 104912 650894 104940 654094
rect 129278 652896 129334 652905
rect 129278 652831 129334 652840
rect 133602 652896 133658 652905
rect 133602 652831 133658 652840
rect 129292 652798 129320 652831
rect 133616 652798 133644 652831
rect 129280 652792 129332 652798
rect 129280 652734 129332 652740
rect 133604 652792 133656 652798
rect 133604 652734 133656 652740
rect 104900 650888 104952 650894
rect 104900 650830 104952 650836
rect 59544 650820 59596 650826
rect 59544 650762 59596 650768
rect 59452 650684 59504 650690
rect 59452 650626 59504 650632
rect 59464 402121 59492 650626
rect 59556 414769 59584 650762
rect 59634 578583 59690 578592
rect 59634 578518 59690 578527
rect 59648 560930 59676 578518
rect 59636 560924 59688 560930
rect 59636 560866 59688 560872
rect 67546 558920 67602 558929
rect 67546 558855 67602 558864
rect 70122 558920 70178 558929
rect 70122 558855 70178 558864
rect 72422 558920 72478 558929
rect 72422 558855 72478 558864
rect 73710 558920 73766 558929
rect 73710 558855 73766 558864
rect 75734 558920 75790 558929
rect 75734 558855 75790 558864
rect 76010 558920 76066 558929
rect 76010 558855 76066 558864
rect 77390 558920 77446 558929
rect 77390 558855 77446 558864
rect 78494 558920 78550 558929
rect 79506 558920 79562 558929
rect 78494 558855 78550 558864
rect 79324 558884 79376 558890
rect 64326 558784 64382 558793
rect 64326 558719 64382 558728
rect 64340 558210 64368 558719
rect 64328 558204 64380 558210
rect 64328 558146 64380 558152
rect 66168 557796 66220 557802
rect 66168 557738 66220 557744
rect 63408 557660 63460 557666
rect 63408 557602 63460 557608
rect 62028 557592 62080 557598
rect 62028 557534 62080 557540
rect 62040 543590 62068 557534
rect 61016 543584 61068 543590
rect 61016 543526 61068 543532
rect 62028 543584 62080 543590
rect 62028 543526 62080 543532
rect 61028 539988 61056 543526
rect 63420 540002 63448 557602
rect 66180 543318 66208 557738
rect 67456 557728 67508 557734
rect 67456 557670 67508 557676
rect 65156 543312 65208 543318
rect 65156 543254 65208 543260
rect 66168 543312 66220 543318
rect 66168 543254 66220 543260
rect 63066 539974 63448 540002
rect 65168 539988 65196 543254
rect 67468 540002 67496 557670
rect 67560 542978 67588 558855
rect 68926 558104 68982 558113
rect 68926 558039 68982 558048
rect 67548 542972 67600 542978
rect 67548 542914 67600 542920
rect 68940 542910 68968 558039
rect 70136 543250 70164 558855
rect 70214 558784 70270 558793
rect 70214 558719 70270 558728
rect 70124 543244 70176 543250
rect 70124 543186 70176 543192
rect 70228 543182 70256 558719
rect 72436 558550 72464 558855
rect 72424 558544 72476 558550
rect 72424 558486 72476 558492
rect 73724 558414 73752 558855
rect 75748 558618 75776 558855
rect 75736 558612 75788 558618
rect 75736 558554 75788 558560
rect 76024 558482 76052 558855
rect 77404 558686 77432 558855
rect 77392 558680 77444 558686
rect 77392 558622 77444 558628
rect 76012 558476 76064 558482
rect 76012 558418 76064 558424
rect 73712 558408 73764 558414
rect 73712 558350 73764 558356
rect 77298 558376 77354 558385
rect 75828 558340 75880 558346
rect 77298 558311 77354 558320
rect 75828 558282 75880 558288
rect 73158 558240 73214 558249
rect 73158 558175 73214 558184
rect 71688 557932 71740 557938
rect 71688 557874 71740 557880
rect 70308 557864 70360 557870
rect 70308 557806 70360 557812
rect 70216 543176 70268 543182
rect 70216 543118 70268 543124
rect 68928 542904 68980 542910
rect 68928 542846 68980 542852
rect 70320 542706 70348 557806
rect 71594 557560 71650 557569
rect 71594 557495 71650 557504
rect 71608 543114 71636 557495
rect 71596 543108 71648 543114
rect 71596 543050 71648 543056
rect 69296 542700 69348 542706
rect 69296 542642 69348 542648
rect 70308 542700 70360 542706
rect 70308 542642 70360 542648
rect 67206 539974 67496 540002
rect 69308 539988 69336 542642
rect 71700 540002 71728 557874
rect 71778 557696 71834 557705
rect 73172 557666 73200 558175
rect 74538 557832 74594 557841
rect 74538 557767 74540 557776
rect 74592 557767 74594 557776
rect 74540 557738 74592 557744
rect 71778 557631 71834 557640
rect 73160 557660 73212 557666
rect 71792 557598 71820 557631
rect 73160 557602 73212 557608
rect 71780 557592 71832 557598
rect 71780 557534 71832 557540
rect 74448 557592 74500 557598
rect 74448 557534 74500 557540
rect 74460 543318 74488 557534
rect 73436 543312 73488 543318
rect 73436 543254 73488 543260
rect 74448 543312 74500 543318
rect 74448 543254 74500 543260
rect 71346 539974 71728 540002
rect 73448 539988 73476 543254
rect 75840 540002 75868 558282
rect 77312 557870 77340 558311
rect 78508 558278 78536 558855
rect 79506 558855 79562 558864
rect 80702 558920 80758 558929
rect 80702 558855 80758 558864
rect 81438 558920 81494 558929
rect 82910 558920 82966 558929
rect 81438 558855 81440 558864
rect 79324 558826 79376 558832
rect 78496 558272 78548 558278
rect 78496 558214 78548 558220
rect 78678 557968 78734 557977
rect 78678 557903 78680 557912
rect 78732 557903 78734 557912
rect 78680 557874 78732 557880
rect 77300 557864 77352 557870
rect 75918 557832 75974 557841
rect 77300 557806 77352 557812
rect 75918 557767 75974 557776
rect 75932 557734 75960 557767
rect 75920 557728 75972 557734
rect 75920 557670 75972 557676
rect 78678 557696 78734 557705
rect 78678 557631 78734 557640
rect 78692 557598 78720 557631
rect 78680 557592 78732 557598
rect 78680 557534 78732 557540
rect 79336 543318 79364 558826
rect 79520 558754 79548 558855
rect 80716 558822 80744 558855
rect 81492 558855 81494 558864
rect 81532 558884 81584 558890
rect 81440 558826 81492 558832
rect 82910 558855 82966 558864
rect 84198 558920 84254 558929
rect 84198 558855 84254 558864
rect 85394 558920 85450 558929
rect 85394 558855 85450 558864
rect 85670 558920 85726 558929
rect 85670 558855 85726 558864
rect 86222 558920 86278 558929
rect 87602 558920 87658 558929
rect 86222 558855 86278 558864
rect 86868 558884 86920 558890
rect 81532 558826 81584 558832
rect 80704 558816 80756 558822
rect 80058 558784 80114 558793
rect 79508 558748 79560 558754
rect 80704 558758 80756 558764
rect 80058 558719 80114 558728
rect 79508 558690 79560 558696
rect 80072 558346 80100 558719
rect 81544 558686 81572 558826
rect 81622 558784 81678 558793
rect 81622 558719 81678 558728
rect 81636 558686 81664 558719
rect 81532 558680 81584 558686
rect 81532 558622 81584 558628
rect 81624 558680 81676 558686
rect 81624 558622 81676 558628
rect 81636 558550 81664 558622
rect 81624 558544 81676 558550
rect 81624 558486 81676 558492
rect 82924 558414 82952 558855
rect 82912 558408 82964 558414
rect 82818 558376 82874 558385
rect 80060 558340 80112 558346
rect 82912 558350 82964 558356
rect 82818 558311 82874 558320
rect 80060 558282 80112 558288
rect 82832 558074 82860 558311
rect 80704 558068 80756 558074
rect 80704 558010 80756 558016
rect 82820 558068 82872 558074
rect 82820 558010 82872 558016
rect 80716 543318 80744 558010
rect 77576 543312 77628 543318
rect 77576 543254 77628 543260
rect 79324 543312 79376 543318
rect 79324 543254 79376 543260
rect 79692 543312 79744 543318
rect 79692 543254 79744 543260
rect 80704 543312 80756 543318
rect 80704 543254 80756 543260
rect 80796 543312 80848 543318
rect 80796 543254 80848 543260
rect 75486 539974 75868 540002
rect 77588 539988 77616 543254
rect 79704 539988 79732 543254
rect 80808 542910 80836 543254
rect 80796 542904 80848 542910
rect 80796 542846 80848 542852
rect 83832 542632 83884 542638
rect 83832 542574 83884 542580
rect 81716 542564 81768 542570
rect 81716 542506 81768 542512
rect 81728 539988 81756 542506
rect 83844 539988 83872 542574
rect 84212 542570 84240 558855
rect 84290 558784 84346 558793
rect 84290 558719 84346 558728
rect 84304 558618 84332 558719
rect 84292 558612 84344 558618
rect 84292 558554 84344 558560
rect 85408 558482 85436 558855
rect 85396 558476 85448 558482
rect 85396 558418 85448 558424
rect 85684 542638 85712 558855
rect 85672 542632 85724 542638
rect 85672 542574 85724 542580
rect 84200 542564 84252 542570
rect 84200 542506 84252 542512
rect 86236 540002 86264 558855
rect 87602 558855 87658 558864
rect 88982 558920 89038 558929
rect 88982 558855 89038 558864
rect 89626 558920 89682 558929
rect 89626 558855 89682 558864
rect 90086 558920 90142 558929
rect 91374 558920 91430 558929
rect 90086 558855 90088 558864
rect 86868 558826 86920 558832
rect 86880 558793 86908 558826
rect 86866 558784 86922 558793
rect 86866 558719 86922 558728
rect 86880 558550 86908 558719
rect 86868 558544 86920 558550
rect 86868 558486 86920 558492
rect 85882 539974 86264 540002
rect 87616 540002 87644 558855
rect 87880 558816 87932 558822
rect 87878 558784 87880 558793
rect 87932 558784 87934 558793
rect 88996 558754 89024 558855
rect 87878 558719 87934 558728
rect 88984 558748 89036 558754
rect 87892 558278 87920 558719
rect 88984 558690 89036 558696
rect 88996 558346 89024 558690
rect 88984 558340 89036 558346
rect 88984 558282 89036 558288
rect 87880 558272 87932 558278
rect 87880 558214 87932 558220
rect 89640 542450 89668 558855
rect 90140 558855 90142 558864
rect 91008 558884 91060 558890
rect 90088 558826 90140 558832
rect 91374 558855 91430 558864
rect 92478 558920 92534 558929
rect 92478 558855 92534 558864
rect 93582 558920 93638 558929
rect 93582 558855 93638 558864
rect 94594 558920 94650 558929
rect 94594 558855 94650 558864
rect 95330 558920 95386 558929
rect 95330 558855 95386 558864
rect 96618 558920 96674 558929
rect 96618 558855 96674 558864
rect 98274 558920 98330 558929
rect 98274 558855 98330 558864
rect 99562 558920 99618 558929
rect 99562 558855 99618 558864
rect 100666 558920 100722 558929
rect 100666 558855 100722 558864
rect 101954 558920 102010 558929
rect 101954 558855 102010 558864
rect 102690 558920 102746 558929
rect 102690 558855 102746 558864
rect 103426 558920 103482 558929
rect 103426 558855 103482 558864
rect 103978 558920 104034 558929
rect 103978 558855 104034 558864
rect 104806 558920 104862 558929
rect 104806 558855 104862 558864
rect 105358 558920 105414 558929
rect 105358 558855 105414 558864
rect 106186 558920 106242 558929
rect 106186 558855 106242 558864
rect 107566 558920 107622 558929
rect 107566 558855 107622 558864
rect 107842 558920 107898 558929
rect 107842 558855 107898 558864
rect 108946 558920 109002 558929
rect 108946 558855 109002 558864
rect 110326 558920 110382 558929
rect 110326 558855 110382 558864
rect 91008 558826 91060 558832
rect 91020 558278 91048 558826
rect 91388 558686 91416 558855
rect 91376 558680 91428 558686
rect 91376 558622 91428 558628
rect 92492 558414 92520 558855
rect 93596 558618 93624 558855
rect 93584 558612 93636 558618
rect 93584 558554 93636 558560
rect 92480 558408 92532 558414
rect 92480 558350 92532 558356
rect 91008 558272 91060 558278
rect 91008 558214 91060 558220
rect 93596 557870 93624 558554
rect 94608 558482 94636 558855
rect 95344 558686 95372 558855
rect 96632 558822 96660 558855
rect 96620 558816 96672 558822
rect 96620 558758 96672 558764
rect 95332 558680 95384 558686
rect 95332 558622 95384 558628
rect 95344 558550 95372 558622
rect 96632 558550 96660 558758
rect 95332 558544 95384 558550
rect 95332 558486 95384 558492
rect 96620 558544 96672 558550
rect 96620 558486 96672 558492
rect 94596 558476 94648 558482
rect 94596 558418 94648 558424
rect 98288 558346 98316 558855
rect 98276 558340 98328 558346
rect 98276 558282 98328 558288
rect 99576 558278 99604 558855
rect 100298 558784 100354 558793
rect 100298 558719 100300 558728
rect 100352 558719 100354 558728
rect 100300 558690 100352 558696
rect 99564 558272 99616 558278
rect 99564 558214 99616 558220
rect 100312 558006 100340 558690
rect 100300 558000 100352 558006
rect 100300 557942 100352 557948
rect 93584 557864 93636 557870
rect 93584 557806 93636 557812
rect 93674 557696 93730 557705
rect 93674 557631 93730 557640
rect 91006 557560 91062 557569
rect 91006 557495 91062 557504
rect 92386 557560 92442 557569
rect 92386 557495 92442 557504
rect 91020 542910 91048 557495
rect 92400 542910 92428 557495
rect 91008 542904 91060 542910
rect 91008 542846 91060 542852
rect 92112 542904 92164 542910
rect 92112 542846 92164 542852
rect 92388 542904 92440 542910
rect 92388 542846 92440 542852
rect 89640 542422 89760 542450
rect 89732 540002 89760 542422
rect 87616 539974 87998 540002
rect 89732 539974 90022 540002
rect 92124 539988 92152 542846
rect 93688 542842 93716 557631
rect 93766 557560 93822 557569
rect 93766 557495 93822 557504
rect 95146 557560 95202 557569
rect 95146 557495 95202 557504
rect 96526 557560 96582 557569
rect 96526 557495 96582 557504
rect 97906 557560 97962 557569
rect 97906 557495 97962 557504
rect 99286 557560 99342 557569
rect 99286 557495 99342 557504
rect 93676 542836 93728 542842
rect 93676 542778 93728 542784
rect 93780 542774 93808 557495
rect 94136 542904 94188 542910
rect 94136 542846 94188 542852
rect 93768 542768 93820 542774
rect 93768 542710 93820 542716
rect 94148 539988 94176 542846
rect 95160 542502 95188 557495
rect 96252 542836 96304 542842
rect 96252 542778 96304 542784
rect 95148 542496 95200 542502
rect 95148 542438 95200 542444
rect 96264 539988 96292 542778
rect 96540 542706 96568 557495
rect 96528 542700 96580 542706
rect 96528 542642 96580 542648
rect 97920 542638 97948 557495
rect 99300 542842 99328 557495
rect 100680 542910 100708 558855
rect 101862 558648 101918 558657
rect 101862 558583 101918 558592
rect 100760 558408 100812 558414
rect 100760 558350 100812 558356
rect 100772 558074 100800 558350
rect 101876 558074 101904 558583
rect 100760 558068 100812 558074
rect 100760 558010 100812 558016
rect 101864 558068 101916 558074
rect 101864 558010 101916 558016
rect 100668 542904 100720 542910
rect 100668 542846 100720 542852
rect 99288 542836 99340 542842
rect 99288 542778 99340 542784
rect 98368 542768 98420 542774
rect 98368 542710 98420 542716
rect 97908 542632 97960 542638
rect 97908 542574 97960 542580
rect 98380 539988 98408 542710
rect 101968 542502 101996 558855
rect 102046 558784 102102 558793
rect 102046 558719 102102 558728
rect 100392 542496 100444 542502
rect 100392 542438 100444 542444
rect 101956 542496 102008 542502
rect 101956 542438 102008 542444
rect 100404 539988 100432 542438
rect 102060 542434 102088 558719
rect 102704 557870 102732 558855
rect 102692 557864 102744 557870
rect 102692 557806 102744 557812
rect 102508 542700 102560 542706
rect 102508 542642 102560 542648
rect 102048 542428 102100 542434
rect 102048 542370 102100 542376
rect 102520 539988 102548 542642
rect 103440 542638 103468 558855
rect 103992 558482 104020 558855
rect 103980 558476 104032 558482
rect 103980 558418 104032 558424
rect 104716 558476 104768 558482
rect 104716 558418 104768 558424
rect 104728 557666 104756 558418
rect 104716 557660 104768 557666
rect 104716 557602 104768 557608
rect 104532 542700 104584 542706
rect 104532 542642 104584 542648
rect 103428 542632 103480 542638
rect 103428 542574 103480 542580
rect 104544 539988 104572 542642
rect 104820 542570 104848 558855
rect 105372 558686 105400 558855
rect 105360 558680 105412 558686
rect 105360 558622 105412 558628
rect 106096 558680 106148 558686
rect 106096 558622 106148 558628
rect 106108 557802 106136 558622
rect 106096 557796 106148 557802
rect 106096 557738 106148 557744
rect 106200 542706 106228 558855
rect 106278 558784 106334 558793
rect 106278 558719 106334 558728
rect 106292 558550 106320 558719
rect 106280 558544 106332 558550
rect 106280 558486 106332 558492
rect 107476 558544 107528 558550
rect 107476 558486 107528 558492
rect 107488 557734 107516 558486
rect 107476 557728 107528 557734
rect 107476 557670 107528 557676
rect 106648 542836 106700 542842
rect 106648 542778 106700 542784
rect 106188 542700 106240 542706
rect 106188 542642 106240 542648
rect 104808 542564 104860 542570
rect 104808 542506 104860 542512
rect 106660 539988 106688 542778
rect 107580 542774 107608 558855
rect 107856 558550 107884 558855
rect 108578 558784 108634 558793
rect 108578 558719 108634 558728
rect 108592 558618 108620 558719
rect 108580 558612 108632 558618
rect 108580 558554 108632 558560
rect 107844 558544 107896 558550
rect 107844 558486 107896 558492
rect 107856 558346 107884 558486
rect 107844 558340 107896 558346
rect 107844 558282 107896 558288
rect 108592 558278 108620 558554
rect 108580 558272 108632 558278
rect 108580 558214 108632 558220
rect 108960 542910 108988 558855
rect 108672 542904 108724 542910
rect 108672 542846 108724 542852
rect 108948 542904 109000 542910
rect 108948 542846 109000 542852
rect 107568 542768 107620 542774
rect 107568 542710 107620 542716
rect 108684 539988 108712 542846
rect 110340 542842 110368 558855
rect 128268 558136 128320 558142
rect 128268 558078 128320 558084
rect 128280 542910 128308 558078
rect 123208 542904 123260 542910
rect 123208 542846 123260 542852
rect 127348 542904 127400 542910
rect 127348 542846 127400 542852
rect 128268 542904 128320 542910
rect 128268 542846 128320 542852
rect 129464 542904 129516 542910
rect 129464 542846 129516 542852
rect 110328 542836 110380 542842
rect 110328 542778 110380 542784
rect 121184 542768 121236 542774
rect 121184 542710 121236 542716
rect 119068 542700 119120 542706
rect 119068 542642 119120 542648
rect 114928 542632 114980 542638
rect 114928 542574 114980 542580
rect 112812 542496 112864 542502
rect 112812 542438 112864 542444
rect 110788 542428 110840 542434
rect 110788 542370 110840 542376
rect 110800 539988 110828 542370
rect 112824 539988 112852 542438
rect 114940 539988 114968 542574
rect 117044 542564 117096 542570
rect 117044 542506 117096 542512
rect 117056 539988 117084 542506
rect 119080 539988 119108 542642
rect 121196 539988 121224 542710
rect 123220 539988 123248 542846
rect 125324 542836 125376 542842
rect 125324 542778 125376 542784
rect 125336 539988 125364 542778
rect 127360 539988 127388 542846
rect 129476 539988 129504 542846
rect 131488 542836 131540 542842
rect 131488 542778 131540 542784
rect 131500 539988 131528 542778
rect 135720 542700 135772 542706
rect 135720 542642 135772 542648
rect 133604 542564 133656 542570
rect 133604 542506 133656 542512
rect 133616 539988 133644 542506
rect 135732 539988 135760 542642
rect 137296 540326 137324 700198
rect 137848 700126 137876 703520
rect 154132 700194 154160 703520
rect 170324 703474 170352 703520
rect 170140 703446 170352 703474
rect 154120 700188 154172 700194
rect 154120 700130 154172 700136
rect 137836 700120 137888 700126
rect 137836 700062 137888 700068
rect 170140 698306 170168 703446
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 218992 700942 219020 703520
rect 218980 700936 219032 700942
rect 218980 700878 219032 700884
rect 235184 700262 235212 703520
rect 267660 700874 267688 703520
rect 267648 700868 267700 700874
rect 267648 700810 267700 700816
rect 283852 700806 283880 703520
rect 283840 700800 283892 700806
rect 283840 700742 283892 700748
rect 235172 700256 235224 700262
rect 235172 700198 235224 700204
rect 170048 698278 170168 698306
rect 154486 697232 154542 697241
rect 154486 697167 154542 697176
rect 166908 697196 166960 697202
rect 154500 697134 154528 697167
rect 166908 697138 166960 697144
rect 147588 697128 147640 697134
rect 147586 697096 147588 697105
rect 154488 697128 154540 697134
rect 147640 697096 147642 697105
rect 166920 697105 166948 697138
rect 154488 697070 154540 697076
rect 166906 697096 166962 697105
rect 147586 697031 147642 697040
rect 166906 697031 166962 697040
rect 170048 695502 170076 698278
rect 172426 697232 172482 697241
rect 172426 697167 172428 697176
rect 172480 697167 172482 697176
rect 193126 697232 193182 697241
rect 193126 697167 193182 697176
rect 212446 697232 212502 697241
rect 212446 697167 212502 697176
rect 231766 697232 231822 697241
rect 231766 697167 231822 697176
rect 251086 697232 251142 697241
rect 251086 697167 251142 697176
rect 270406 697232 270462 697241
rect 270406 697167 270462 697176
rect 289726 697232 289782 697241
rect 289726 697167 289782 697176
rect 172428 697138 172480 697144
rect 193140 697134 193168 697167
rect 212460 697134 212488 697167
rect 231780 697134 231808 697167
rect 251100 697134 251128 697167
rect 270420 697134 270448 697167
rect 289740 697134 289768 697167
rect 186228 697128 186280 697134
rect 186226 697096 186228 697105
rect 193128 697128 193180 697134
rect 186280 697096 186282 697105
rect 205548 697128 205600 697134
rect 193128 697070 193180 697076
rect 205546 697096 205548 697105
rect 212448 697128 212500 697134
rect 205600 697096 205602 697105
rect 186226 697031 186282 697040
rect 224868 697128 224920 697134
rect 212448 697070 212500 697076
rect 224866 697096 224868 697105
rect 231768 697128 231820 697134
rect 224920 697096 224922 697105
rect 205546 697031 205602 697040
rect 244188 697128 244240 697134
rect 231768 697070 231820 697076
rect 244186 697096 244188 697105
rect 251088 697128 251140 697134
rect 244240 697096 244242 697105
rect 224866 697031 224922 697040
rect 263508 697128 263560 697134
rect 251088 697070 251140 697076
rect 263506 697096 263508 697105
rect 270408 697128 270460 697134
rect 263560 697096 263562 697105
rect 244186 697031 244242 697040
rect 282828 697128 282880 697134
rect 270408 697070 270460 697076
rect 282826 697096 282828 697105
rect 289728 697128 289780 697134
rect 282880 697096 282882 697105
rect 263506 697031 263562 697040
rect 289728 697070 289780 697076
rect 282826 697031 282882 697040
rect 169760 695496 169812 695502
rect 169760 695438 169812 695444
rect 170036 695496 170088 695502
rect 170036 695438 170088 695444
rect 166906 686352 166962 686361
rect 167090 686352 167146 686361
rect 166962 686310 167090 686338
rect 166906 686287 166962 686296
rect 167090 686287 167146 686296
rect 154578 686216 154634 686225
rect 154578 686151 154580 686160
rect 154632 686151 154634 686160
rect 162216 686180 162268 686186
rect 154580 686122 154632 686128
rect 162216 686122 162268 686128
rect 162228 685953 162256 686122
rect 162214 685944 162270 685953
rect 169772 685914 169800 695438
rect 188342 686488 188398 686497
rect 188342 686423 188398 686432
rect 173898 686352 173954 686361
rect 173898 686287 173900 686296
rect 173952 686287 173954 686296
rect 178776 686316 178828 686322
rect 173900 686258 173952 686264
rect 178776 686258 178828 686264
rect 178788 686225 178816 686258
rect 188356 686225 188384 686423
rect 178774 686216 178830 686225
rect 178774 686151 178830 686160
rect 188342 686216 188398 686225
rect 188342 686151 188398 686160
rect 289818 686216 289874 686225
rect 289818 686151 289820 686160
rect 289872 686151 289874 686160
rect 294512 686180 294564 686186
rect 289820 686122 289872 686128
rect 294512 686122 294564 686128
rect 294524 685953 294552 686122
rect 294510 685944 294566 685953
rect 162214 685879 162270 685888
rect 169760 685908 169812 685914
rect 169760 685850 169812 685856
rect 169944 685908 169996 685914
rect 300136 685914 300164 703520
rect 332520 700738 332548 703520
rect 332508 700732 332560 700738
rect 332508 700674 332560 700680
rect 348804 700670 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365116 703474
rect 348792 700664 348844 700670
rect 348792 700606 348844 700612
rect 365088 698290 365116 703446
rect 397472 700602 397500 703520
rect 397460 700596 397512 700602
rect 397460 700538 397512 700544
rect 413664 700534 413692 703520
rect 429856 703474 429884 703520
rect 429856 703446 429976 703474
rect 413652 700528 413704 700534
rect 413652 700470 413704 700476
rect 364432 698284 364484 698290
rect 364432 698226 364484 698232
rect 365076 698284 365128 698290
rect 365076 698226 365128 698232
rect 309046 697232 309102 697241
rect 309046 697167 309102 697176
rect 328366 697232 328422 697241
rect 328366 697167 328422 697176
rect 309060 697134 309088 697167
rect 328380 697134 328408 697167
rect 302148 697128 302200 697134
rect 302146 697096 302148 697105
rect 309048 697128 309100 697134
rect 302200 697096 302202 697105
rect 321468 697128 321520 697134
rect 309048 697070 309100 697076
rect 321466 697096 321468 697105
rect 328368 697128 328420 697134
rect 321520 697096 321522 697105
rect 302146 697031 302202 697040
rect 328368 697070 328420 697076
rect 321466 697031 321522 697040
rect 364444 688650 364472 698226
rect 429948 692850 429976 703446
rect 429200 692844 429252 692850
rect 429200 692786 429252 692792
rect 429936 692844 429988 692850
rect 429936 692786 429988 692792
rect 364352 688622 364472 688650
rect 364352 688514 364380 688622
rect 364352 688486 364472 688514
rect 360106 686352 360162 686361
rect 360290 686352 360346 686361
rect 360162 686310 360290 686338
rect 360106 686287 360162 686296
rect 360290 686287 360346 686296
rect 347778 686216 347834 686225
rect 347778 686151 347780 686160
rect 347832 686151 347834 686160
rect 355416 686180 355468 686186
rect 347780 686122 347832 686128
rect 355416 686122 355468 686128
rect 355428 685953 355456 686122
rect 355414 685944 355470 685953
rect 294510 685879 294566 685888
rect 299572 685908 299624 685914
rect 169944 685850 169996 685856
rect 299572 685850 299624 685856
rect 300124 685908 300176 685914
rect 355414 685879 355470 685888
rect 300124 685850 300176 685856
rect 169956 678994 169984 685850
rect 299584 684486 299612 685850
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 299664 684480 299716 684486
rect 299664 684422 299716 684428
rect 299676 679046 299704 684422
rect 169864 678966 169984 678994
rect 299664 679040 299716 679046
rect 299664 678982 299716 678988
rect 299572 678972 299624 678978
rect 166998 673976 167054 673985
rect 166998 673911 167054 673920
rect 154578 673840 154634 673849
rect 154578 673775 154580 673784
rect 154632 673775 154634 673784
rect 162216 673804 162268 673810
rect 154580 673746 154632 673752
rect 162216 673746 162268 673752
rect 162228 673577 162256 673746
rect 162214 673568 162270 673577
rect 162214 673503 162270 673512
rect 166906 673568 166962 673577
rect 167012 673554 167040 673911
rect 166962 673526 167040 673554
rect 166906 673503 166962 673512
rect 169864 666641 169892 678966
rect 299572 678914 299624 678920
rect 188342 674112 188398 674121
rect 188342 674047 188398 674056
rect 173898 673976 173954 673985
rect 173898 673911 173900 673920
rect 173952 673911 173954 673920
rect 178776 673940 178828 673946
rect 173900 673882 173952 673888
rect 178776 673882 178828 673888
rect 178788 673849 178816 673882
rect 188356 673849 188384 674047
rect 178774 673840 178830 673849
rect 178774 673775 178830 673784
rect 188342 673840 188398 673849
rect 188342 673775 188398 673784
rect 289818 673840 289874 673849
rect 289818 673775 289820 673784
rect 289872 673775 289874 673784
rect 292672 673804 292724 673810
rect 289820 673746 289872 673752
rect 292672 673746 292724 673752
rect 292684 673577 292712 673746
rect 292670 673568 292726 673577
rect 292670 673503 292726 673512
rect 169850 666632 169906 666641
rect 169850 666567 169906 666576
rect 170034 666632 170090 666641
rect 299584 666602 299612 678914
rect 360106 673976 360162 673985
rect 360290 673976 360346 673985
rect 360162 673934 360290 673962
rect 360106 673911 360162 673920
rect 360290 673911 360346 673920
rect 347778 673840 347834 673849
rect 347778 673775 347780 673784
rect 347832 673775 347834 673784
rect 355416 673804 355468 673810
rect 347780 673746 347832 673752
rect 355416 673746 355468 673752
rect 355428 673577 355456 673746
rect 355414 673568 355470 673577
rect 355414 673503 355470 673512
rect 364444 669458 364472 688486
rect 379518 686488 379574 686497
rect 379518 686423 379574 686432
rect 367098 686352 367154 686361
rect 367098 686287 367100 686296
rect 367152 686287 367154 686296
rect 371976 686316 372028 686322
rect 367100 686258 367152 686264
rect 371976 686258 372028 686264
rect 371988 686225 372016 686258
rect 379532 686225 379560 686423
rect 371974 686216 372030 686225
rect 371974 686151 372030 686160
rect 379518 686216 379574 686225
rect 379518 686151 379574 686160
rect 427542 686216 427598 686225
rect 427726 686216 427782 686225
rect 427598 686174 427726 686202
rect 427542 686151 427598 686160
rect 427726 686151 427782 686160
rect 429212 676190 429240 692786
rect 441526 686488 441582 686497
rect 441526 686423 441582 686432
rect 441540 686225 441568 686423
rect 441526 686216 441582 686225
rect 441526 686151 441582 686160
rect 429200 676184 429252 676190
rect 429200 676126 429252 676132
rect 429292 676184 429344 676190
rect 429292 676126 429344 676132
rect 379518 674112 379574 674121
rect 379518 674047 379574 674056
rect 367098 673976 367154 673985
rect 367098 673911 367100 673920
rect 367152 673911 367154 673920
rect 371976 673940 372028 673946
rect 367100 673882 367152 673888
rect 371976 673882 372028 673888
rect 371988 673849 372016 673882
rect 379532 673849 379560 674047
rect 371974 673840 372030 673849
rect 371974 673775 372030 673784
rect 379518 673840 379574 673849
rect 379518 673775 379574 673784
rect 364432 669452 364484 669458
rect 364432 669394 364484 669400
rect 364432 669316 364484 669322
rect 364432 669258 364484 669264
rect 170034 666567 170090 666576
rect 299572 666596 299624 666602
rect 170048 659734 170076 666567
rect 299572 666538 299624 666544
rect 299756 666596 299808 666602
rect 299756 666538 299808 666544
rect 299768 659734 299796 666538
rect 170036 659728 170088 659734
rect 170036 659670 170088 659676
rect 299756 659728 299808 659734
rect 299756 659670 299808 659676
rect 364444 659682 364472 669258
rect 429304 666602 429332 676126
rect 429292 666596 429344 666602
rect 429292 666538 429344 666544
rect 429384 666596 429436 666602
rect 429384 666538 429436 666544
rect 429396 659734 429424 666538
rect 429384 659728 429436 659734
rect 169944 659660 169996 659666
rect 169944 659602 169996 659608
rect 299572 659660 299624 659666
rect 364444 659654 364564 659682
rect 429384 659670 429436 659676
rect 299572 659602 299624 659608
rect 169956 655518 169984 659602
rect 169760 655512 169812 655518
rect 169760 655454 169812 655460
rect 169944 655512 169996 655518
rect 169944 655454 169996 655460
rect 139584 652792 139636 652798
rect 139584 652734 139636 652740
rect 139400 650412 139452 650418
rect 139400 650354 139452 650360
rect 139412 649913 139440 650354
rect 139398 649904 139454 649913
rect 139398 649839 139454 649848
rect 139596 649754 139624 652734
rect 139412 649726 139624 649754
rect 137928 643136 137980 643142
rect 137928 643078 137980 643084
rect 137284 540320 137336 540326
rect 137284 540262 137336 540268
rect 137940 540002 137968 643078
rect 139412 589665 139440 649726
rect 169772 645969 169800 655454
rect 259182 652896 259238 652905
rect 259182 652831 259238 652840
rect 263782 652896 263838 652905
rect 263782 652831 263838 652840
rect 259196 652798 259224 652831
rect 263796 652798 263824 652831
rect 259184 652792 259236 652798
rect 259184 652734 259236 652740
rect 263784 652792 263836 652798
rect 263784 652734 263836 652740
rect 269120 652792 269172 652798
rect 269120 652734 269172 652740
rect 266360 650412 266412 650418
rect 266360 650354 266412 650360
rect 266372 650078 266400 650354
rect 266360 650072 266412 650078
rect 266360 650014 266412 650020
rect 266372 649890 266400 650014
rect 266450 649904 266506 649913
rect 266372 649862 266450 649890
rect 266450 649839 266506 649848
rect 187698 646232 187754 646241
rect 187698 646167 187754 646176
rect 169758 645960 169814 645969
rect 142068 645924 142120 645930
rect 169758 645895 169814 645904
rect 170034 645960 170090 645969
rect 187712 645930 187740 646167
rect 170034 645895 170090 645904
rect 187700 645924 187752 645930
rect 142068 645866 142120 645872
rect 140688 644496 140740 644502
rect 140688 644438 140740 644444
rect 139398 589656 139454 589665
rect 139398 589591 139454 589600
rect 140700 542774 140728 644438
rect 139860 542768 139912 542774
rect 139860 542710 139912 542716
rect 140688 542768 140740 542774
rect 140688 542710 140740 542716
rect 140780 542768 140832 542774
rect 140780 542710 140832 542716
rect 137770 539974 137968 540002
rect 139872 539988 139900 542710
rect 140792 542570 140820 542710
rect 140780 542564 140832 542570
rect 140780 542506 140832 542512
rect 142080 540002 142108 645866
rect 160744 641776 160796 641782
rect 160744 641718 160796 641724
rect 159364 640348 159416 640354
rect 159364 640290 159416 640296
rect 146024 543720 146076 543726
rect 146024 543662 146076 543668
rect 144000 542972 144052 542978
rect 144000 542914 144052 542920
rect 141910 539974 142108 540002
rect 144012 539988 144040 542914
rect 146036 539988 146064 543662
rect 148140 543652 148192 543658
rect 148140 543594 148192 543600
rect 148152 539988 148180 543594
rect 150164 543584 150216 543590
rect 150164 543526 150216 543532
rect 150176 539988 150204 543526
rect 152280 543516 152332 543522
rect 152280 543458 152332 543464
rect 152292 539988 152320 543458
rect 154396 543448 154448 543454
rect 154396 543390 154448 543396
rect 154408 539988 154436 543390
rect 156420 543380 156472 543386
rect 156420 543322 156472 543328
rect 156432 539988 156460 543322
rect 158534 543008 158590 543017
rect 158534 542943 158590 542952
rect 158548 539988 158576 542943
rect 159376 542774 159404 640290
rect 160560 543516 160612 543522
rect 160560 543458 160612 543464
rect 159364 542768 159416 542774
rect 159364 542710 159416 542716
rect 160572 539988 160600 543458
rect 160756 542706 160784 641718
rect 170048 640642 170076 645895
rect 187700 645866 187752 645872
rect 187698 644872 187754 644881
rect 187698 644807 187754 644816
rect 187712 644502 187740 644807
rect 187700 644496 187752 644502
rect 187700 644438 187752 644444
rect 187698 643240 187754 643249
rect 187698 643175 187754 643184
rect 187712 643142 187740 643175
rect 187700 643136 187752 643142
rect 187700 643078 187752 643084
rect 187698 642016 187754 642025
rect 187698 641951 187754 641960
rect 187712 641782 187740 641951
rect 187700 641776 187752 641782
rect 187700 641718 187752 641724
rect 169956 640614 170076 640642
rect 169956 636274 169984 640614
rect 187698 640384 187754 640393
rect 187698 640319 187700 640328
rect 187752 640319 187754 640328
rect 187700 640290 187752 640296
rect 188342 639296 188398 639305
rect 188342 639231 188398 639240
rect 169668 636268 169720 636274
rect 169668 636210 169720 636216
rect 169944 636268 169996 636274
rect 169944 636210 169996 636216
rect 169680 627978 169708 636210
rect 169668 627972 169720 627978
rect 169668 627914 169720 627920
rect 170036 627972 170088 627978
rect 170036 627914 170088 627920
rect 170048 618322 170076 627914
rect 169852 618316 169904 618322
rect 169852 618258 169904 618264
rect 170036 618316 170088 618322
rect 170036 618258 170088 618264
rect 169864 618202 169892 618258
rect 169864 618174 169984 618202
rect 169956 611454 169984 618174
rect 169944 611448 169996 611454
rect 169944 611390 169996 611396
rect 170036 611244 170088 611250
rect 170036 611186 170088 611192
rect 170048 599010 170076 611186
rect 169852 599004 169904 599010
rect 169852 598946 169904 598952
rect 170036 599004 170088 599010
rect 170036 598946 170088 598952
rect 169864 598890 169892 598946
rect 169864 598862 169984 598890
rect 169956 592142 169984 598862
rect 169944 592136 169996 592142
rect 169944 592078 169996 592084
rect 170036 591932 170088 591938
rect 170036 591874 170088 591880
rect 170048 587897 170076 591874
rect 170034 587888 170090 587897
rect 170034 587823 170090 587832
rect 170310 587888 170366 587897
rect 170310 587823 170366 587832
rect 170324 578270 170352 587823
rect 187698 579728 187754 579737
rect 177948 579692 178000 579698
rect 187698 579663 187700 579672
rect 177948 579634 178000 579640
rect 187752 579663 187754 579672
rect 187700 579634 187752 579640
rect 170128 578264 170180 578270
rect 170128 578206 170180 578212
rect 170312 578264 170364 578270
rect 170312 578206 170364 578212
rect 170140 572762 170168 578206
rect 170128 572756 170180 572762
rect 170128 572698 170180 572704
rect 170128 572620 170180 572626
rect 170128 572562 170180 572568
rect 170140 563174 170168 572562
rect 170128 563168 170180 563174
rect 170128 563110 170180 563116
rect 170036 563032 170088 563038
rect 170036 562974 170088 562980
rect 166908 558476 166960 558482
rect 166908 558418 166960 558424
rect 165528 558408 165580 558414
rect 165528 558350 165580 558356
rect 162768 558340 162820 558346
rect 162768 558282 162820 558288
rect 161388 558272 161440 558278
rect 161388 558214 161440 558220
rect 161400 543522 161428 558214
rect 161388 543516 161440 543522
rect 161388 543458 161440 543464
rect 160744 542700 160796 542706
rect 160744 542642 160796 542648
rect 162780 540002 162808 558282
rect 165540 543590 165568 558350
rect 164700 543584 164752 543590
rect 164700 543526 164752 543532
rect 165528 543584 165580 543590
rect 165528 543526 165580 543532
rect 162702 539974 162808 540002
rect 164712 539988 164740 543526
rect 166920 540002 166948 558418
rect 170048 553450 170076 562974
rect 169852 553444 169904 553450
rect 169852 553386 169904 553392
rect 170036 553444 170088 553450
rect 170036 553386 170088 553392
rect 169864 553330 169892 553386
rect 169864 553302 169984 553330
rect 169956 543810 169984 553302
rect 169956 543782 170076 543810
rect 168840 543312 168892 543318
rect 168840 543254 168892 543260
rect 166842 539974 166948 540002
rect 168852 539988 168880 543254
rect 170048 540258 170076 543782
rect 177960 543590 177988 579634
rect 177212 543584 177264 543590
rect 177212 543526 177264 543532
rect 177948 543584 178000 543590
rect 177948 543526 178000 543532
rect 170956 543244 171008 543250
rect 170956 543186 171008 543192
rect 170036 540252 170088 540258
rect 170036 540194 170088 540200
rect 170968 539988 170996 543186
rect 173072 543176 173124 543182
rect 173072 543118 173124 543124
rect 173084 539988 173112 543118
rect 175096 543108 175148 543114
rect 175096 543050 175148 543056
rect 175108 539988 175136 543050
rect 177224 539988 177252 543526
rect 187516 543244 187568 543250
rect 187516 543186 187568 543192
rect 185492 543176 185544 543182
rect 185492 543118 185544 543124
rect 183376 543108 183428 543114
rect 183376 543050 183428 543056
rect 179236 543040 179288 543046
rect 179236 542982 179288 542988
rect 181352 543040 181404 543046
rect 181352 542982 181404 542988
rect 179248 539988 179276 542982
rect 181364 539988 181392 542982
rect 183388 539988 183416 543050
rect 185504 539988 185532 543118
rect 187528 539988 187556 543186
rect 188356 542842 188384 639231
rect 188434 637664 188490 637673
rect 188434 637599 188490 637608
rect 188448 542910 188476 637599
rect 269132 589393 269160 652734
rect 282000 650412 282052 650418
rect 282000 650354 282052 650360
rect 282012 650078 282040 650354
rect 281540 650072 281592 650078
rect 281540 650014 281592 650020
rect 282000 650072 282052 650078
rect 282000 650014 282052 650020
rect 269118 589384 269174 589393
rect 269118 589319 269174 589328
rect 269132 587761 269160 589319
rect 269118 587752 269174 587761
rect 269118 587687 269174 587696
rect 270038 580952 270094 580961
rect 270038 580887 270094 580896
rect 270052 580310 270080 580887
rect 270040 580304 270092 580310
rect 270040 580246 270092 580252
rect 188986 578368 189042 578377
rect 188986 578303 189042 578312
rect 189000 560930 189028 578303
rect 188988 560924 189040 560930
rect 188988 560866 189040 560872
rect 211066 560008 211122 560017
rect 211066 559943 211122 559952
rect 210422 559872 210478 559881
rect 210422 559807 210478 559816
rect 193770 558920 193826 558929
rect 193770 558855 193826 558864
rect 202786 558920 202842 558929
rect 202786 558855 202842 558864
rect 204166 558920 204222 558929
rect 204166 558855 204222 558864
rect 205546 558920 205602 558929
rect 205546 558855 205602 558864
rect 193784 558210 193812 558855
rect 195978 558784 196034 558793
rect 195978 558719 196034 558728
rect 201498 558784 201554 558793
rect 201498 558719 201554 558728
rect 202142 558784 202198 558793
rect 202142 558719 202198 558728
rect 193772 558204 193824 558210
rect 193772 558146 193824 558152
rect 195992 558142 196020 558719
rect 197358 558648 197414 558657
rect 197358 558583 197414 558592
rect 197372 558278 197400 558583
rect 198738 558512 198794 558521
rect 198738 558447 198794 558456
rect 200210 558512 200266 558521
rect 201512 558482 201540 558719
rect 200210 558447 200266 558456
rect 201500 558476 201552 558482
rect 198752 558346 198780 558447
rect 200224 558414 200252 558447
rect 201500 558418 201552 558424
rect 200212 558408 200264 558414
rect 200212 558350 200264 558356
rect 198740 558340 198792 558346
rect 198740 558282 198792 558288
rect 197360 558272 197412 558278
rect 197360 558214 197412 558220
rect 195980 558136 196032 558142
rect 195980 558078 196032 558084
rect 198740 558068 198792 558074
rect 198740 558010 198792 558016
rect 197360 558000 197412 558006
rect 197360 557942 197412 557948
rect 193772 543516 193824 543522
rect 193772 543458 193824 543464
rect 189632 543380 189684 543386
rect 189632 543322 189684 543328
rect 188436 542904 188488 542910
rect 188436 542846 188488 542852
rect 188344 542836 188396 542842
rect 188344 542778 188396 542784
rect 189644 539988 189672 543322
rect 191748 543312 191800 543318
rect 191748 543254 191800 543260
rect 191760 539988 191788 543254
rect 193784 539988 193812 543458
rect 195888 543448 195940 543454
rect 195888 543390 195940 543396
rect 195900 539988 195928 543390
rect 197372 539866 197400 557942
rect 198752 539866 198780 558010
rect 202156 557938 202184 558719
rect 202144 557932 202196 557938
rect 202144 557874 202196 557880
rect 201500 557864 201552 557870
rect 201500 557806 201552 557812
rect 201512 539866 201540 557806
rect 202156 543046 202184 557874
rect 202800 543046 202828 558855
rect 203522 558648 203578 558657
rect 203522 558583 203578 558592
rect 203536 557870 203564 558583
rect 203524 557864 203576 557870
rect 203524 557806 203576 557812
rect 202880 557660 202932 557666
rect 202880 557602 202932 557608
rect 202144 543040 202196 543046
rect 202144 542982 202196 542988
rect 202788 543040 202840 543046
rect 202788 542982 202840 542988
rect 202892 540138 202920 557602
rect 203536 543114 203564 557806
rect 203524 543108 203576 543114
rect 203524 543050 203576 543056
rect 204180 542978 204208 558855
rect 204902 558784 204958 558793
rect 204902 558719 204958 558728
rect 204916 558142 204944 558719
rect 204904 558136 204956 558142
rect 204904 558078 204956 558084
rect 204916 543182 204944 558078
rect 205560 543658 205588 558855
rect 209042 558648 209098 558657
rect 209042 558583 209098 558592
rect 206282 558104 206338 558113
rect 206282 558039 206284 558048
rect 206336 558039 206338 558048
rect 206284 558010 206336 558016
rect 205640 557796 205692 557802
rect 205640 557738 205692 557744
rect 205548 543652 205600 543658
rect 205548 543594 205600 543600
rect 204904 543176 204956 543182
rect 204904 543118 204956 543124
rect 204168 542972 204220 542978
rect 204168 542914 204220 542920
rect 202892 540110 203840 540138
rect 203812 540002 203840 540110
rect 203812 539974 204194 540002
rect 205652 539866 205680 557738
rect 206296 543250 206324 558010
rect 207676 557734 207704 557765
rect 207020 557728 207072 557734
rect 207664 557728 207716 557734
rect 207020 557670 207072 557676
rect 207662 557696 207664 557705
rect 207716 557696 207718 557705
rect 206926 557560 206982 557569
rect 206926 557495 206982 557504
rect 206940 543726 206968 557495
rect 206928 543720 206980 543726
rect 206928 543662 206980 543668
rect 206284 543244 206336 543250
rect 206284 543186 206336 543192
rect 207032 540138 207060 557670
rect 209056 557666 209084 558583
rect 209780 558544 209832 558550
rect 209780 558486 209832 558492
rect 209228 558000 209280 558006
rect 209228 557942 209280 557948
rect 209240 557705 209268 557942
rect 209226 557696 209282 557705
rect 207662 557631 207718 557640
rect 209044 557660 209096 557666
rect 207676 543386 207704 557631
rect 209226 557631 209282 557640
rect 209044 557602 209096 557608
rect 208306 557560 208362 557569
rect 208306 557495 208362 557504
rect 208320 543590 208348 557495
rect 208308 543584 208360 543590
rect 208308 543526 208360 543532
rect 209056 543522 209084 557602
rect 209044 543516 209096 543522
rect 209044 543458 209096 543464
rect 207664 543380 207716 543386
rect 207664 543322 207716 543328
rect 209240 543318 209268 557631
rect 209686 557560 209742 557569
rect 209686 557495 209742 557504
rect 209700 543522 209728 557495
rect 209688 543516 209740 543522
rect 209688 543458 209740 543464
rect 209228 543312 209280 543318
rect 209228 543254 209280 543260
rect 207032 540110 207888 540138
rect 207860 540002 207888 540110
rect 207860 539974 208334 540002
rect 209792 539866 209820 558486
rect 210436 557598 210464 559807
rect 210974 557696 211030 557705
rect 210974 557631 211030 557640
rect 210424 557592 210476 557598
rect 210424 557534 210476 557540
rect 210436 543454 210464 557534
rect 210988 543454 211016 557631
rect 210424 543448 210476 543454
rect 210424 543390 210476 543396
rect 210976 543448 211028 543454
rect 210976 543390 211028 543396
rect 211080 543318 211108 559943
rect 211894 558920 211950 558929
rect 211894 558855 211950 558864
rect 213182 558920 213238 558929
rect 213182 558855 213238 558864
rect 213918 558920 213974 558929
rect 213918 558855 213974 558864
rect 216586 558920 216642 558929
rect 216586 558855 216642 558864
rect 217598 558920 217654 558929
rect 217598 558855 217654 558864
rect 217874 558920 217930 558929
rect 217874 558855 217930 558864
rect 218886 558920 218942 558929
rect 218886 558855 218942 558864
rect 219346 558920 219402 558929
rect 219346 558855 219402 558864
rect 220082 558920 220138 558929
rect 220082 558855 220138 558864
rect 220726 558920 220782 558929
rect 220726 558855 220782 558864
rect 221094 558920 221150 558929
rect 221094 558855 221150 558864
rect 222106 558920 222162 558929
rect 222106 558855 222162 558864
rect 222290 558920 222346 558929
rect 222290 558855 222346 558864
rect 223486 558920 223542 558929
rect 223486 558855 223542 558864
rect 224866 558920 224922 558929
rect 224866 558855 224922 558864
rect 225786 558920 225842 558929
rect 225786 558855 225842 558864
rect 226246 558920 226302 558929
rect 226246 558855 226302 558864
rect 227166 558920 227222 558929
rect 227166 558855 227222 558864
rect 227626 558920 227682 558929
rect 227626 558855 227682 558864
rect 229006 558920 229062 558929
rect 229006 558855 229062 558864
rect 229466 558920 229522 558929
rect 229466 558855 229522 558864
rect 230386 558920 230442 558929
rect 230386 558855 230442 558864
rect 231766 558920 231822 558929
rect 231766 558855 231822 558864
rect 231950 558920 232006 558929
rect 231950 558855 232006 558864
rect 233146 558920 233202 558929
rect 233146 558855 233202 558864
rect 234526 558920 234582 558929
rect 234526 558855 234582 558864
rect 235906 558920 235962 558929
rect 235906 558855 235962 558864
rect 237286 558920 237342 558929
rect 237286 558855 237342 558864
rect 240046 558920 240102 558929
rect 240046 558855 240102 558864
rect 211344 558612 211396 558618
rect 211344 558554 211396 558560
rect 211160 558544 211212 558550
rect 211160 558486 211212 558492
rect 211172 557938 211200 558486
rect 211160 557932 211212 557938
rect 211160 557874 211212 557880
rect 211356 553330 211384 558554
rect 211908 558550 211936 558855
rect 213196 558618 213224 558855
rect 212540 558612 212592 558618
rect 212540 558554 212592 558560
rect 213184 558612 213236 558618
rect 213184 558554 213236 558560
rect 211896 558544 211948 558550
rect 211896 558486 211948 558492
rect 212552 557870 212580 558554
rect 213932 558346 213960 558855
rect 215298 558784 215354 558793
rect 215298 558719 215354 558728
rect 215312 558686 215340 558719
rect 215300 558680 215352 558686
rect 215300 558622 215352 558628
rect 213920 558340 213972 558346
rect 213920 558282 213972 558288
rect 213932 558142 213960 558282
rect 213920 558136 213972 558142
rect 213920 558078 213972 558084
rect 215312 558074 215340 558622
rect 215300 558068 215352 558074
rect 215300 558010 215352 558016
rect 212540 557864 212592 557870
rect 212540 557806 212592 557812
rect 212446 557560 212502 557569
rect 212446 557495 212502 557504
rect 213826 557560 213882 557569
rect 213826 557495 213882 557504
rect 215206 557560 215262 557569
rect 215206 557495 215262 557504
rect 211264 553302 211384 553330
rect 211264 550633 211292 553302
rect 211250 550624 211306 550633
rect 211250 550559 211306 550568
rect 211434 550624 211490 550633
rect 211434 550559 211490 550568
rect 211068 543312 211120 543318
rect 211068 543254 211120 543260
rect 211448 541006 211476 550559
rect 212460 543386 212488 557495
rect 212448 543380 212500 543386
rect 212448 543322 212500 543328
rect 213840 543250 213868 557495
rect 213828 543244 213880 543250
rect 213828 543186 213880 543192
rect 215220 543114 215248 557495
rect 216600 543182 216628 558855
rect 216770 558784 216826 558793
rect 216770 558719 216772 558728
rect 216824 558719 216826 558728
rect 216772 558690 216824 558696
rect 216680 558272 216732 558278
rect 216680 558214 216732 558220
rect 216692 558006 216720 558214
rect 216680 558000 216732 558006
rect 216680 557942 216732 557948
rect 216784 557734 216812 558690
rect 217612 558278 217640 558855
rect 217600 558272 217652 558278
rect 217600 558214 217652 558220
rect 216772 557728 216824 557734
rect 216772 557670 216824 557676
rect 216588 543176 216640 543182
rect 216588 543118 216640 543124
rect 215208 543108 215260 543114
rect 215208 543050 215260 543056
rect 214564 543040 214616 543046
rect 214564 542982 214616 542988
rect 211160 541000 211212 541006
rect 211160 540942 211212 540948
rect 211436 541000 211488 541006
rect 211436 540942 211488 540948
rect 211172 540138 211200 540942
rect 211172 540110 212028 540138
rect 212000 539866 212028 540110
rect 214576 539988 214604 542982
rect 216588 542972 216640 542978
rect 216588 542914 216640 542920
rect 216600 539988 216628 542914
rect 217888 542570 217916 558855
rect 217966 558784 218022 558793
rect 217966 558719 218022 558728
rect 217980 543046 218008 558719
rect 218900 558414 218928 558855
rect 218060 558408 218112 558414
rect 218060 558350 218112 558356
rect 218888 558408 218940 558414
rect 218888 558350 218940 558356
rect 218072 557666 218100 558350
rect 218060 557660 218112 557666
rect 218060 557602 218112 557608
rect 218704 543652 218756 543658
rect 218704 543594 218756 543600
rect 217968 543040 218020 543046
rect 217968 542982 218020 542988
rect 217876 542564 217928 542570
rect 217876 542506 217928 542512
rect 218716 539988 218744 543594
rect 219360 542502 219388 558855
rect 220096 557598 220124 558855
rect 220084 557592 220136 557598
rect 220084 557534 220136 557540
rect 220740 545306 220768 558855
rect 221108 558550 221136 558855
rect 221096 558544 221148 558550
rect 221096 558486 221148 558492
rect 220556 545278 220768 545306
rect 220556 542706 220584 545278
rect 220728 543720 220780 543726
rect 220728 543662 220780 543668
rect 220544 542700 220596 542706
rect 220544 542642 220596 542648
rect 219348 542496 219400 542502
rect 219348 542438 219400 542444
rect 220740 539988 220768 543662
rect 222120 542638 222148 558855
rect 222304 558618 222332 558855
rect 222292 558612 222344 558618
rect 222292 558554 222344 558560
rect 222844 543584 222896 543590
rect 222844 543526 222896 543532
rect 222108 542632 222160 542638
rect 222108 542574 222160 542580
rect 222856 539988 222884 543526
rect 223500 542842 223528 558855
rect 223592 558822 223620 558853
rect 223580 558816 223632 558822
rect 223578 558784 223580 558793
rect 223632 558784 223634 558793
rect 223578 558719 223634 558728
rect 224406 558784 224462 558793
rect 224406 558719 224462 558728
rect 223592 558346 223620 558719
rect 224420 558686 224448 558719
rect 224408 558680 224460 558686
rect 224408 558622 224460 558628
rect 223580 558340 223632 558346
rect 223580 558282 223632 558288
rect 224880 545306 224908 558855
rect 225800 558754 225828 558855
rect 226154 558784 226210 558793
rect 225788 558748 225840 558754
rect 226154 558719 226210 558728
rect 225788 558690 225840 558696
rect 225800 558346 225828 558690
rect 225788 558340 225840 558346
rect 225788 558282 225840 558288
rect 224696 545278 224908 545306
rect 223488 542836 223540 542842
rect 223488 542778 223540 542784
rect 224696 542774 224724 545278
rect 224868 543516 224920 543522
rect 224868 543458 224920 543464
rect 224684 542768 224736 542774
rect 224684 542710 224736 542716
rect 224880 539988 224908 543458
rect 226168 542910 226196 558719
rect 226260 542978 226288 558855
rect 227180 558754 227208 558855
rect 226340 558748 226392 558754
rect 226340 558690 226392 558696
rect 227168 558748 227220 558754
rect 227168 558690 227220 558696
rect 226352 558278 226380 558690
rect 226340 558272 226392 558278
rect 226340 558214 226392 558220
rect 227640 543658 227668 558855
rect 227718 558784 227774 558793
rect 227718 558719 227774 558728
rect 227732 558414 227760 558719
rect 227720 558408 227772 558414
rect 227720 558350 227772 558356
rect 227812 558408 227864 558414
rect 227812 558350 227864 558356
rect 227732 558278 227760 558350
rect 227720 558272 227772 558278
rect 227720 558214 227772 558220
rect 227824 557598 227852 558350
rect 227812 557592 227864 557598
rect 227812 557534 227864 557540
rect 229020 543726 229048 558855
rect 229480 558414 229508 558855
rect 229468 558408 229520 558414
rect 229468 558350 229520 558356
rect 229008 543720 229060 543726
rect 229008 543662 229060 543668
rect 227628 543652 227680 543658
rect 227628 543594 227680 543600
rect 230400 543522 230428 558855
rect 230478 558648 230534 558657
rect 230478 558583 230534 558592
rect 230492 558550 230520 558583
rect 230480 558544 230532 558550
rect 230480 558486 230532 558492
rect 231780 543590 231808 558855
rect 231964 558822 231992 558855
rect 231952 558816 232004 558822
rect 231952 558758 232004 558764
rect 233054 558784 233110 558793
rect 233054 558719 233110 558728
rect 231858 558648 231914 558657
rect 231858 558583 231860 558592
rect 231912 558583 231914 558592
rect 231860 558554 231912 558560
rect 231768 543584 231820 543590
rect 231768 543526 231820 543532
rect 230388 543516 230440 543522
rect 230388 543458 230440 543464
rect 233068 543454 233096 558719
rect 226984 543448 227036 543454
rect 226984 543390 227036 543396
rect 233056 543448 233108 543454
rect 233056 543390 233108 543396
rect 226248 542972 226300 542978
rect 226248 542914 226300 542920
rect 226156 542904 226208 542910
rect 226156 542846 226208 542852
rect 226996 539988 227024 543390
rect 233160 543386 233188 558855
rect 233238 558784 233294 558793
rect 233238 558719 233294 558728
rect 233252 558686 233280 558719
rect 233240 558680 233292 558686
rect 233240 558622 233292 558628
rect 231124 543380 231176 543386
rect 231124 543322 231176 543328
rect 233148 543380 233200 543386
rect 233148 543322 233200 543328
rect 229100 543312 229152 543318
rect 229100 543254 229152 543260
rect 229112 539988 229140 543254
rect 231136 539988 231164 543322
rect 234540 543318 234568 558855
rect 234618 558648 234674 558657
rect 234618 558583 234674 558592
rect 234632 558346 234660 558583
rect 234620 558340 234672 558346
rect 234620 558282 234672 558288
rect 234528 543312 234580 543318
rect 234528 543254 234580 543260
rect 235920 543250 235948 558855
rect 235998 558784 236054 558793
rect 235998 558719 236000 558728
rect 236052 558719 236054 558728
rect 236000 558690 236052 558696
rect 233240 543244 233292 543250
rect 233240 543186 233292 543192
rect 235908 543244 235960 543250
rect 235908 543186 235960 543192
rect 233252 539988 233280 543186
rect 237300 543114 237328 558855
rect 237378 558512 237434 558521
rect 237378 558447 237434 558456
rect 238758 558512 238814 558521
rect 238758 558447 238814 558456
rect 237392 558278 237420 558447
rect 238772 558414 238800 558447
rect 238760 558408 238812 558414
rect 238760 558350 238812 558356
rect 237380 558272 237432 558278
rect 237380 558214 237432 558220
rect 238666 558104 238722 558113
rect 238666 558039 238722 558048
rect 238680 543182 238708 558039
rect 237380 543176 237432 543182
rect 237380 543118 237432 543124
rect 238668 543176 238720 543182
rect 238668 543118 238720 543124
rect 235264 543108 235316 543114
rect 235264 543050 235316 543056
rect 237288 543108 237340 543114
rect 237288 543050 237340 543056
rect 235276 539988 235304 543050
rect 237392 539988 237420 543118
rect 240060 543046 240088 558855
rect 260196 543720 260248 543726
rect 260196 543662 260248 543668
rect 258080 543652 258132 543658
rect 258080 543594 258132 543600
rect 239404 543040 239456 543046
rect 239404 542982 239456 542988
rect 240048 543040 240100 543046
rect 240048 542982 240100 542988
rect 239416 539988 239444 542982
rect 256056 542972 256108 542978
rect 256056 542914 256108 542920
rect 253940 542904 253992 542910
rect 253940 542846 253992 542852
rect 249800 542836 249852 542842
rect 249800 542778 249852 542784
rect 245660 542700 245712 542706
rect 245660 542642 245712 542648
rect 241520 542564 241572 542570
rect 241520 542506 241572 542512
rect 241532 539988 241560 542506
rect 243544 542496 243596 542502
rect 243544 542438 243596 542444
rect 243556 539988 243584 542438
rect 245672 539988 245700 542642
rect 247776 542632 247828 542638
rect 247776 542574 247828 542580
rect 247788 539988 247816 542574
rect 249812 539988 249840 542778
rect 251916 542768 251968 542774
rect 251916 542710 251968 542716
rect 251928 539988 251956 542710
rect 253952 539988 253980 542846
rect 256068 539988 256096 542914
rect 258092 539988 258120 543594
rect 260208 539988 260236 543662
rect 264336 543584 264388 543590
rect 264336 543526 264388 543532
rect 262220 543516 262272 543522
rect 262220 543458 262272 543464
rect 262232 539988 262260 543458
rect 264348 539988 264376 543526
rect 266452 543448 266504 543454
rect 266452 543390 266504 543396
rect 266464 539988 266492 543390
rect 268476 543380 268528 543386
rect 268476 543322 268528 543328
rect 268488 539988 268516 543322
rect 270592 543312 270644 543318
rect 270592 543254 270644 543260
rect 270604 539988 270632 543254
rect 272616 543244 272668 543250
rect 272616 543186 272668 543192
rect 272628 539988 272656 543186
rect 276756 543176 276808 543182
rect 276756 543118 276808 543124
rect 274732 543108 274784 543114
rect 274732 543050 274784 543056
rect 274744 539988 274772 543050
rect 276768 539988 276796 543118
rect 278872 543040 278924 543046
rect 278872 542982 278924 542988
rect 278884 539988 278912 542982
rect 197372 539838 197938 539866
rect 198752 539838 200054 539866
rect 201512 539838 202078 539866
rect 205652 539838 206218 539866
rect 209792 539838 210450 539866
rect 212000 539838 212474 539866
rect 59728 539164 59780 539170
rect 59728 539106 59780 539112
rect 59636 539096 59688 539102
rect 59636 539038 59688 539044
rect 59542 414760 59598 414769
rect 59542 414695 59598 414704
rect 59450 402112 59506 402121
rect 59450 402047 59506 402056
rect 59358 399936 59414 399945
rect 59358 399871 59414 399880
rect 59266 397896 59322 397905
rect 59266 397831 59322 397840
rect 59648 395729 59676 539038
rect 59740 408377 59768 539106
rect 60740 538416 60792 538422
rect 60740 538358 60792 538364
rect 60004 538348 60056 538354
rect 60004 538290 60056 538296
rect 60016 429214 60044 538290
rect 60752 536858 60780 538358
rect 60096 536852 60148 536858
rect 60096 536794 60148 536800
rect 60740 536852 60792 536858
rect 60740 536794 60792 536800
rect 60108 434042 60136 536794
rect 60096 434036 60148 434042
rect 60096 433978 60148 433984
rect 60004 429208 60056 429214
rect 60004 429150 60056 429156
rect 59726 408368 59782 408377
rect 59726 408303 59782 408312
rect 59634 395720 59690 395729
rect 59634 395655 59690 395664
rect 58622 385248 58678 385257
rect 58622 385183 58678 385192
rect 58254 372600 58310 372609
rect 58254 372535 58310 372544
rect 58162 370424 58218 370433
rect 58162 370359 58218 370368
rect 57702 364168 57758 364177
rect 57702 364103 57758 364112
rect 57702 359952 57758 359961
rect 57702 359887 57758 359896
rect 57426 357912 57482 357921
rect 57426 357847 57482 357856
rect 57334 349480 57390 349489
rect 57334 349415 57390 349424
rect 57348 330546 57376 349415
rect 57336 330540 57388 330546
rect 57336 330482 57388 330488
rect 57334 330440 57390 330449
rect 57334 330375 57390 330384
rect 57348 316033 57376 330375
rect 57440 328438 57468 357847
rect 57518 351520 57574 351529
rect 57518 351455 57574 351464
rect 57428 328432 57480 328438
rect 57428 328374 57480 328380
rect 57426 326224 57482 326233
rect 57426 326159 57482 326168
rect 57334 316024 57390 316033
rect 57334 315959 57390 315968
rect 57334 306504 57390 306513
rect 57334 306439 57390 306448
rect 57348 296682 57376 306439
rect 57336 296676 57388 296682
rect 57336 296618 57388 296624
rect 57244 295316 57296 295322
rect 57244 295258 57296 295264
rect 57336 287088 57388 287094
rect 57336 287030 57388 287036
rect 57348 277409 57376 287030
rect 57334 277400 57390 277409
rect 57244 277364 57296 277370
rect 57334 277335 57390 277344
rect 57244 277306 57296 277312
rect 57256 263634 57284 277306
rect 57336 268456 57388 268462
rect 57336 268398 57388 268404
rect 57244 263628 57296 263634
rect 57244 263570 57296 263576
rect 57152 229084 57204 229090
rect 57152 229026 57204 229032
rect 57348 218006 57376 268398
rect 57336 218000 57388 218006
rect 57336 217942 57388 217948
rect 57440 205630 57468 326159
rect 57532 317422 57560 351455
rect 57610 345264 57666 345273
rect 57610 345199 57666 345208
rect 57624 322114 57652 345199
rect 57716 336734 57744 359887
rect 57794 347304 57850 347313
rect 57794 347239 57850 347248
rect 57704 336728 57756 336734
rect 57704 336670 57756 336676
rect 57704 330540 57756 330546
rect 57704 330482 57756 330488
rect 57716 327078 57744 330482
rect 57704 327072 57756 327078
rect 57704 327014 57756 327020
rect 57702 324184 57758 324193
rect 57702 324119 57758 324128
rect 57612 322108 57664 322114
rect 57612 322050 57664 322056
rect 57520 317416 57572 317422
rect 57520 317358 57572 317364
rect 57520 317280 57572 317286
rect 57520 317222 57572 317228
rect 57532 315994 57560 317222
rect 57520 315988 57572 315994
rect 57520 315930 57572 315936
rect 57716 315858 57744 324119
rect 57808 322998 57836 347239
rect 57886 341048 57942 341057
rect 57886 340983 57942 340992
rect 57796 322992 57848 322998
rect 57796 322934 57848 322940
rect 57794 322008 57850 322017
rect 57794 321943 57850 321952
rect 57808 317898 57836 321943
rect 57796 317892 57848 317898
rect 57796 317834 57848 317840
rect 57794 317792 57850 317801
rect 57794 317727 57850 317736
rect 57704 315852 57756 315858
rect 57704 315794 57756 315800
rect 57702 315752 57758 315761
rect 57702 315687 57758 315696
rect 57520 306400 57572 306406
rect 57520 306342 57572 306348
rect 57612 306400 57664 306406
rect 57612 306342 57664 306348
rect 57532 296682 57560 306342
rect 57624 296721 57652 306342
rect 57610 296712 57666 296721
rect 57520 296676 57572 296682
rect 57610 296647 57666 296656
rect 57520 296618 57572 296624
rect 57612 287156 57664 287162
rect 57612 287098 57664 287104
rect 57520 287088 57572 287094
rect 57520 287030 57572 287036
rect 57532 277370 57560 287030
rect 57624 277370 57652 287098
rect 57520 277364 57572 277370
rect 57520 277306 57572 277312
rect 57612 277364 57664 277370
rect 57612 277306 57664 277312
rect 57612 268456 57664 268462
rect 57612 268398 57664 268404
rect 57520 263628 57572 263634
rect 57520 263570 57572 263576
rect 57428 205624 57480 205630
rect 57428 205566 57480 205572
rect 57532 182170 57560 263570
rect 57520 182164 57572 182170
rect 57520 182106 57572 182112
rect 57624 171086 57652 268398
rect 57612 171080 57664 171086
rect 57612 171022 57664 171028
rect 57716 135250 57744 315687
rect 57704 135244 57756 135250
rect 57704 135186 57756 135192
rect 57808 124166 57836 317727
rect 57900 300830 57928 340983
rect 58716 339448 58768 339454
rect 58716 339390 58768 339396
rect 58624 336728 58676 336734
rect 58624 336670 58676 336676
rect 58532 320136 58584 320142
rect 58532 320078 58584 320084
rect 58440 317416 58492 317422
rect 58440 317358 58492 317364
rect 57980 315852 58032 315858
rect 57980 315794 58032 315800
rect 57992 306406 58020 315794
rect 57980 306400 58032 306406
rect 57980 306342 58032 306348
rect 57888 300824 57940 300830
rect 57888 300766 57940 300772
rect 58452 300422 58480 317358
rect 58440 300416 58492 300422
rect 58440 300358 58492 300364
rect 58544 300150 58572 320078
rect 58636 300490 58664 336670
rect 58728 304366 58756 339390
rect 58808 331628 58860 331634
rect 58808 331570 58860 331576
rect 58716 304360 58768 304366
rect 58716 304302 58768 304308
rect 58820 303482 58848 331570
rect 58900 328432 58952 328438
rect 58900 328374 58952 328380
rect 58808 303476 58860 303482
rect 58808 303418 58860 303424
rect 58624 300484 58676 300490
rect 58624 300426 58676 300432
rect 58912 300218 58940 328374
rect 58992 327072 59044 327078
rect 58992 327014 59044 327020
rect 59004 300286 59032 327014
rect 59084 322992 59136 322998
rect 59084 322934 59136 322940
rect 59096 314702 59124 322934
rect 59268 322108 59320 322114
rect 59268 322050 59320 322056
rect 59084 314696 59136 314702
rect 59084 314638 59136 314644
rect 59082 313576 59138 313585
rect 59082 313511 59138 313520
rect 58992 300280 59044 300286
rect 58992 300222 59044 300228
rect 58900 300212 58952 300218
rect 58900 300154 58952 300160
rect 58532 300144 58584 300150
rect 58532 300086 58584 300092
rect 57888 296676 57940 296682
rect 57888 296618 57940 296624
rect 57900 287094 57928 296618
rect 57888 287088 57940 287094
rect 57888 287030 57940 287036
rect 57888 277364 57940 277370
rect 57888 277306 57940 277312
rect 57900 268462 57928 277306
rect 57888 268456 57940 268462
rect 57888 268398 57940 268404
rect 57796 124160 57848 124166
rect 57796 124102 57848 124108
rect 59096 111790 59124 313511
rect 59174 307320 59230 307329
rect 59174 307255 59230 307264
rect 59084 111784 59136 111790
rect 59084 111726 59136 111732
rect 56600 88324 56652 88330
rect 56600 88266 56652 88272
rect 59188 64870 59216 307255
rect 59280 304502 59308 322050
rect 59358 319968 59414 319977
rect 59358 319903 59414 319912
rect 59268 304496 59320 304502
rect 59268 304438 59320 304444
rect 59266 301064 59322 301073
rect 59266 300999 59322 301008
rect 53104 64864 53156 64870
rect 53104 64806 53156 64812
rect 59176 64864 59228 64870
rect 59176 64806 59228 64812
rect 59280 17950 59308 300999
rect 59372 158710 59400 319903
rect 60004 314696 60056 314702
rect 60004 314638 60056 314644
rect 59452 304496 59504 304502
rect 59452 304438 59504 304444
rect 59464 300694 59492 304438
rect 59544 304360 59596 304366
rect 59544 304302 59596 304308
rect 59452 300688 59504 300694
rect 59452 300630 59504 300636
rect 59556 300354 59584 304302
rect 60016 300626 60044 314638
rect 60648 303476 60700 303482
rect 60648 303418 60700 303424
rect 60004 300620 60056 300626
rect 60004 300562 60056 300568
rect 60660 300558 60688 303418
rect 281552 303385 281580 650014
rect 299584 650010 299612 659602
rect 364536 654158 364564 659654
rect 429292 659660 429344 659666
rect 429292 659602 429344 659608
rect 364340 654152 364392 654158
rect 364340 654094 364392 654100
rect 364524 654152 364576 654158
rect 364524 654094 364576 654100
rect 364352 650826 364380 654094
rect 378506 652896 378562 652905
rect 378506 652831 378562 652840
rect 383474 652896 383530 652905
rect 383474 652831 383530 652840
rect 378520 652798 378548 652831
rect 383488 652798 383516 652831
rect 378508 652792 378560 652798
rect 378508 652734 378560 652740
rect 383476 652792 383528 652798
rect 383476 652734 383528 652740
rect 389364 652792 389416 652798
rect 389364 652734 389416 652740
rect 364340 650820 364392 650826
rect 364340 650762 364392 650768
rect 389180 650412 389232 650418
rect 389180 650354 389232 650360
rect 299572 650004 299624 650010
rect 299572 649946 299624 649952
rect 299756 650004 299808 650010
rect 299756 649946 299808 649952
rect 291936 645924 291988 645930
rect 291936 645866 291988 645872
rect 290556 644496 290608 644502
rect 290556 644438 290608 644444
rect 287704 643136 287756 643142
rect 287704 643078 287756 643084
rect 286324 641776 286376 641782
rect 286324 641718 286376 641724
rect 284944 640348 284996 640354
rect 284944 640290 284996 640296
rect 283564 638988 283616 638994
rect 283564 638930 283616 638936
rect 281632 580304 281684 580310
rect 281632 580246 281684 580252
rect 281538 303376 281594 303385
rect 281538 303311 281594 303320
rect 281644 301209 281672 580246
rect 282184 578264 282236 578270
rect 282184 578206 282236 578212
rect 282196 561678 282224 578206
rect 281724 561672 281776 561678
rect 281724 561614 281776 561620
rect 282184 561672 282236 561678
rect 282184 561614 282236 561620
rect 281736 560930 281764 561614
rect 281724 560924 281776 560930
rect 281724 560866 281776 560872
rect 281736 538937 281764 560866
rect 281722 538928 281778 538937
rect 281722 538863 281778 538872
rect 282828 536784 282880 536790
rect 282826 536752 282828 536761
rect 282880 536752 282882 536761
rect 282826 536687 282882 536696
rect 282828 535424 282880 535430
rect 282828 535366 282880 535372
rect 282840 534585 282868 535366
rect 282826 534576 282882 534585
rect 282826 534511 282882 534520
rect 282828 532704 282880 532710
rect 282828 532646 282880 532652
rect 282840 532409 282868 532646
rect 282826 532400 282882 532409
rect 282826 532335 282882 532344
rect 282828 531276 282880 531282
rect 282828 531218 282880 531224
rect 282840 530233 282868 531218
rect 282826 530224 282882 530233
rect 282826 530159 282882 530168
rect 282828 528556 282880 528562
rect 282828 528498 282880 528504
rect 282840 527921 282868 528498
rect 282826 527912 282882 527921
rect 282826 527847 282882 527856
rect 282828 525768 282880 525774
rect 282826 525736 282828 525745
rect 282880 525736 282882 525745
rect 282826 525671 282882 525680
rect 282828 524408 282880 524414
rect 282828 524350 282880 524356
rect 282840 523569 282868 524350
rect 282826 523560 282882 523569
rect 282826 523495 282882 523504
rect 282828 521620 282880 521626
rect 282828 521562 282880 521568
rect 282840 521393 282868 521562
rect 282826 521384 282882 521393
rect 282826 521319 282882 521328
rect 282828 520260 282880 520266
rect 282828 520202 282880 520208
rect 282840 519217 282868 520202
rect 282826 519208 282882 519217
rect 282826 519143 282882 519152
rect 281908 517472 281960 517478
rect 281908 517414 281960 517420
rect 281920 516905 281948 517414
rect 281906 516896 281962 516905
rect 281906 516831 281962 516840
rect 282828 514752 282880 514758
rect 282826 514720 282828 514729
rect 282880 514720 282882 514729
rect 282826 514655 282882 514664
rect 282092 513324 282144 513330
rect 282092 513266 282144 513272
rect 282104 512553 282132 513266
rect 282090 512544 282146 512553
rect 282090 512479 282146 512488
rect 282828 510604 282880 510610
rect 282828 510546 282880 510552
rect 282840 510377 282868 510546
rect 282826 510368 282882 510377
rect 282826 510303 282882 510312
rect 282276 509244 282328 509250
rect 282276 509186 282328 509192
rect 282288 508201 282316 509186
rect 282274 508192 282330 508201
rect 282274 508127 282330 508136
rect 281908 506456 281960 506462
rect 281908 506398 281960 506404
rect 281920 505889 281948 506398
rect 281906 505880 281962 505889
rect 281906 505815 281962 505824
rect 282826 503704 282882 503713
rect 282826 503639 282828 503648
rect 282880 503639 282882 503648
rect 282828 503610 282880 503616
rect 282092 502308 282144 502314
rect 282092 502250 282144 502256
rect 282104 501537 282132 502250
rect 282090 501528 282146 501537
rect 282090 501463 282146 501472
rect 282828 499520 282880 499526
rect 282828 499462 282880 499468
rect 282840 499361 282868 499462
rect 282826 499352 282882 499361
rect 282826 499287 282882 499296
rect 282276 498160 282328 498166
rect 282276 498102 282328 498108
rect 282288 497185 282316 498102
rect 282274 497176 282330 497185
rect 282274 497111 282330 497120
rect 281908 495440 281960 495446
rect 281908 495382 281960 495388
rect 281920 494873 281948 495382
rect 281906 494864 281962 494873
rect 281906 494799 281962 494808
rect 282460 494012 282512 494018
rect 282460 493954 282512 493960
rect 282472 492697 282500 493954
rect 282458 492688 282514 492697
rect 282458 492623 282514 492632
rect 282092 491292 282144 491298
rect 282092 491234 282144 491240
rect 282104 490521 282132 491234
rect 282090 490512 282146 490521
rect 282090 490447 282146 490456
rect 282828 488504 282880 488510
rect 282828 488446 282880 488452
rect 282840 488345 282868 488446
rect 282826 488336 282882 488345
rect 282826 488271 282882 488280
rect 282828 487144 282880 487150
rect 282828 487086 282880 487092
rect 282840 486169 282868 487086
rect 282826 486160 282882 486169
rect 282826 486095 282882 486104
rect 282828 484356 282880 484362
rect 282828 484298 282880 484304
rect 282840 483857 282868 484298
rect 282826 483848 282882 483857
rect 282826 483783 282882 483792
rect 282460 482996 282512 483002
rect 282460 482938 282512 482944
rect 282472 481681 282500 482938
rect 282458 481672 282514 481681
rect 282458 481607 282514 481616
rect 282092 480208 282144 480214
rect 282092 480150 282144 480156
rect 282104 479505 282132 480150
rect 282090 479496 282146 479505
rect 282090 479431 282146 479440
rect 282828 477488 282880 477494
rect 282828 477430 282880 477436
rect 282840 477329 282868 477430
rect 282826 477320 282882 477329
rect 282826 477255 282882 477264
rect 282552 476060 282604 476066
rect 282552 476002 282604 476008
rect 282564 475153 282592 476002
rect 282550 475144 282606 475153
rect 282550 475079 282606 475088
rect 282092 473340 282144 473346
rect 282092 473282 282144 473288
rect 282104 472977 282132 473282
rect 282090 472968 282146 472977
rect 282090 472903 282146 472912
rect 282460 471980 282512 471986
rect 282460 471922 282512 471928
rect 282472 470665 282500 471922
rect 282458 470656 282514 470665
rect 282458 470591 282514 470600
rect 282092 469192 282144 469198
rect 282092 469134 282144 469140
rect 282104 468489 282132 469134
rect 282090 468480 282146 468489
rect 282090 468415 282146 468424
rect 282828 466404 282880 466410
rect 282828 466346 282880 466352
rect 282840 466313 282868 466346
rect 282826 466304 282882 466313
rect 282826 466239 282882 466248
rect 282276 465044 282328 465050
rect 282276 464986 282328 464992
rect 282288 464137 282316 464986
rect 282274 464128 282330 464137
rect 282274 464063 282330 464072
rect 282828 462324 282880 462330
rect 282828 462266 282880 462272
rect 282840 461961 282868 462266
rect 282826 461952 282882 461961
rect 282826 461887 282882 461896
rect 282460 460896 282512 460902
rect 282460 460838 282512 460844
rect 282472 459649 282500 460838
rect 282458 459640 282514 459649
rect 282458 459575 282514 459584
rect 282092 458176 282144 458182
rect 282092 458118 282144 458124
rect 282104 457473 282132 458118
rect 282090 457464 282146 457473
rect 282090 457399 282146 457408
rect 282828 455388 282880 455394
rect 282828 455330 282880 455336
rect 282840 455297 282868 455330
rect 282826 455288 282882 455297
rect 282826 455223 282882 455232
rect 282828 454028 282880 454034
rect 282828 453970 282880 453976
rect 282840 453121 282868 453970
rect 282826 453112 282882 453121
rect 282826 453047 282882 453056
rect 282828 451240 282880 451246
rect 282828 451182 282880 451188
rect 282840 450945 282868 451182
rect 282826 450936 282882 450945
rect 282826 450871 282882 450880
rect 282460 449880 282512 449886
rect 282460 449822 282512 449828
rect 282472 448633 282500 449822
rect 282458 448624 282514 448633
rect 282458 448559 282514 448568
rect 282828 447092 282880 447098
rect 282828 447034 282880 447040
rect 282840 446457 282868 447034
rect 282826 446448 282882 446457
rect 282826 446383 282882 446392
rect 282828 444372 282880 444378
rect 282828 444314 282880 444320
rect 282840 444281 282868 444314
rect 282826 444272 282882 444281
rect 282826 444207 282882 444216
rect 282828 442944 282880 442950
rect 282828 442886 282880 442892
rect 282840 442105 282868 442886
rect 282826 442096 282882 442105
rect 282826 442031 282882 442040
rect 282828 440224 282880 440230
rect 282828 440166 282880 440172
rect 282840 439929 282868 440166
rect 282826 439920 282882 439929
rect 282826 439855 282882 439864
rect 282460 438864 282512 438870
rect 282460 438806 282512 438812
rect 282472 437617 282500 438806
rect 282458 437608 282514 437617
rect 282458 437543 282514 437552
rect 282828 436076 282880 436082
rect 282828 436018 282880 436024
rect 282840 435441 282868 436018
rect 282826 435432 282882 435441
rect 282826 435367 282882 435376
rect 282828 433288 282880 433294
rect 282826 433256 282828 433265
rect 282880 433256 282882 433265
rect 282826 433191 282882 433200
rect 282828 431928 282880 431934
rect 282828 431870 282880 431876
rect 282840 431089 282868 431870
rect 282826 431080 282882 431089
rect 282826 431015 282882 431024
rect 282828 429140 282880 429146
rect 282828 429082 282880 429088
rect 282840 428913 282868 429082
rect 282826 428904 282882 428913
rect 282826 428839 282882 428848
rect 282828 426624 282880 426630
rect 282826 426592 282828 426601
rect 282880 426592 282882 426601
rect 282826 426527 282882 426536
rect 282460 425060 282512 425066
rect 282460 425002 282512 425008
rect 282472 424425 282500 425002
rect 282458 424416 282514 424425
rect 282458 424351 282514 424360
rect 282092 422272 282144 422278
rect 282090 422240 282092 422249
rect 282144 422240 282146 422249
rect 282090 422175 282146 422184
rect 283576 420850 283604 638930
rect 284956 422278 284984 640290
rect 285036 579692 285088 579698
rect 285036 579634 285088 579640
rect 284944 422272 284996 422278
rect 284944 422214 284996 422220
rect 281724 420844 281776 420850
rect 281724 420786 281776 420792
rect 283564 420844 283616 420850
rect 283564 420786 283616 420792
rect 281736 420073 281764 420786
rect 281722 420064 281778 420073
rect 281722 419999 281778 420008
rect 282828 418124 282880 418130
rect 282828 418066 282880 418072
rect 282840 417897 282868 418066
rect 282826 417888 282882 417897
rect 282826 417823 282882 417832
rect 282828 416764 282880 416770
rect 282828 416706 282880 416712
rect 282840 415721 282868 416706
rect 282826 415712 282882 415721
rect 282826 415647 282882 415656
rect 281908 413976 281960 413982
rect 281908 413918 281960 413924
rect 281920 413409 281948 413918
rect 281906 413400 281962 413409
rect 281906 413335 281962 413344
rect 282828 411256 282880 411262
rect 282826 411224 282828 411233
rect 282880 411224 282882 411233
rect 282826 411159 282882 411168
rect 282092 409828 282144 409834
rect 282092 409770 282144 409776
rect 282104 409057 282132 409770
rect 282090 409048 282146 409057
rect 282090 408983 282146 408992
rect 282828 407108 282880 407114
rect 282828 407050 282880 407056
rect 282840 406881 282868 407050
rect 282826 406872 282882 406881
rect 282826 406807 282882 406816
rect 282828 405680 282880 405686
rect 282828 405622 282880 405628
rect 282840 404705 282868 405622
rect 282826 404696 282882 404705
rect 282826 404631 282882 404640
rect 281908 402960 281960 402966
rect 281908 402902 281960 402908
rect 281920 402393 281948 402902
rect 281906 402384 281962 402393
rect 281906 402319 281962 402328
rect 282826 400208 282882 400217
rect 282826 400143 282828 400152
rect 282880 400143 282882 400152
rect 282828 400114 282880 400120
rect 282092 398812 282144 398818
rect 282092 398754 282144 398760
rect 282104 398041 282132 398754
rect 282090 398032 282146 398041
rect 282090 397967 282146 397976
rect 285048 395894 285076 579634
rect 286336 425066 286364 641718
rect 286416 557728 286468 557734
rect 286416 557670 286468 557676
rect 286324 425060 286376 425066
rect 286324 425002 286376 425008
rect 282092 395888 282144 395894
rect 282090 395856 282092 395865
rect 285036 395888 285088 395894
rect 282144 395856 282146 395865
rect 285036 395830 285088 395836
rect 282090 395791 282146 395800
rect 282276 394664 282328 394670
rect 282276 394606 282328 394612
rect 282288 393689 282316 394606
rect 282274 393680 282330 393689
rect 282274 393615 282330 393624
rect 281908 391944 281960 391950
rect 281908 391886 281960 391892
rect 281920 391377 281948 391886
rect 281906 391368 281962 391377
rect 281906 391303 281962 391312
rect 286428 389842 286456 557670
rect 287716 426630 287744 643078
rect 290464 558136 290516 558142
rect 290464 558078 290516 558084
rect 287796 557796 287848 557802
rect 287796 557738 287848 557744
rect 287704 426624 287756 426630
rect 287704 426566 287756 426572
rect 282460 389836 282512 389842
rect 282460 389778 282512 389784
rect 286416 389836 286468 389842
rect 286416 389778 286468 389784
rect 282472 389201 282500 389778
rect 282458 389192 282514 389201
rect 282458 389127 282514 389136
rect 282092 387796 282144 387802
rect 282092 387738 282144 387744
rect 282104 387025 282132 387738
rect 282090 387016 282146 387025
rect 282090 386951 282146 386960
rect 282826 384840 282882 384849
rect 282826 384775 282882 384784
rect 282840 384674 282868 384775
rect 287808 384674 287836 557738
rect 282828 384668 282880 384674
rect 282828 384610 282880 384616
rect 287796 384668 287848 384674
rect 287796 384610 287848 384616
rect 282828 383648 282880 383654
rect 282828 383590 282880 383596
rect 282840 382673 282868 383590
rect 282826 382664 282882 382673
rect 282826 382599 282882 382608
rect 282828 380860 282880 380866
rect 282828 380802 282880 380808
rect 282840 380361 282868 380802
rect 282826 380352 282882 380361
rect 282826 380287 282882 380296
rect 282460 379500 282512 379506
rect 282460 379442 282512 379448
rect 282472 378185 282500 379442
rect 282458 378176 282514 378185
rect 282458 378111 282514 378120
rect 282092 376712 282144 376718
rect 282092 376654 282144 376660
rect 282104 376009 282132 376654
rect 282090 376000 282146 376009
rect 282090 375935 282146 375944
rect 282828 373992 282880 373998
rect 282828 373934 282880 373940
rect 282840 373833 282868 373934
rect 282826 373824 282882 373833
rect 282826 373759 282882 373768
rect 282552 372564 282604 372570
rect 282552 372506 282604 372512
rect 282564 371657 282592 372506
rect 282550 371648 282606 371657
rect 282550 371583 282606 371592
rect 282828 369844 282880 369850
rect 282828 369786 282880 369792
rect 282840 369345 282868 369786
rect 282826 369336 282882 369345
rect 282826 369271 282882 369280
rect 282460 368484 282512 368490
rect 282460 368426 282512 368432
rect 282472 367169 282500 368426
rect 282458 367160 282514 367169
rect 282458 367095 282514 367104
rect 282092 365696 282144 365702
rect 282092 365638 282144 365644
rect 282104 364993 282132 365638
rect 282090 364984 282146 364993
rect 282090 364919 282146 364928
rect 282828 362908 282880 362914
rect 282828 362850 282880 362856
rect 282840 362817 282868 362850
rect 282826 362808 282882 362817
rect 282826 362743 282882 362752
rect 282552 361548 282604 361554
rect 282552 361490 282604 361496
rect 282564 360641 282592 361490
rect 282550 360632 282606 360641
rect 282550 360567 282606 360576
rect 282828 358760 282880 358766
rect 282828 358702 282880 358708
rect 282840 358465 282868 358702
rect 282826 358456 282882 358465
rect 282826 358391 282882 358400
rect 282460 357400 282512 357406
rect 282460 357342 282512 357348
rect 282472 356153 282500 357342
rect 282458 356144 282514 356153
rect 282458 356079 282514 356088
rect 282092 354680 282144 354686
rect 282092 354622 282144 354628
rect 282104 353977 282132 354622
rect 282090 353968 282146 353977
rect 282090 353903 282146 353912
rect 282828 351892 282880 351898
rect 282828 351834 282880 351840
rect 282840 351801 282868 351834
rect 282826 351792 282882 351801
rect 282826 351727 282882 351736
rect 282552 350532 282604 350538
rect 282552 350474 282604 350480
rect 282564 349625 282592 350474
rect 282550 349616 282606 349625
rect 282550 349551 282606 349560
rect 282828 347744 282880 347750
rect 282828 347686 282880 347692
rect 282840 347449 282868 347686
rect 282826 347440 282882 347449
rect 282826 347375 282882 347384
rect 282460 346384 282512 346390
rect 282460 346326 282512 346332
rect 282472 345137 282500 346326
rect 282458 345128 282514 345137
rect 282458 345063 282514 345072
rect 282828 343596 282880 343602
rect 282828 343538 282880 343544
rect 282840 342961 282868 343538
rect 282826 342952 282882 342961
rect 282826 342887 282882 342896
rect 282828 340876 282880 340882
rect 282828 340818 282880 340824
rect 282840 340785 282868 340818
rect 282826 340776 282882 340785
rect 282826 340711 282882 340720
rect 282828 339448 282880 339454
rect 282828 339390 282880 339396
rect 282840 338609 282868 339390
rect 282826 338600 282882 338609
rect 282826 338535 282882 338544
rect 282828 336728 282880 336734
rect 282828 336670 282880 336676
rect 282840 336433 282868 336670
rect 282826 336424 282882 336433
rect 282826 336359 282882 336368
rect 282368 335300 282420 335306
rect 282368 335242 282420 335248
rect 282380 334121 282408 335242
rect 282366 334112 282422 334121
rect 282366 334047 282422 334056
rect 282828 332580 282880 332586
rect 282828 332522 282880 332528
rect 282840 331945 282868 332522
rect 282826 331936 282882 331945
rect 282826 331871 282882 331880
rect 282828 329792 282880 329798
rect 282826 329760 282828 329769
rect 282880 329760 282882 329769
rect 282826 329695 282882 329704
rect 282828 328432 282880 328438
rect 282828 328374 282880 328380
rect 282840 327593 282868 328374
rect 282826 327584 282882 327593
rect 282826 327519 282882 327528
rect 282828 325644 282880 325650
rect 282828 325586 282880 325592
rect 282840 325417 282868 325586
rect 282826 325408 282882 325417
rect 282826 325343 282882 325352
rect 290476 324290 290504 558078
rect 290568 429146 290596 644438
rect 291844 558272 291896 558278
rect 291844 558214 291896 558220
rect 290556 429140 290608 429146
rect 290556 429082 290608 429088
rect 282368 324284 282420 324290
rect 282368 324226 282420 324232
rect 290464 324284 290516 324290
rect 290464 324226 290516 324232
rect 282380 323105 282408 324226
rect 282366 323096 282422 323105
rect 282366 323031 282422 323040
rect 282828 321564 282880 321570
rect 282828 321506 282880 321512
rect 282840 320929 282868 321506
rect 282826 320920 282882 320929
rect 282826 320855 282882 320864
rect 291856 318782 291884 558214
rect 291948 431934 291976 645866
rect 299768 642394 299796 649946
rect 389192 649913 389220 650354
rect 389178 649904 389234 649913
rect 389178 649839 389234 649848
rect 389376 649754 389404 652734
rect 429304 650010 429332 659602
rect 462332 650758 462360 703520
rect 478524 700466 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 494900 692850 494928 703446
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 553306 697368 553362 697377
rect 553490 697368 553546 697377
rect 553362 697326 553490 697354
rect 553306 697303 553362 697312
rect 553490 697303 553546 697312
rect 540978 697232 541034 697241
rect 540978 697167 540980 697176
rect 541032 697167 541034 697176
rect 548616 697196 548668 697202
rect 540980 697138 541032 697144
rect 548616 697138 548668 697144
rect 548628 696969 548656 697138
rect 548614 696960 548670 696969
rect 548614 696895 548670 696904
rect 494060 692844 494112 692850
rect 494060 692786 494112 692792
rect 494888 692844 494940 692850
rect 494888 692786 494940 692792
rect 494072 683074 494100 692786
rect 553306 686352 553362 686361
rect 553490 686352 553546 686361
rect 553362 686310 553490 686338
rect 553306 686287 553362 686296
rect 553490 686287 553546 686296
rect 540978 686216 541034 686225
rect 540978 686151 540980 686160
rect 541032 686151 541034 686160
rect 548616 686180 548668 686186
rect 540980 686122 541032 686128
rect 548616 686122 548668 686128
rect 548628 685953 548656 686122
rect 548614 685944 548670 685953
rect 548614 685879 548670 685888
rect 559668 684554 559696 703520
rect 560298 697368 560354 697377
rect 560298 697303 560300 697312
rect 560352 697303 560354 697312
rect 565176 697332 565228 697338
rect 560300 697274 560352 697280
rect 565176 697274 565228 697280
rect 565188 697241 565216 697274
rect 565174 697232 565230 697241
rect 572718 697232 572774 697241
rect 565174 697167 565230 697176
rect 572640 697190 572718 697218
rect 572640 697105 572668 697190
rect 572718 697167 572774 697176
rect 572626 697096 572682 697105
rect 572626 697031 572682 697040
rect 560298 686352 560354 686361
rect 560298 686287 560300 686296
rect 560352 686287 560354 686296
rect 565176 686316 565228 686322
rect 560300 686258 560352 686264
rect 565176 686258 565228 686264
rect 565188 686225 565216 686258
rect 565174 686216 565230 686225
rect 572718 686216 572774 686225
rect 565174 686151 565230 686160
rect 572640 686174 572718 686202
rect 572640 686089 572668 686174
rect 572718 686151 572774 686160
rect 572626 686080 572682 686089
rect 572626 686015 572682 686024
rect 559012 684548 559064 684554
rect 559012 684490 559064 684496
rect 559656 684548 559708 684554
rect 559656 684490 559708 684496
rect 559024 684457 559052 684490
rect 559010 684448 559066 684457
rect 559010 684383 559066 684392
rect 559010 684312 559066 684321
rect 559010 684247 559066 684256
rect 494072 683046 494284 683074
rect 494256 673538 494284 683046
rect 559024 674898 559052 684247
rect 559012 674892 559064 674898
rect 559012 674834 559064 674840
rect 559380 674892 559432 674898
rect 559380 674834 559432 674840
rect 553398 673976 553454 673985
rect 553398 673911 553454 673920
rect 540978 673840 541034 673849
rect 540978 673775 540980 673784
rect 541032 673775 541034 673784
rect 548616 673804 548668 673810
rect 540980 673746 541032 673752
rect 548616 673746 548668 673752
rect 548628 673577 548656 673746
rect 548614 673568 548670 673577
rect 494060 673532 494112 673538
rect 494060 673474 494112 673480
rect 494244 673532 494296 673538
rect 548614 673503 548670 673512
rect 553306 673568 553362 673577
rect 553412 673554 553440 673911
rect 553362 673526 553440 673554
rect 553306 673503 553362 673512
rect 494244 673474 494296 673480
rect 494072 663762 494100 673474
rect 494072 663734 494284 663762
rect 494256 654158 494284 663734
rect 559392 661774 559420 674834
rect 560298 673976 560354 673985
rect 560298 673911 560300 673920
rect 560352 673911 560354 673920
rect 565176 673940 565228 673946
rect 560300 673882 560352 673888
rect 565176 673882 565228 673888
rect 565188 673849 565216 673882
rect 565174 673840 565230 673849
rect 572718 673840 572774 673849
rect 565174 673775 565230 673784
rect 572640 673798 572718 673826
rect 572640 673713 572668 673798
rect 572718 673775 572774 673784
rect 572626 673704 572682 673713
rect 572626 673639 572682 673648
rect 559104 661768 559156 661774
rect 559104 661710 559156 661716
rect 559380 661768 559432 661774
rect 559380 661710 559432 661716
rect 559116 656946 559144 661710
rect 559104 656940 559156 656946
rect 559104 656882 559156 656888
rect 559196 656940 559248 656946
rect 559196 656882 559248 656888
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 462320 650752 462372 650758
rect 462320 650694 462372 650700
rect 494072 650690 494100 654094
rect 507860 653404 507912 653410
rect 507860 653346 507912 653352
rect 513380 653404 513432 653410
rect 513380 653346 513432 653352
rect 507872 652905 507900 653346
rect 513392 652905 513420 653346
rect 507858 652896 507914 652905
rect 507858 652831 507914 652840
rect 513378 652896 513434 652905
rect 513378 652831 513380 652840
rect 507872 652798 507900 652831
rect 513432 652831 513434 652840
rect 518900 652860 518952 652866
rect 513380 652802 513432 652808
rect 518900 652802 518952 652808
rect 507860 652792 507912 652798
rect 513392 652771 513420 652802
rect 507860 652734 507912 652740
rect 494060 650684 494112 650690
rect 494060 650626 494112 650632
rect 516416 650412 516468 650418
rect 516416 650354 516468 650360
rect 429292 650004 429344 650010
rect 429292 649946 429344 649952
rect 429476 650004 429528 650010
rect 429476 649946 429528 649952
rect 389192 649726 389404 649754
rect 307390 646096 307446 646105
rect 307390 646031 307446 646040
rect 307404 645930 307432 646031
rect 307392 645924 307444 645930
rect 307392 645866 307444 645872
rect 307114 645008 307170 645017
rect 307114 644943 307170 644952
rect 307128 644502 307156 644943
rect 307116 644496 307168 644502
rect 307116 644438 307168 644444
rect 307114 643512 307170 643521
rect 307114 643447 307170 643456
rect 307128 643142 307156 643447
rect 307116 643136 307168 643142
rect 307116 643078 307168 643084
rect 299480 642388 299532 642394
rect 299480 642330 299532 642336
rect 299756 642388 299808 642394
rect 299756 642330 299808 642336
rect 299492 637702 299520 642330
rect 307666 642152 307722 642161
rect 307666 642087 307722 642096
rect 307680 641782 307708 642087
rect 307668 641776 307720 641782
rect 307668 641718 307720 641724
rect 307666 640520 307722 640529
rect 307666 640455 307722 640464
rect 307680 640354 307708 640455
rect 307668 640348 307720 640354
rect 307668 640290 307720 640296
rect 306654 639432 306710 639441
rect 306654 639367 306710 639376
rect 306668 638994 306696 639367
rect 306656 638988 306708 638994
rect 306656 638930 306708 638936
rect 299570 637936 299626 637945
rect 299570 637871 299626 637880
rect 299480 637696 299532 637702
rect 299480 637638 299532 637644
rect 299584 637634 299612 637871
rect 294604 637628 294656 637634
rect 294604 637570 294656 637576
rect 299572 637628 299624 637634
rect 299572 637570 299624 637576
rect 299664 637628 299716 637634
rect 299664 637570 299716 637576
rect 388444 637628 388496 637634
rect 388444 637570 388496 637576
rect 291936 431928 291988 431934
rect 291936 431870 291988 431876
rect 294616 418130 294644 637570
rect 299676 637537 299704 637570
rect 299662 637528 299718 637537
rect 299662 637463 299718 637472
rect 300030 637528 300086 637537
rect 300030 637463 300086 637472
rect 300044 627978 300072 637463
rect 299848 627972 299900 627978
rect 299848 627914 299900 627920
rect 300032 627972 300084 627978
rect 300032 627914 300084 627920
rect 299860 621110 299888 627914
rect 299848 621104 299900 621110
rect 299848 621046 299900 621052
rect 299756 620968 299808 620974
rect 299756 620910 299808 620916
rect 299768 611386 299796 620910
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 299572 608592 299624 608598
rect 299572 608534 299624 608540
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 299584 601730 299612 608534
rect 299572 601724 299624 601730
rect 299572 601666 299624 601672
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299664 598936 299716 598942
rect 299664 598878 299716 598884
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 299676 589354 299704 598878
rect 299664 589348 299716 589354
rect 299664 589290 299716 589296
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 299952 582486 299980 589290
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 306930 580000 306986 580009
rect 306930 579935 306986 579944
rect 306944 579698 306972 579935
rect 306932 579692 306984 579698
rect 306932 579634 306984 579640
rect 306378 578368 306434 578377
rect 306378 578303 306434 578312
rect 306392 578270 306420 578303
rect 306380 578264 306432 578270
rect 299676 572614 299888 572642
rect 306300 578212 306380 578218
rect 306300 578206 306432 578212
rect 306300 578190 306420 578206
rect 299676 563122 299704 572614
rect 299584 563094 299704 563122
rect 299584 562986 299612 563094
rect 299584 562958 299704 562986
rect 299676 553466 299704 562958
rect 306300 560930 306328 578190
rect 306392 578141 306420 578190
rect 306288 560924 306340 560930
rect 306288 560866 306340 560872
rect 347962 559328 348018 559337
rect 347962 559263 348018 559272
rect 357714 559328 357770 559337
rect 357714 559263 357770 559272
rect 313738 558920 313794 558929
rect 313738 558855 313794 558864
rect 316038 558920 316094 558929
rect 316038 558855 316094 558864
rect 318798 558920 318854 558929
rect 318798 558855 318854 558864
rect 320270 558920 320326 558929
rect 320270 558855 320326 558864
rect 321558 558920 321614 558929
rect 321558 558855 321614 558864
rect 323582 558920 323638 558929
rect 323582 558855 323638 558864
rect 325698 558920 325754 558929
rect 325698 558855 325754 558864
rect 327078 558920 327134 558929
rect 327078 558855 327134 558864
rect 329930 558920 329986 558929
rect 329930 558855 329986 558864
rect 331770 558920 331826 558929
rect 331770 558855 331826 558864
rect 332598 558920 332654 558929
rect 332598 558855 332654 558864
rect 333978 558920 334034 558929
rect 333978 558855 334034 558864
rect 335358 558920 335414 558929
rect 336738 558920 336794 558929
rect 335358 558855 335414 558864
rect 335452 558884 335504 558890
rect 313752 558210 313780 558855
rect 313740 558204 313792 558210
rect 313740 558146 313792 558152
rect 302884 557864 302936 557870
rect 302884 557806 302936 557812
rect 299676 553438 299796 553466
rect 299768 539238 299796 553438
rect 299756 539232 299808 539238
rect 299756 539174 299808 539180
rect 294604 418124 294656 418130
rect 294604 418066 294656 418072
rect 282828 318776 282880 318782
rect 282826 318744 282828 318753
rect 291844 318776 291896 318782
rect 282880 318744 282882 318753
rect 291844 318718 291896 318724
rect 282826 318679 282882 318688
rect 282828 317416 282880 317422
rect 282828 317358 282880 317364
rect 282840 316577 282868 317358
rect 282826 316568 282882 316577
rect 282826 316503 282882 316512
rect 282828 314628 282880 314634
rect 282828 314570 282880 314576
rect 282840 314401 282868 314570
rect 282826 314392 282882 314401
rect 282826 314327 282882 314336
rect 282368 313268 282420 313274
rect 282368 313210 282420 313216
rect 282380 312089 282408 313210
rect 282366 312080 282422 312089
rect 282366 312015 282422 312024
rect 281908 310480 281960 310486
rect 281908 310422 281960 310428
rect 281920 309913 281948 310422
rect 281906 309904 281962 309913
rect 281906 309839 281962 309848
rect 302896 307766 302924 557806
rect 316052 416770 316080 558855
rect 317418 558512 317474 558521
rect 317418 558447 317474 558456
rect 317432 557802 317460 558447
rect 317420 557796 317472 557802
rect 317420 557738 317472 557744
rect 316040 416764 316092 416770
rect 316040 416706 316092 416712
rect 318812 387802 318840 558855
rect 320178 557832 320234 557841
rect 320178 557767 320234 557776
rect 320192 557734 320220 557767
rect 320180 557728 320232 557734
rect 320180 557670 320232 557676
rect 320284 391950 320312 558855
rect 320272 391944 320324 391950
rect 320272 391886 320324 391892
rect 318800 387796 318852 387802
rect 318800 387738 318852 387744
rect 282828 307760 282880 307766
rect 282826 307728 282828 307737
rect 302884 307760 302936 307766
rect 282880 307728 282882 307737
rect 302884 307702 302936 307708
rect 282826 307663 282882 307672
rect 321572 306338 321600 558855
rect 322294 558784 322350 558793
rect 322294 558719 322350 558728
rect 322204 558068 322256 558074
rect 322204 558010 322256 558016
rect 322216 317422 322244 558010
rect 322308 557938 322336 558719
rect 322938 557968 322994 557977
rect 322296 557932 322348 557938
rect 322938 557903 322994 557912
rect 322296 557874 322348 557880
rect 322308 451246 322336 557874
rect 322952 557870 322980 557903
rect 322940 557864 322992 557870
rect 322940 557806 322992 557812
rect 322296 451240 322348 451246
rect 322296 451182 322348 451188
rect 322204 317416 322256 317422
rect 322204 317358 322256 317364
rect 323596 310486 323624 558855
rect 323674 558648 323730 558657
rect 323674 558583 323730 558592
rect 324962 558648 325018 558657
rect 324962 558583 325018 558592
rect 323688 557870 323716 558583
rect 323676 557864 323728 557870
rect 323676 557806 323728 557812
rect 323688 454034 323716 557806
rect 324976 557802 325004 558583
rect 324964 557796 325016 557802
rect 324964 557738 325016 557744
rect 324976 455394 325004 557738
rect 324964 455388 325016 455394
rect 324964 455330 325016 455336
rect 323676 454028 323728 454034
rect 323676 453970 323728 453976
rect 325712 313274 325740 558855
rect 326342 558648 326398 558657
rect 326342 558583 326398 558592
rect 326356 557734 326384 558583
rect 326344 557728 326396 557734
rect 326344 557670 326396 557676
rect 326356 458182 326384 557670
rect 326344 458176 326396 458182
rect 326344 458118 326396 458124
rect 327092 314634 327120 558855
rect 327722 558784 327778 558793
rect 327722 558719 327778 558728
rect 329102 558784 329158 558793
rect 329102 558719 329158 558728
rect 327736 558006 327764 558719
rect 328458 558240 328514 558249
rect 328458 558175 328514 558184
rect 328472 558074 328500 558175
rect 329116 558074 329144 558719
rect 329286 558648 329342 558657
rect 329286 558583 329342 558592
rect 328460 558068 328512 558074
rect 328460 558010 328512 558016
rect 329104 558068 329156 558074
rect 329104 558010 329156 558016
rect 327724 558000 327776 558006
rect 327724 557942 327776 557948
rect 327736 460902 327764 557942
rect 329116 462330 329144 558010
rect 329300 557666 329328 558583
rect 329838 558376 329894 558385
rect 329838 558311 329894 558320
rect 329852 558278 329880 558311
rect 329840 558272 329892 558278
rect 329840 558214 329892 558220
rect 329288 557660 329340 557666
rect 329288 557602 329340 557608
rect 329300 465050 329328 557602
rect 329288 465044 329340 465050
rect 329288 464986 329340 464992
rect 329104 462324 329156 462330
rect 329104 462266 329156 462272
rect 327724 460896 327776 460902
rect 327724 460838 327776 460844
rect 329944 321570 329972 558855
rect 330482 558648 330538 558657
rect 330482 558583 330538 558592
rect 330496 557598 330524 558583
rect 331784 558482 331812 558855
rect 331312 558476 331364 558482
rect 331312 558418 331364 558424
rect 331772 558476 331824 558482
rect 331772 558418 331824 558424
rect 331218 558240 331274 558249
rect 331218 558175 331274 558184
rect 331232 558142 331260 558175
rect 331220 558136 331272 558142
rect 331220 558078 331272 558084
rect 331324 557938 331352 558418
rect 331312 557932 331364 557938
rect 331312 557874 331364 557880
rect 330484 557592 330536 557598
rect 330484 557534 330536 557540
rect 330496 466410 330524 557534
rect 330484 466404 330536 466410
rect 330484 466346 330536 466352
rect 332612 325650 332640 558855
rect 332690 558784 332746 558793
rect 332690 558719 332746 558728
rect 332704 558414 332732 558719
rect 332692 558408 332744 558414
rect 332692 558350 332744 558356
rect 332704 557870 332732 558350
rect 332692 557864 332744 557870
rect 332692 557806 332744 557812
rect 333992 328438 334020 558855
rect 334070 558784 334126 558793
rect 334070 558719 334126 558728
rect 334084 558278 334112 558719
rect 334072 558272 334124 558278
rect 334072 558214 334124 558220
rect 334084 557802 334112 558214
rect 334072 557796 334124 557802
rect 334072 557738 334124 557744
rect 335372 329798 335400 558855
rect 336738 558855 336794 558864
rect 337382 558920 337438 558929
rect 337382 558855 337438 558864
rect 338118 558920 338174 558929
rect 338118 558855 338174 558864
rect 339498 558920 339554 558929
rect 339498 558855 339554 558864
rect 340878 558920 340934 558929
rect 340878 558855 340934 558864
rect 342258 558920 342314 558929
rect 342258 558855 342314 558864
rect 343638 558920 343694 558929
rect 343638 558855 343694 558864
rect 344282 558920 344338 558929
rect 344282 558855 344284 558864
rect 335452 558826 335504 558832
rect 335464 558793 335492 558826
rect 335450 558784 335506 558793
rect 335450 558719 335506 558728
rect 336646 558784 336702 558793
rect 336646 558719 336702 558728
rect 335464 557734 335492 558719
rect 336660 558618 336688 558719
rect 336648 558612 336700 558618
rect 336648 558554 336700 558560
rect 336660 558006 336688 558554
rect 336648 558000 336700 558006
rect 336648 557942 336700 557948
rect 335452 557728 335504 557734
rect 335452 557670 335504 557676
rect 336752 332586 336780 558855
rect 337396 558550 337424 558855
rect 337384 558544 337436 558550
rect 336830 558512 336886 558521
rect 337384 558486 337436 558492
rect 336830 558447 336886 558456
rect 336844 335306 336872 558447
rect 337396 558074 337424 558486
rect 337384 558068 337436 558074
rect 337384 558010 337436 558016
rect 338132 336734 338160 558855
rect 338946 558784 339002 558793
rect 338946 558719 339002 558728
rect 338960 558686 338988 558719
rect 338948 558680 339000 558686
rect 338948 558622 339000 558628
rect 338960 557666 338988 558622
rect 338948 557660 339000 557666
rect 338948 557602 339000 557608
rect 339512 339454 339540 558855
rect 339866 558784 339922 558793
rect 339866 558719 339922 558728
rect 339880 558346 339908 558719
rect 339868 558340 339920 558346
rect 339868 558282 339920 558288
rect 339880 557598 339908 558282
rect 339868 557592 339920 557598
rect 339868 557534 339920 557540
rect 340892 340882 340920 558855
rect 340970 558784 341026 558793
rect 340970 558719 341026 558728
rect 340984 558482 341012 558719
rect 340972 558476 341024 558482
rect 340972 558418 341024 558424
rect 342272 343602 342300 558855
rect 342534 558784 342590 558793
rect 342534 558719 342590 558728
rect 342548 558414 342576 558719
rect 342536 558408 342588 558414
rect 342536 558350 342588 558356
rect 343652 346390 343680 558855
rect 344336 558855 344338 558864
rect 345018 558920 345074 558929
rect 345018 558855 345074 558864
rect 346398 558920 346454 558929
rect 346398 558855 346454 558864
rect 347778 558920 347834 558929
rect 347778 558855 347834 558864
rect 344284 558826 344336 558832
rect 343732 558816 343784 558822
rect 343730 558784 343732 558793
rect 343784 558784 343786 558793
rect 344296 558754 344324 558826
rect 343730 558719 343786 558728
rect 344284 558748 344336 558754
rect 343744 558278 343772 558719
rect 344284 558690 344336 558696
rect 343732 558272 343784 558278
rect 343732 558214 343784 558220
rect 343730 557696 343786 557705
rect 343730 557631 343786 557640
rect 343744 347750 343772 557631
rect 345032 350538 345060 558855
rect 346306 558784 346362 558793
rect 346306 558719 346362 558728
rect 346320 558618 346348 558719
rect 346308 558612 346360 558618
rect 346308 558554 346360 558560
rect 346320 558278 346348 558554
rect 346308 558272 346360 558278
rect 346308 558214 346360 558220
rect 346412 351898 346440 558855
rect 346950 558784 347006 558793
rect 346950 558719 347006 558728
rect 346964 558618 346992 558719
rect 346952 558612 347004 558618
rect 346952 558554 347004 558560
rect 347792 354686 347820 558855
rect 347976 558414 348004 559263
rect 349158 558920 349214 558929
rect 349158 558855 349214 558864
rect 351918 558920 351974 558929
rect 351918 558855 351974 558864
rect 355324 558884 355376 558890
rect 348330 558784 348386 558793
rect 348330 558719 348386 558728
rect 348344 558686 348372 558719
rect 348332 558680 348384 558686
rect 348332 558622 348384 558628
rect 347964 558408 348016 558414
rect 347964 558350 348016 558356
rect 349172 357406 349200 558855
rect 351932 558822 351960 558855
rect 355324 558826 355376 558832
rect 351920 558816 351972 558822
rect 349526 558784 349582 558793
rect 351920 558758 351972 558764
rect 353298 558784 353354 558793
rect 349526 558719 349582 558728
rect 353298 558719 353300 558728
rect 349540 558346 349568 558719
rect 353352 558719 353354 558728
rect 353300 558690 353352 558696
rect 350538 558512 350594 558521
rect 350538 558447 350540 558456
rect 350592 558447 350594 558456
rect 350540 558418 350592 558424
rect 354678 558376 354734 558385
rect 349528 558340 349580 558346
rect 354678 558311 354734 558320
rect 349528 558282 349580 558288
rect 354692 558278 354720 558311
rect 354680 558272 354732 558278
rect 354680 558214 354732 558220
rect 349804 558136 349856 558142
rect 349804 558078 349856 558084
rect 349816 471986 349844 558078
rect 352564 558068 352616 558074
rect 352564 558010 352616 558016
rect 352010 557696 352066 557705
rect 352010 557631 352066 557640
rect 350538 557560 350594 557569
rect 350538 557495 350594 557504
rect 349804 471980 349856 471986
rect 349804 471922 349856 471928
rect 350552 358766 350580 557495
rect 352024 362914 352052 557631
rect 352194 555520 352250 555529
rect 352194 555455 352250 555464
rect 352012 362908 352064 362914
rect 352012 362850 352064 362856
rect 352208 361554 352236 555455
rect 352576 514758 352604 558010
rect 352656 558000 352708 558006
rect 352656 557942 352708 557948
rect 352668 517478 352696 557942
rect 352748 557932 352800 557938
rect 352748 557874 352800 557880
rect 352760 520266 352788 557874
rect 353944 557864 353996 557870
rect 353944 557806 353996 557812
rect 353298 557560 353354 557569
rect 353298 557495 353354 557504
rect 352748 520260 352800 520266
rect 352748 520202 352800 520208
rect 352656 517472 352708 517478
rect 352656 517414 352708 517420
rect 352564 514752 352616 514758
rect 352564 514694 352616 514700
rect 353312 365702 353340 557495
rect 353956 521626 353984 557806
rect 354036 557728 354088 557734
rect 354036 557670 354088 557676
rect 354048 524414 354076 557670
rect 354770 557560 354826 557569
rect 354770 557495 354826 557504
rect 354036 524408 354088 524414
rect 354036 524350 354088 524356
rect 353944 521620 353996 521626
rect 353944 521562 353996 521568
rect 354784 368490 354812 557495
rect 355336 525774 355364 558826
rect 357438 558784 357494 558793
rect 357438 558719 357494 558728
rect 357452 558686 357480 558719
rect 357440 558680 357492 558686
rect 356058 558648 356114 558657
rect 357440 558622 357492 558628
rect 356058 558583 356060 558592
rect 356112 558583 356114 558592
rect 356796 558612 356848 558618
rect 356060 558554 356112 558560
rect 356796 558554 356848 558560
rect 356704 557796 356756 557802
rect 356704 557738 356756 557744
rect 356058 557560 356114 557569
rect 356058 557495 356114 557504
rect 355324 525768 355376 525774
rect 355324 525710 355376 525716
rect 356072 369850 356100 557495
rect 356716 528562 356744 557738
rect 356808 531282 356836 558554
rect 357728 558346 357756 559263
rect 358176 558408 358228 558414
rect 358176 558350 358228 558356
rect 357716 558340 357768 558346
rect 357716 558282 357768 558288
rect 358084 557660 358136 557666
rect 358084 557602 358136 557608
rect 357438 557560 357494 557569
rect 357438 557495 357494 557504
rect 356796 531276 356848 531282
rect 356796 531218 356848 531224
rect 356704 528556 356756 528562
rect 356704 528498 356756 528504
rect 357452 372570 357480 557495
rect 358096 473346 358124 557602
rect 358188 476066 358216 558350
rect 359464 558340 359516 558346
rect 359464 558282 359516 558288
rect 358818 555520 358874 555529
rect 358818 555455 358874 555464
rect 358176 476060 358228 476066
rect 358176 476002 358228 476008
rect 358084 473340 358136 473346
rect 358084 473282 358136 473288
rect 358832 373998 358860 555455
rect 359476 477494 359504 558282
rect 359556 558272 359608 558278
rect 359556 558214 359608 558220
rect 359568 480214 359596 558214
rect 359556 480208 359608 480214
rect 359556 480150 359608 480156
rect 359464 477488 359516 477494
rect 359464 477430 359516 477436
rect 388456 400178 388484 637570
rect 389192 589665 389220 649726
rect 399484 645924 399536 645930
rect 399484 645866 399536 645872
rect 398104 644496 398156 644502
rect 398104 644438 398156 644444
rect 395344 643136 395396 643142
rect 395344 643078 395396 643084
rect 393964 641776 394016 641782
rect 393964 641718 394016 641724
rect 392584 640348 392636 640354
rect 392584 640290 392636 640296
rect 391204 638988 391256 638994
rect 391204 638930 391256 638936
rect 389178 589656 389234 589665
rect 389178 589591 389234 589600
rect 391216 402966 391244 638930
rect 392596 405686 392624 640290
rect 393976 407114 394004 641718
rect 395356 409834 395384 643078
rect 398116 411262 398144 644438
rect 399496 413982 399524 645866
rect 429488 642410 429516 649946
rect 516428 649913 516456 650354
rect 516414 649904 516470 649913
rect 516414 649839 516470 649848
rect 437478 646232 437534 646241
rect 437478 646167 437534 646176
rect 437492 645930 437520 646167
rect 437480 645924 437532 645930
rect 437480 645866 437532 645872
rect 437478 644872 437534 644881
rect 437478 644807 437534 644816
rect 437492 644502 437520 644807
rect 437480 644496 437532 644502
rect 437480 644438 437532 644444
rect 437478 643240 437534 643249
rect 437478 643175 437534 643184
rect 437492 643142 437520 643175
rect 437480 643136 437532 643142
rect 437480 643078 437532 643084
rect 429304 642382 429516 642410
rect 429304 637650 429332 642382
rect 437478 642016 437534 642025
rect 437478 641951 437534 641960
rect 437492 641782 437520 641951
rect 437480 641776 437532 641782
rect 437480 641718 437532 641724
rect 437478 640384 437534 640393
rect 437478 640319 437480 640328
rect 437532 640319 437534 640328
rect 437480 640290 437532 640296
rect 437478 639296 437534 639305
rect 437478 639231 437534 639240
rect 437492 638994 437520 639231
rect 437480 638988 437532 638994
rect 437480 638930 437532 638936
rect 437478 637664 437534 637673
rect 429304 637622 429424 637650
rect 429396 637566 429424 637622
rect 437478 637599 437480 637608
rect 437532 637599 437534 637608
rect 437480 637570 437532 637576
rect 429200 637560 429252 637566
rect 429200 637502 429252 637508
rect 429384 637560 429436 637566
rect 429384 637502 429436 637508
rect 429212 627978 429240 637502
rect 429200 627972 429252 627978
rect 429200 627914 429252 627920
rect 429568 627972 429620 627978
rect 429568 627914 429620 627920
rect 429580 621110 429608 627914
rect 429568 621104 429620 621110
rect 429568 621046 429620 621052
rect 429476 620968 429528 620974
rect 429476 620910 429528 620916
rect 429488 611386 429516 620910
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 429396 608598 429424 611238
rect 429292 608592 429344 608598
rect 429292 608534 429344 608540
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 429304 601730 429332 608534
rect 429292 601724 429344 601730
rect 429292 601666 429344 601672
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429384 598936 429436 598942
rect 429384 598878 429436 598884
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 429396 589354 429424 598878
rect 518912 589393 518940 652802
rect 559208 647290 559236 656882
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650350 580212 651063
rect 580172 650344 580224 650350
rect 580172 650286 580224 650292
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 559208 630698 559236 640358
rect 580262 639432 580318 639441
rect 580262 639367 580318 639376
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 559116 621058 559144 630550
rect 559116 621030 559236 621058
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559012 608592 559064 608598
rect 559012 608534 559064 608540
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 559024 601730 559052 608534
rect 559012 601724 559064 601730
rect 559012 601666 559064 601672
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559104 598936 559156 598942
rect 559104 598878 559156 598884
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 518898 589384 518954 589393
rect 429384 589348 429436 589354
rect 429384 589290 429436 589296
rect 429660 589348 429712 589354
rect 559116 589354 559144 598878
rect 518898 589319 518954 589328
rect 559104 589348 559156 589354
rect 429660 589290 429712 589296
rect 429672 582486 429700 589290
rect 518912 587761 518940 589319
rect 559104 589290 559156 589296
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 518898 587752 518954 587761
rect 518898 587687 518954 587696
rect 559392 582486 559420 589290
rect 429660 582480 429712 582486
rect 429660 582422 429712 582428
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 429568 582344 429620 582350
rect 429568 582286 429620 582292
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 402244 579692 402296 579698
rect 402244 579634 402296 579640
rect 399484 413976 399536 413982
rect 399484 413918 399536 413924
rect 398104 411256 398156 411262
rect 398104 411198 398156 411204
rect 395344 409828 395396 409834
rect 395344 409770 395396 409776
rect 393964 407108 394016 407114
rect 393964 407050 394016 407056
rect 392584 405680 392636 405686
rect 392584 405622 392636 405628
rect 391204 402960 391256 402966
rect 391204 402902 391256 402908
rect 388444 400172 388496 400178
rect 388444 400114 388496 400120
rect 402256 394670 402284 579634
rect 429580 572642 429608 582286
rect 437478 579728 437534 579737
rect 437478 579663 437480 579672
rect 437532 579663 437534 579672
rect 437480 579634 437532 579640
rect 438122 578368 438178 578377
rect 438122 578303 438178 578312
rect 429396 572614 429608 572642
rect 429396 563122 429424 572614
rect 429304 563094 429424 563122
rect 429304 562986 429332 563094
rect 429304 562958 429424 562986
rect 429396 553466 429424 562958
rect 438136 560930 438164 578303
rect 559300 572642 559328 582286
rect 559116 572614 559328 572642
rect 438124 560924 438176 560930
rect 438124 560866 438176 560872
rect 559116 560318 559144 572614
rect 559012 560312 559064 560318
rect 559012 560254 559064 560260
rect 559104 560312 559156 560318
rect 559104 560254 559156 560260
rect 443090 558920 443146 558929
rect 443090 558855 443146 558864
rect 445758 558920 445814 558929
rect 445758 558855 445814 558864
rect 446402 558920 446458 558929
rect 446402 558855 446458 558864
rect 447782 558920 447838 558929
rect 447782 558855 447838 558864
rect 449162 558920 449218 558929
rect 449162 558855 449218 558864
rect 452750 558920 452806 558929
rect 452750 558855 452806 558864
rect 453486 558920 453542 558929
rect 453486 558855 453542 558864
rect 454682 558920 454738 558929
rect 454682 558855 454738 558864
rect 458822 558920 458878 558929
rect 458822 558855 458878 558864
rect 460938 558920 460994 558929
rect 460938 558855 460994 558864
rect 461766 558920 461822 558929
rect 461766 558855 461822 558864
rect 462318 558920 462374 558929
rect 462318 558855 462374 558864
rect 463698 558920 463754 558929
rect 463698 558855 463754 558864
rect 465078 558920 465134 558929
rect 465078 558855 465134 558864
rect 466458 558920 466514 558929
rect 466458 558855 466514 558864
rect 467838 558920 467894 558929
rect 467838 558855 467894 558864
rect 468574 558920 468630 558929
rect 468574 558855 468630 558864
rect 469218 558920 469274 558929
rect 469218 558855 469274 558864
rect 470598 558920 470654 558929
rect 470598 558855 470654 558864
rect 471978 558920 472034 558929
rect 471978 558855 472034 558864
rect 473358 558920 473414 558929
rect 473358 558855 473414 558864
rect 474738 558920 474794 558929
rect 474738 558855 474794 558864
rect 476210 558920 476266 558929
rect 476210 558855 476266 558864
rect 477130 558920 477186 558929
rect 477130 558855 477186 558864
rect 478326 558920 478382 558929
rect 478326 558855 478382 558864
rect 479430 558920 479486 558929
rect 479430 558855 479486 558864
rect 480534 558920 480590 558929
rect 480534 558855 480590 558864
rect 483018 558920 483074 558929
rect 483018 558855 483020 558864
rect 443104 558210 443132 558855
rect 443092 558204 443144 558210
rect 443092 558146 443144 558152
rect 443644 558204 443696 558210
rect 443644 558146 443696 558152
rect 429396 553438 429516 553466
rect 429488 539170 429516 553438
rect 429476 539164 429528 539170
rect 429476 539106 429528 539112
rect 443656 483002 443684 558146
rect 443644 482996 443696 483002
rect 443644 482938 443696 482944
rect 445772 398818 445800 558855
rect 445760 398812 445812 398818
rect 445760 398754 445812 398760
rect 402244 394664 402296 394670
rect 402244 394606 402296 394612
rect 446416 376718 446444 558855
rect 447796 379506 447824 558855
rect 449176 380866 449204 558855
rect 452658 558240 452714 558249
rect 452658 558175 452714 558184
rect 452672 558142 452700 558175
rect 452660 558136 452712 558142
rect 452660 558078 452712 558084
rect 451370 557696 451426 557705
rect 451370 557631 451426 557640
rect 451384 557598 451412 557631
rect 450544 557592 450596 557598
rect 450544 557534 450596 557540
rect 451372 557592 451424 557598
rect 451372 557534 451424 557540
rect 450556 383654 450584 557534
rect 452764 469198 452792 558855
rect 453302 558784 453358 558793
rect 453302 558719 453358 558728
rect 453316 558482 453344 558719
rect 453500 558618 453528 558855
rect 453488 558612 453540 558618
rect 453488 558554 453540 558560
rect 453304 558476 453356 558482
rect 453304 558418 453356 558424
rect 452752 469192 452804 469198
rect 452752 469134 452804 469140
rect 453316 433294 453344 558418
rect 453500 436082 453528 558554
rect 454038 558376 454094 558385
rect 454038 558311 454094 558320
rect 454052 557666 454080 558311
rect 454696 558142 454724 558855
rect 458836 558822 458864 558855
rect 458824 558816 458876 558822
rect 458824 558758 458876 558764
rect 460202 558784 460258 558793
rect 456062 558648 456118 558657
rect 456062 558583 456118 558592
rect 457442 558648 457498 558657
rect 457442 558583 457498 558592
rect 455418 558512 455474 558521
rect 455418 558447 455474 558456
rect 455432 558414 455460 558447
rect 455420 558408 455472 558414
rect 455420 558350 455472 558356
rect 454684 558136 454736 558142
rect 454684 558078 454736 558084
rect 454040 557660 454092 557666
rect 454040 557602 454092 557608
rect 454696 438870 454724 558078
rect 456076 557666 456104 558583
rect 456798 558376 456854 558385
rect 456798 558311 456800 558320
rect 456852 558311 456854 558320
rect 456800 558282 456852 558288
rect 456064 557660 456116 557666
rect 456064 557602 456116 557608
rect 456076 440230 456104 557602
rect 457456 557598 457484 558583
rect 458178 558376 458234 558385
rect 458178 558311 458234 558320
rect 458192 558278 458220 558311
rect 458180 558272 458232 558278
rect 458180 558214 458232 558220
rect 457444 557592 457496 557598
rect 457444 557534 457496 557540
rect 457456 442950 457484 557534
rect 458836 444378 458864 558758
rect 460202 558719 460258 558728
rect 460662 558784 460718 558793
rect 460662 558719 460664 558728
rect 459558 558240 459614 558249
rect 459558 558175 459560 558184
rect 459612 558175 459614 558184
rect 459560 558146 459612 558152
rect 460216 447098 460244 558719
rect 460716 558719 460718 558728
rect 460664 558690 460716 558696
rect 460846 558648 460902 558657
rect 460846 558583 460902 558592
rect 460860 558550 460888 558583
rect 460388 558544 460440 558550
rect 460388 558486 460440 558492
rect 460848 558544 460900 558550
rect 460848 558486 460900 558492
rect 460400 449886 460428 558486
rect 460952 484362 460980 558855
rect 461030 558784 461086 558793
rect 461030 558719 461086 558728
rect 461044 487150 461072 558719
rect 461780 558482 461808 558855
rect 461768 558476 461820 558482
rect 461768 558418 461820 558424
rect 462332 488510 462360 558855
rect 462962 558784 463018 558793
rect 462962 558719 463018 558728
rect 462976 558618 463004 558719
rect 462964 558612 463016 558618
rect 462964 558554 463016 558560
rect 463608 558612 463660 558618
rect 463608 558554 463660 558560
rect 463620 558414 463648 558554
rect 463608 558408 463660 558414
rect 463608 558350 463660 558356
rect 463712 491298 463740 558855
rect 464342 558784 464398 558793
rect 464342 558719 464398 558728
rect 464356 558618 464384 558719
rect 464344 558612 464396 558618
rect 464344 558554 464396 558560
rect 464356 558226 464384 558554
rect 464264 558198 464384 558226
rect 464264 558142 464292 558198
rect 464252 558136 464304 558142
rect 464252 558078 464304 558084
rect 464344 558136 464396 558142
rect 464344 558078 464396 558084
rect 464356 532710 464384 558078
rect 464344 532704 464396 532710
rect 464344 532646 464396 532652
rect 465092 494018 465120 558855
rect 465170 558784 465226 558793
rect 465170 558719 465226 558728
rect 465184 558346 465212 558719
rect 465172 558340 465224 558346
rect 465172 558282 465224 558288
rect 465184 557666 465212 558282
rect 465724 558204 465776 558210
rect 465724 558146 465776 558152
rect 465172 557660 465224 557666
rect 465172 557602 465224 557608
rect 465736 535430 465764 558146
rect 465724 535424 465776 535430
rect 465724 535366 465776 535372
rect 466472 495446 466500 558855
rect 466550 558648 466606 558657
rect 466550 558583 466606 558592
rect 466564 557598 466592 558583
rect 467104 558272 467156 558278
rect 467104 558214 467156 558220
rect 466552 557592 466604 557598
rect 466552 557534 466604 557540
rect 467116 536790 467144 558214
rect 467104 536784 467156 536790
rect 467104 536726 467156 536732
rect 467852 498166 467880 558855
rect 468024 558816 468076 558822
rect 467930 558784 467986 558793
rect 468024 558758 468076 558764
rect 467930 558719 467986 558728
rect 467944 499526 467972 558719
rect 468036 558657 468064 558758
rect 468588 558754 468616 558855
rect 468576 558748 468628 558754
rect 468576 558690 468628 558696
rect 468022 558648 468078 558657
rect 468022 558583 468078 558592
rect 468588 557666 468616 558690
rect 468576 557660 468628 557666
rect 468576 557602 468628 557608
rect 469232 502314 469260 558855
rect 470046 558784 470102 558793
rect 470046 558719 470102 558728
rect 470060 558550 470088 558719
rect 470048 558544 470100 558550
rect 470048 558486 470100 558492
rect 470612 503674 470640 558855
rect 471242 558784 471298 558793
rect 471242 558719 471298 558728
rect 471256 558482 471284 558719
rect 471244 558476 471296 558482
rect 471244 558418 471296 558424
rect 471992 506462 472020 558855
rect 472254 558784 472310 558793
rect 472254 558719 472310 558728
rect 472268 558414 472296 558719
rect 472256 558408 472308 558414
rect 472256 558350 472308 558356
rect 473372 509250 473400 558855
rect 473542 558784 473598 558793
rect 473542 558719 473598 558728
rect 473556 558618 473584 558719
rect 473544 558612 473596 558618
rect 473544 558554 473596 558560
rect 474646 557696 474702 557705
rect 474646 557631 474702 557640
rect 474660 557598 474688 557631
rect 474648 557592 474700 557598
rect 474648 557534 474700 557540
rect 474752 510610 474780 558855
rect 474830 558784 474886 558793
rect 474830 558719 474886 558728
rect 475566 558784 475622 558793
rect 475566 558719 475568 558728
rect 474844 558346 474872 558719
rect 475620 558719 475622 558728
rect 475568 558690 475620 558696
rect 474832 558340 474884 558346
rect 474832 558282 474884 558288
rect 474844 557598 474872 558282
rect 476118 558104 476174 558113
rect 476118 558039 476120 558048
rect 476172 558039 476174 558048
rect 476120 558010 476172 558016
rect 474832 557592 474884 557598
rect 474832 557534 474884 557540
rect 476224 513330 476252 558855
rect 477144 558822 477172 558855
rect 477132 558816 477184 558822
rect 477132 558758 477184 558764
rect 478340 558346 478368 558855
rect 479444 558550 479472 558855
rect 480442 558784 480498 558793
rect 480442 558719 480498 558728
rect 479432 558544 479484 558550
rect 479432 558486 479484 558492
rect 480456 558482 480484 558719
rect 480444 558476 480496 558482
rect 480444 558418 480496 558424
rect 477592 558340 477644 558346
rect 477592 558282 477644 558288
rect 478328 558340 478380 558346
rect 478328 558282 478380 558288
rect 477498 558104 477554 558113
rect 477498 558039 477554 558048
rect 477512 558006 477540 558039
rect 477500 558000 477552 558006
rect 477500 557942 477552 557948
rect 477604 557666 477632 558282
rect 478878 557968 478934 557977
rect 478878 557903 478880 557912
rect 478932 557903 478934 557912
rect 478880 557874 478932 557880
rect 480548 557870 480576 558855
rect 483072 558855 483074 558864
rect 484490 558920 484546 558929
rect 484490 558855 484546 558864
rect 485778 558920 485834 558929
rect 485778 558855 485834 558864
rect 483020 558826 483072 558832
rect 484398 558784 484454 558793
rect 484398 558719 484400 558728
rect 484452 558719 484454 558728
rect 484400 558690 484452 558696
rect 484504 558686 484532 558855
rect 485792 558822 485820 558855
rect 485780 558816 485832 558822
rect 485780 558758 485832 558764
rect 484492 558680 484544 558686
rect 483018 558648 483074 558657
rect 484492 558622 484544 558628
rect 488538 558648 488594 558657
rect 483018 558583 483020 558592
rect 483072 558583 483074 558592
rect 488538 558583 488594 558592
rect 483020 558554 483072 558560
rect 488552 558550 488580 558583
rect 488540 558544 488592 558550
rect 481638 558512 481694 558521
rect 481638 558447 481694 558456
rect 487158 558512 487214 558521
rect 488540 558486 488592 558492
rect 487158 558447 487214 558456
rect 481652 558414 481680 558447
rect 481640 558408 481692 558414
rect 481640 558350 481692 558356
rect 487172 558346 487200 558447
rect 488538 558376 488594 558385
rect 487160 558340 487212 558346
rect 488538 558311 488594 558320
rect 487160 558282 487212 558288
rect 488552 558278 488580 558311
rect 488540 558272 488592 558278
rect 483018 558240 483074 558249
rect 483018 558175 483074 558184
rect 485778 558240 485834 558249
rect 485778 558175 485834 558184
rect 487158 558240 487214 558249
rect 488540 558214 488592 558220
rect 487158 558175 487160 558184
rect 480536 557864 480588 557870
rect 480536 557806 480588 557812
rect 481638 557832 481694 557841
rect 483032 557802 483060 558175
rect 485792 558142 485820 558175
rect 487212 558175 487214 558184
rect 487160 558146 487212 558152
rect 485780 558136 485832 558142
rect 485780 558078 485832 558084
rect 481638 557767 481694 557776
rect 483020 557796 483072 557802
rect 481652 557734 481680 557767
rect 483020 557738 483072 557744
rect 481640 557728 481692 557734
rect 481640 557670 481692 557676
rect 483018 557696 483074 557705
rect 477592 557660 477644 557666
rect 483018 557631 483074 557640
rect 477592 557602 477644 557608
rect 483032 557598 483060 557631
rect 483020 557592 483072 557598
rect 483020 557534 483072 557540
rect 559024 553330 559052 560254
rect 579618 557288 579674 557297
rect 579618 557223 579674 557232
rect 579632 556238 579660 557223
rect 579620 556232 579672 556238
rect 579620 556174 579672 556180
rect 559024 553302 559144 553330
rect 559116 543810 559144 553302
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 559116 543782 559236 543810
rect 559208 539102 559236 543782
rect 580276 539209 580304 639367
rect 580354 627736 580410 627745
rect 580354 627671 580410 627680
rect 580262 539200 580318 539209
rect 580262 539135 580318 539144
rect 559196 539096 559248 539102
rect 559196 539038 559248 539044
rect 580368 539034 580396 627671
rect 580446 604208 580502 604217
rect 580446 604143 580502 604152
rect 580460 539073 580488 604143
rect 580538 592512 580594 592521
rect 580538 592447 580594 592456
rect 580446 539064 580502 539073
rect 580356 539028 580408 539034
rect 580446 538999 580502 539008
rect 580356 538970 580408 538976
rect 580552 538898 580580 592447
rect 580630 580816 580686 580825
rect 580630 580751 580686 580760
rect 580644 538966 580672 580751
rect 580632 538960 580684 538966
rect 580632 538902 580684 538908
rect 580540 538892 580592 538898
rect 580540 538834 580592 538840
rect 541624 538416 541676 538422
rect 541624 538358 541676 538364
rect 541636 530602 541664 538358
rect 563704 538348 563756 538354
rect 563704 538290 563756 538296
rect 541624 530596 541676 530602
rect 541624 530538 541676 530544
rect 556160 530596 556212 530602
rect 556160 530538 556212 530544
rect 556172 529242 556200 530538
rect 563716 530058 563744 538290
rect 579804 538280 579856 538286
rect 579804 538222 579856 538228
rect 579816 533905 579844 538222
rect 580264 537940 580316 537946
rect 580264 537882 580316 537888
rect 579802 533896 579858 533905
rect 579802 533831 579858 533840
rect 563704 530052 563756 530058
rect 563704 529994 563756 530000
rect 569224 529916 569276 529922
rect 569224 529858 569276 529864
rect 556160 529236 556212 529242
rect 556160 529178 556212 529184
rect 568488 529236 568540 529242
rect 568488 529178 568540 529184
rect 568500 525842 568528 529178
rect 568488 525836 568540 525842
rect 568488 525778 568540 525784
rect 569236 521626 569264 529858
rect 571984 525768 572036 525774
rect 571984 525710 572036 525716
rect 569224 521620 569276 521626
rect 569224 521562 569276 521568
rect 570972 521620 571024 521626
rect 570972 521562 571024 521568
rect 570984 517546 571012 521562
rect 570972 517540 571024 517546
rect 570972 517482 571024 517488
rect 571996 513330 572024 525710
rect 573364 517472 573416 517478
rect 573364 517414 573416 517420
rect 476212 513324 476264 513330
rect 476212 513266 476264 513272
rect 571984 513324 572036 513330
rect 571984 513266 572036 513272
rect 474740 510604 474792 510610
rect 474740 510546 474792 510552
rect 473360 509244 473412 509250
rect 473360 509186 473412 509192
rect 471980 506456 472032 506462
rect 471980 506398 472032 506404
rect 470600 503668 470652 503674
rect 470600 503610 470652 503616
rect 469220 502308 469272 502314
rect 469220 502250 469272 502256
rect 573376 499594 573404 517414
rect 574744 513324 574796 513330
rect 574744 513266 574796 513272
rect 574756 507822 574784 513266
rect 580276 510377 580304 537882
rect 580262 510368 580318 510377
rect 580262 510303 580318 510312
rect 574744 507816 574796 507822
rect 574744 507758 574796 507764
rect 577964 507816 578016 507822
rect 577964 507758 578016 507764
rect 577976 506326 578004 507758
rect 577964 506320 578016 506326
rect 577964 506262 578016 506268
rect 580264 506320 580316 506326
rect 580264 506262 580316 506268
rect 573364 499588 573416 499594
rect 573364 499530 573416 499536
rect 467932 499520 467984 499526
rect 467932 499462 467984 499468
rect 576768 499520 576820 499526
rect 576768 499462 576820 499468
rect 467840 498160 467892 498166
rect 467840 498102 467892 498108
rect 576780 496754 576808 499462
rect 580276 498681 580304 506262
rect 580262 498672 580318 498681
rect 580262 498607 580318 498616
rect 576780 496726 576900 496754
rect 466460 495440 466512 495446
rect 466460 495382 466512 495388
rect 465080 494012 465132 494018
rect 465080 493954 465132 493960
rect 576872 493882 576900 496726
rect 576860 493876 576912 493882
rect 576860 493818 576912 493824
rect 578884 493876 578936 493882
rect 578884 493818 578936 493824
rect 463700 491292 463752 491298
rect 463700 491234 463752 491240
rect 462320 488504 462372 488510
rect 462320 488446 462372 488452
rect 461032 487144 461084 487150
rect 461032 487086 461084 487092
rect 578896 486849 578924 493818
rect 578882 486840 578938 486849
rect 578882 486775 578938 486784
rect 460940 484356 460992 484362
rect 460940 484298 460992 484304
rect 579986 463448 580042 463457
rect 579986 463383 580042 463392
rect 580000 462058 580028 463383
rect 576860 462052 576912 462058
rect 576860 461994 576912 462000
rect 579988 462052 580040 462058
rect 579988 461994 580040 462000
rect 576872 459610 576900 461994
rect 571800 459604 571852 459610
rect 571800 459546 571852 459552
rect 576860 459604 576912 459610
rect 576860 459546 576912 459552
rect 571812 456074 571840 459546
rect 566464 456068 566516 456074
rect 566464 456010 566516 456016
rect 571800 456068 571852 456074
rect 571800 456010 571852 456016
rect 460388 449880 460440 449886
rect 460388 449822 460440 449828
rect 460204 447092 460256 447098
rect 460204 447034 460256 447040
rect 566476 445806 566504 456010
rect 580262 451752 580318 451761
rect 580262 451687 580318 451696
rect 566464 445800 566516 445806
rect 566464 445742 566516 445748
rect 563244 445732 563296 445738
rect 563244 445674 563296 445680
rect 458824 444372 458876 444378
rect 458824 444314 458876 444320
rect 457444 442944 457496 442950
rect 457444 442886 457496 442892
rect 563256 442202 563284 445674
rect 562416 442196 562468 442202
rect 562416 442138 562468 442144
rect 563244 442196 563296 442202
rect 563244 442138 563296 442144
rect 456064 440224 456116 440230
rect 456064 440166 456116 440172
rect 562428 438938 562456 442138
rect 580276 440298 580304 451687
rect 578608 440292 578660 440298
rect 578608 440234 578660 440240
rect 580264 440292 580316 440298
rect 580264 440234 580316 440240
rect 578620 438938 578648 440234
rect 579618 439920 579674 439929
rect 579618 439855 579674 439864
rect 560944 438932 560996 438938
rect 560944 438874 560996 438880
rect 562416 438932 562468 438938
rect 562416 438874 562468 438880
rect 576124 438932 576176 438938
rect 576124 438874 576176 438880
rect 578608 438932 578660 438938
rect 578608 438874 578660 438880
rect 454684 438864 454736 438870
rect 454684 438806 454736 438812
rect 453488 436076 453540 436082
rect 453488 436018 453540 436024
rect 453304 433288 453356 433294
rect 453304 433230 453356 433236
rect 560956 418198 560984 438874
rect 575848 435532 575900 435538
rect 575848 435474 575900 435480
rect 575860 432546 575888 435474
rect 574744 432540 574796 432546
rect 574744 432482 574796 432488
rect 575848 432540 575900 432546
rect 575848 432482 575900 432488
rect 570604 426828 570656 426834
rect 570604 426770 570656 426776
rect 567844 419552 567896 419558
rect 567844 419494 567896 419500
rect 558184 418192 558236 418198
rect 558184 418134 558236 418140
rect 560944 418192 560996 418198
rect 560944 418134 560996 418140
rect 558196 399702 558224 418134
rect 556804 399696 556856 399702
rect 556804 399638 556856 399644
rect 558184 399696 558236 399702
rect 558184 399638 558236 399644
rect 556816 387802 556844 399638
rect 567856 392018 567884 419494
rect 570616 394670 570644 426770
rect 574756 422754 574784 432482
rect 576136 426834 576164 438874
rect 579632 437646 579660 439855
rect 577964 437640 578016 437646
rect 577964 437582 578016 437588
rect 579620 437640 579672 437646
rect 579620 437582 579672 437588
rect 577976 435538 578004 437582
rect 577964 435532 578016 435538
rect 577964 435474 578016 435480
rect 576124 426828 576176 426834
rect 576124 426770 576176 426776
rect 570788 422748 570840 422754
rect 570788 422690 570840 422696
rect 574744 422748 574796 422754
rect 574744 422690 574796 422696
rect 570800 419558 570828 422690
rect 570788 419552 570840 419558
rect 570788 419494 570840 419500
rect 580262 416528 580318 416537
rect 580262 416463 580318 416472
rect 580276 405754 580304 416463
rect 578976 405748 579028 405754
rect 578976 405690 579028 405696
rect 580264 405748 580316 405754
rect 580264 405690 580316 405696
rect 578988 403578 579016 405690
rect 580906 404832 580962 404841
rect 580906 404767 580962 404776
rect 577596 403572 577648 403578
rect 577596 403514 577648 403520
rect 578976 403572 579028 403578
rect 578976 403514 579028 403520
rect 577504 400240 577556 400246
rect 577504 400182 577556 400188
rect 569224 394664 569276 394670
rect 569224 394606 569276 394612
rect 570604 394664 570656 394670
rect 570604 394606 570656 394612
rect 566556 392012 566608 392018
rect 566556 391954 566608 391960
rect 567844 392012 567896 392018
rect 567844 391954 567896 391960
rect 555424 387796 555476 387802
rect 555424 387738 555476 387744
rect 556804 387796 556856 387802
rect 556804 387738 556856 387744
rect 450544 383648 450596 383654
rect 450544 383590 450596 383596
rect 449164 380860 449216 380866
rect 449164 380802 449216 380808
rect 447784 379500 447836 379506
rect 447784 379442 447836 379448
rect 446404 376712 446456 376718
rect 446404 376654 446456 376660
rect 358820 373992 358872 373998
rect 358820 373934 358872 373940
rect 357440 372564 357492 372570
rect 357440 372506 357492 372512
rect 356060 369844 356112 369850
rect 356060 369786 356112 369792
rect 354772 368484 354824 368490
rect 354772 368426 354824 368432
rect 353300 365696 353352 365702
rect 353300 365638 353352 365644
rect 352196 361548 352248 361554
rect 352196 361490 352248 361496
rect 553308 360868 553360 360874
rect 553308 360810 553360 360816
rect 350540 358760 350592 358766
rect 350540 358702 350592 358708
rect 349160 357400 349212 357406
rect 349160 357342 349212 357348
rect 553320 356658 553348 360810
rect 551284 356652 551336 356658
rect 551284 356594 551336 356600
rect 553308 356652 553360 356658
rect 553308 356594 553360 356600
rect 347780 354680 347832 354686
rect 347780 354622 347832 354628
rect 551296 351966 551324 356594
rect 555436 351966 555464 387738
rect 566464 371748 566516 371754
rect 566464 371690 566516 371696
rect 565268 369912 565320 369918
rect 565268 369854 565320 369860
rect 564072 369844 564124 369850
rect 564072 369786 564124 369792
rect 563704 368484 563756 368490
rect 563704 368426 563756 368432
rect 560944 367124 560996 367130
rect 560944 367066 560996 367072
rect 549260 351960 549312 351966
rect 549260 351902 549312 351908
rect 551284 351960 551336 351966
rect 551284 351902 551336 351908
rect 554044 351960 554096 351966
rect 554044 351902 554096 351908
rect 555424 351960 555476 351966
rect 555424 351902 555476 351908
rect 346400 351892 346452 351898
rect 346400 351834 346452 351840
rect 345020 350532 345072 350538
rect 345020 350474 345072 350480
rect 343732 347744 343784 347750
rect 343732 347686 343784 347692
rect 343640 346384 343692 346390
rect 343640 346326 343692 346332
rect 549272 345914 549300 351902
rect 548524 345908 548576 345914
rect 548524 345850 548576 345856
rect 549260 345908 549312 345914
rect 549260 345850 549312 345856
rect 342260 343596 342312 343602
rect 342260 343538 342312 343544
rect 340880 340876 340932 340882
rect 340880 340818 340932 340824
rect 339500 339448 339552 339454
rect 339500 339390 339552 339396
rect 338120 336728 338172 336734
rect 338120 336670 338172 336676
rect 336832 335300 336884 335306
rect 336832 335242 336884 335248
rect 336740 332580 336792 332586
rect 336740 332522 336792 332528
rect 548536 331226 548564 345850
rect 554056 342310 554084 351902
rect 560956 348430 560984 367066
rect 563716 357066 563744 368426
rect 563796 368076 563848 368082
rect 563796 368018 563848 368024
rect 563808 360874 563836 368018
rect 564084 367130 564112 369786
rect 565280 368082 565308 369854
rect 565268 368076 565320 368082
rect 565268 368018 565320 368024
rect 564072 367124 564124 367130
rect 564072 367066 564124 367072
rect 563796 360868 563848 360874
rect 563796 360810 563848 360816
rect 562416 357060 562468 357066
rect 562416 357002 562468 357008
rect 563704 357060 563756 357066
rect 563704 357002 563756 357008
rect 562428 350606 562456 357002
rect 561036 350600 561088 350606
rect 561036 350542 561088 350548
rect 562416 350600 562468 350606
rect 562416 350542 562468 350548
rect 559564 348424 559616 348430
rect 559564 348366 559616 348372
rect 560944 348424 560996 348430
rect 560944 348366 560996 348372
rect 558460 343596 558512 343602
rect 558460 343538 558512 343544
rect 552664 342304 552716 342310
rect 552664 342246 552716 342252
rect 554044 342304 554096 342310
rect 554044 342246 554096 342252
rect 551376 338156 551428 338162
rect 551376 338098 551428 338104
rect 551284 334008 551336 334014
rect 551284 333950 551336 333956
rect 546500 331220 546552 331226
rect 546500 331162 546552 331168
rect 548524 331220 548576 331226
rect 548524 331162 548576 331168
rect 335360 329792 335412 329798
rect 335360 329734 335412 329740
rect 333980 328432 334032 328438
rect 333980 328374 334032 328380
rect 546512 325718 546540 331162
rect 549352 328160 549404 328166
rect 549352 328102 549404 328108
rect 549260 327752 549312 327758
rect 549260 327694 549312 327700
rect 546500 325712 546552 325718
rect 546500 325654 546552 325660
rect 332600 325644 332652 325650
rect 332600 325586 332652 325592
rect 543740 325644 543792 325650
rect 543740 325586 543792 325592
rect 543752 323610 543780 325586
rect 545120 324352 545172 324358
rect 545120 324294 545172 324300
rect 535460 323604 535512 323610
rect 535460 323546 535512 323552
rect 543740 323604 543792 323610
rect 543740 323546 543792 323552
rect 535472 321638 535500 323546
rect 532884 321632 532936 321638
rect 532884 321574 532936 321580
rect 535460 321632 535512 321638
rect 535460 321574 535512 321580
rect 329932 321564 329984 321570
rect 329932 321506 329984 321512
rect 532896 319258 532924 321574
rect 544108 321496 544160 321502
rect 544108 321438 544160 321444
rect 543004 320204 543056 320210
rect 543004 320146 543056 320152
rect 529572 319252 529624 319258
rect 529572 319194 529624 319200
rect 532884 319252 532936 319258
rect 532884 319194 532936 319200
rect 529584 316062 529612 319194
rect 542084 317008 542136 317014
rect 542084 316950 542136 316956
rect 529572 316056 529624 316062
rect 529572 315998 529624 316004
rect 523500 315988 523552 315994
rect 523500 315930 523552 315936
rect 327080 314628 327132 314634
rect 327080 314570 327132 314576
rect 325700 313268 325752 313274
rect 325700 313210 325752 313216
rect 323584 310480 323636 310486
rect 323584 310422 323636 310428
rect 519544 309800 519596 309806
rect 519544 309742 519596 309748
rect 282092 306332 282144 306338
rect 282092 306274 282144 306280
rect 321560 306332 321612 306338
rect 321560 306274 321612 306280
rect 282104 305561 282132 306274
rect 517520 305652 517572 305658
rect 517520 305594 517572 305600
rect 282090 305552 282146 305561
rect 282090 305487 282146 305496
rect 516140 305040 516192 305046
rect 516140 304982 516192 304988
rect 281630 301200 281686 301209
rect 281630 301135 281686 301144
rect 514760 300892 514812 300898
rect 514760 300834 514812 300840
rect 60844 300750 60950 300778
rect 60844 300665 60872 300750
rect 60830 300656 60886 300665
rect 60830 300591 60886 300600
rect 60648 300552 60700 300558
rect 60648 300494 60700 300500
rect 59544 300348 59596 300354
rect 59544 300290 59596 300296
rect 514772 300150 514800 300834
rect 516152 300218 516180 304982
rect 517532 300898 517560 305594
rect 519556 305046 519584 309742
rect 523512 307154 523540 315930
rect 542096 311982 542124 316950
rect 539968 311976 540020 311982
rect 539968 311918 540020 311924
rect 542084 311976 542136 311982
rect 542084 311918 542136 311924
rect 535460 311160 535512 311166
rect 535460 311102 535512 311108
rect 535472 309194 535500 311102
rect 539980 309806 540008 311918
rect 543016 311166 543044 320146
rect 544120 317014 544148 321438
rect 545132 320210 545160 324294
rect 549168 322992 549220 322998
rect 549168 322934 549220 322940
rect 548524 320748 548576 320754
rect 548524 320690 548576 320696
rect 545120 320204 545172 320210
rect 545120 320146 545172 320152
rect 546500 319796 546552 319802
rect 546500 319738 546552 319744
rect 544108 317008 544160 317014
rect 544108 316950 544160 316956
rect 546512 316674 546540 319738
rect 545212 316668 545264 316674
rect 545212 316610 545264 316616
rect 546500 316668 546552 316674
rect 546500 316610 546552 316616
rect 545224 311914 545252 316610
rect 545212 311908 545264 311914
rect 545212 311850 545264 311856
rect 543096 311840 543148 311846
rect 543096 311782 543148 311788
rect 543004 311160 543056 311166
rect 543004 311102 543056 311108
rect 539968 309800 540020 309806
rect 539968 309742 540020 309748
rect 535460 309188 535512 309194
rect 535460 309130 535512 309136
rect 532332 309120 532384 309126
rect 532332 309062 532384 309068
rect 522488 307148 522540 307154
rect 522488 307090 522540 307096
rect 523500 307148 523552 307154
rect 523500 307090 523552 307096
rect 522500 305658 522528 307090
rect 522488 305652 522540 305658
rect 522488 305594 522540 305600
rect 519544 305040 519596 305046
rect 519544 304982 519596 304988
rect 517520 300892 517572 300898
rect 517520 300834 517572 300840
rect 532344 300286 532372 309062
rect 539692 308712 539744 308718
rect 539692 308654 539744 308660
rect 539704 301034 539732 308654
rect 543108 305046 543136 311782
rect 545120 311024 545172 311030
rect 545120 310966 545172 310972
rect 545132 308718 545160 310966
rect 545120 308712 545172 308718
rect 545120 308654 545172 308660
rect 548536 305046 548564 320690
rect 549180 319802 549208 322934
rect 549272 321638 549300 327694
rect 549364 324358 549392 328102
rect 549352 324352 549404 324358
rect 549352 324294 549404 324300
rect 549260 321632 549312 321638
rect 549260 321574 549312 321580
rect 551296 320754 551324 333950
rect 551388 328166 551416 338098
rect 552676 334014 552704 342246
rect 558472 340950 558500 343538
rect 553400 340944 553452 340950
rect 553400 340886 553452 340892
rect 558460 340944 558512 340950
rect 558460 340886 558512 340892
rect 553412 338162 553440 340886
rect 553400 338156 553452 338162
rect 553400 338098 553452 338104
rect 552664 334008 552716 334014
rect 552664 333950 552716 333956
rect 558828 334008 558880 334014
rect 558828 333950 558880 333956
rect 558840 331498 558868 333950
rect 556804 331492 556856 331498
rect 556804 331434 556856 331440
rect 558828 331492 558880 331498
rect 558828 331434 558880 331440
rect 551376 328160 551428 328166
rect 551376 328102 551428 328108
rect 552664 325372 552716 325378
rect 552664 325314 552716 325320
rect 552676 322998 552704 325314
rect 556816 324358 556844 331434
rect 559576 325378 559604 348366
rect 561048 343670 561076 350542
rect 564440 349852 564492 349858
rect 564440 349794 564492 349800
rect 564452 347478 564480 349794
rect 561680 347472 561732 347478
rect 561680 347414 561732 347420
rect 564440 347472 564492 347478
rect 564440 347414 564492 347420
rect 561692 343670 561720 347414
rect 559656 343664 559708 343670
rect 559656 343606 559708 343612
rect 561036 343664 561088 343670
rect 561036 343606 561088 343612
rect 561680 343664 561732 343670
rect 561680 343606 561732 343612
rect 559668 327758 559696 343606
rect 566476 338706 566504 371690
rect 566568 368490 566596 391954
rect 567384 382288 567436 382294
rect 567384 382230 567436 382236
rect 567396 377738 567424 382230
rect 566648 377732 566700 377738
rect 566648 377674 566700 377680
rect 567384 377732 567436 377738
rect 567384 377674 567436 377680
rect 566660 369918 566688 377674
rect 569236 371754 569264 394606
rect 574100 390652 574152 390658
rect 574100 390594 574152 390600
rect 574112 387190 574140 390594
rect 571984 387184 572036 387190
rect 571984 387126 572036 387132
rect 574100 387184 574152 387190
rect 574100 387126 574152 387132
rect 571996 382294 572024 387126
rect 576216 385076 576268 385082
rect 576216 385018 576268 385024
rect 576228 382294 576256 385018
rect 571984 382288 572036 382294
rect 571984 382230 572036 382236
rect 574100 382288 574152 382294
rect 574100 382230 574152 382236
rect 576216 382288 576268 382294
rect 576216 382230 576268 382236
rect 574112 376378 574140 382230
rect 570972 376372 571024 376378
rect 570972 376314 571024 376320
rect 574100 376372 574152 376378
rect 574100 376314 574152 376320
rect 569224 371748 569276 371754
rect 569224 371690 569276 371696
rect 570984 371618 571012 376314
rect 568764 371612 568816 371618
rect 568764 371554 568816 371560
rect 570972 371612 571024 371618
rect 570972 371554 571024 371560
rect 568776 369918 568804 371554
rect 566648 369912 566700 369918
rect 566648 369854 566700 369860
rect 568764 369912 568816 369918
rect 568764 369854 568816 369860
rect 566556 368484 566608 368490
rect 566556 368426 566608 368432
rect 576860 356108 576912 356114
rect 576860 356050 576912 356056
rect 574744 354748 574796 354754
rect 574744 354690 574796 354696
rect 571984 353456 572036 353462
rect 571984 353398 572036 353404
rect 571996 349858 572024 353398
rect 571984 349852 572036 349858
rect 571984 349794 572036 349800
rect 574756 347478 574784 354690
rect 576872 353462 576900 356050
rect 577516 354754 577544 400182
rect 577608 390658 577636 403514
rect 580920 400246 580948 404767
rect 580908 400240 580960 400246
rect 580908 400182 580960 400188
rect 579618 393000 579674 393009
rect 579618 392935 579674 392944
rect 579632 392018 579660 392935
rect 577872 392012 577924 392018
rect 577872 391954 577924 391960
rect 579620 392012 579672 392018
rect 579620 391954 579672 391960
rect 577596 390652 577648 390658
rect 577596 390594 577648 390600
rect 577884 385082 577912 391954
rect 577872 385076 577924 385082
rect 577872 385018 577924 385024
rect 579526 369608 579582 369617
rect 579526 369543 579582 369552
rect 579540 367130 579568 369543
rect 577596 367124 577648 367130
rect 577596 367066 577648 367072
rect 579528 367124 579580 367130
rect 579528 367066 579580 367072
rect 577504 354748 577556 354754
rect 577504 354690 577556 354696
rect 576860 353456 576912 353462
rect 576860 353398 576912 353404
rect 573364 347472 573416 347478
rect 573364 347414 573416 347420
rect 574744 347472 574796 347478
rect 574744 347414 574796 347420
rect 571432 340944 571484 340950
rect 571432 340886 571484 340892
rect 563428 338700 563480 338706
rect 563428 338642 563480 338648
rect 566464 338700 566516 338706
rect 566464 338642 566516 338648
rect 563440 336666 563468 338642
rect 561772 336660 561824 336666
rect 561772 336602 561824 336608
rect 563428 336660 563480 336666
rect 563428 336602 563480 336608
rect 561784 334014 561812 336602
rect 571444 336394 571472 340886
rect 570972 336388 571024 336394
rect 570972 336330 571024 336336
rect 571432 336388 571484 336394
rect 571432 336330 571484 336336
rect 561772 334008 561824 334014
rect 561772 333950 561824 333956
rect 570984 331362 571012 336330
rect 567844 331356 567896 331362
rect 567844 331298 567896 331304
rect 570972 331356 571024 331362
rect 570972 331298 571024 331304
rect 567856 330138 567884 331298
rect 565084 330132 565136 330138
rect 565084 330074 565136 330080
rect 567844 330132 567896 330138
rect 567844 330074 567896 330080
rect 559656 327752 559708 327758
rect 559656 327694 559708 327700
rect 559564 325372 559616 325378
rect 559564 325314 559616 325320
rect 553400 324352 553452 324358
rect 553400 324294 553452 324300
rect 556804 324352 556856 324358
rect 556804 324294 556856 324300
rect 552664 322992 552716 322998
rect 552664 322934 552716 322940
rect 551284 320748 551336 320754
rect 551284 320690 551336 320696
rect 549168 319796 549220 319802
rect 549168 319738 549220 319744
rect 553412 319530 553440 324294
rect 549904 319524 549956 319530
rect 549904 319466 549956 319472
rect 553400 319524 553452 319530
rect 553400 319466 553452 319472
rect 549916 311030 549944 319466
rect 565096 314702 565124 330074
rect 572720 317076 572772 317082
rect 572720 317018 572772 317024
rect 560944 314696 560996 314702
rect 560944 314638 560996 314644
rect 565084 314696 565136 314702
rect 565084 314638 565136 314644
rect 549904 311024 549956 311030
rect 549904 310966 549956 310972
rect 557540 307760 557592 307766
rect 557540 307702 557592 307708
rect 540980 305040 541032 305046
rect 540980 304982 541032 304988
rect 543096 305040 543148 305046
rect 543096 304982 543148 304988
rect 546500 305040 546552 305046
rect 546500 304982 546552 304988
rect 548524 305040 548576 305046
rect 548524 304982 548576 304988
rect 540992 302274 541020 304982
rect 540900 302246 541020 302274
rect 536840 301028 536892 301034
rect 536840 300970 536892 300976
rect 539692 301028 539744 301034
rect 539692 300970 539744 300976
rect 536852 300354 536880 300970
rect 540900 300422 540928 302246
rect 546512 300490 546540 304982
rect 557552 302802 557580 307702
rect 553400 302796 553452 302802
rect 553400 302738 553452 302744
rect 557540 302796 557592 302802
rect 557540 302738 557592 302744
rect 553412 300558 553440 302738
rect 560956 302394 560984 314638
rect 567936 311840 567988 311846
rect 567936 311782 567988 311788
rect 567948 310010 567976 311782
rect 563060 310004 563112 310010
rect 563060 309946 563112 309952
rect 567936 310004 567988 310010
rect 567936 309946 567988 309952
rect 563072 307834 563100 309946
rect 572732 309194 572760 317018
rect 573376 311914 573404 347414
rect 577608 345098 577636 367066
rect 579526 357912 579582 357921
rect 579526 357847 579582 357856
rect 579540 356114 579568 357847
rect 579528 356108 579580 356114
rect 579528 356050 579580 356056
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 574100 345092 574152 345098
rect 574100 345034 574152 345040
rect 577596 345092 577648 345098
rect 577596 345034 577648 345040
rect 574112 340950 574140 345034
rect 574100 340944 574152 340950
rect 574100 340886 574152 340892
rect 580184 340202 580212 346015
rect 578884 340196 578936 340202
rect 578884 340138 578936 340144
rect 580172 340196 580224 340202
rect 580172 340138 580224 340144
rect 578896 328438 578924 340138
rect 576860 328432 576912 328438
rect 576860 328374 576912 328380
rect 578884 328432 578936 328438
rect 578884 328374 578936 328380
rect 576872 321586 576900 328374
rect 580262 322688 580318 322697
rect 580262 322623 580318 322632
rect 576780 321558 576900 321586
rect 576780 318850 576808 321558
rect 574836 318844 574888 318850
rect 574836 318786 574888 318792
rect 576768 318844 576820 318850
rect 576768 318786 576820 318792
rect 574848 317082 574876 318786
rect 574836 317076 574888 317082
rect 574836 317018 574888 317024
rect 573364 311908 573416 311914
rect 573364 311850 573416 311856
rect 569960 309188 570012 309194
rect 569960 309130 570012 309136
rect 572720 309188 572772 309194
rect 572720 309130 572772 309136
rect 569972 308446 570000 309130
rect 565084 308440 565136 308446
rect 565084 308382 565136 308388
rect 569960 308440 570012 308446
rect 569960 308382 570012 308388
rect 563060 307828 563112 307834
rect 563060 307770 563112 307776
rect 559104 302388 559156 302394
rect 559104 302330 559156 302336
rect 560944 302388 560996 302394
rect 560944 302330 560996 302336
rect 559116 300626 559144 302330
rect 565096 300694 565124 308382
rect 580276 300830 580304 322623
rect 580354 310856 580410 310865
rect 580354 310791 580410 310800
rect 580264 300824 580316 300830
rect 580264 300766 580316 300772
rect 580368 300762 580396 310791
rect 580356 300756 580408 300762
rect 580356 300698 580408 300704
rect 565084 300688 565136 300694
rect 565084 300630 565136 300636
rect 559104 300620 559156 300626
rect 559104 300562 559156 300568
rect 553400 300552 553452 300558
rect 553400 300494 553452 300500
rect 546500 300484 546552 300490
rect 546500 300426 546552 300432
rect 540888 300416 540940 300422
rect 540888 300358 540940 300364
rect 536840 300348 536892 300354
rect 536840 300290 536892 300296
rect 532332 300280 532384 300286
rect 532332 300222 532384 300228
rect 516140 300212 516192 300218
rect 516140 300154 516192 300160
rect 514760 300144 514812 300150
rect 62224 300070 62882 300098
rect 61106 299568 61162 299577
rect 61106 299503 61162 299512
rect 61120 298058 61148 299503
rect 61028 298030 61148 298058
rect 61028 292602 61056 298030
rect 62028 297016 62080 297022
rect 62028 296958 62080 296964
rect 61016 292596 61068 292602
rect 61016 292538 61068 292544
rect 61108 292528 61160 292534
rect 61108 292470 61160 292476
rect 61120 288454 61148 292470
rect 61016 288448 61068 288454
rect 61016 288390 61068 288396
rect 61108 288448 61160 288454
rect 61108 288390 61160 288396
rect 61028 285002 61056 288390
rect 61028 284974 61148 285002
rect 61120 273290 61148 284974
rect 60740 273284 60792 273290
rect 60740 273226 60792 273232
rect 61108 273284 61160 273290
rect 61108 273226 61160 273232
rect 60752 273170 60780 273226
rect 60752 273142 60872 273170
rect 60844 263650 60872 273142
rect 60844 263622 60964 263650
rect 60936 263566 60964 263622
rect 60924 263560 60976 263566
rect 60924 263502 60976 263508
rect 61108 263560 61160 263566
rect 61108 263502 61160 263508
rect 61120 260846 61148 263502
rect 60832 260840 60884 260846
rect 60832 260782 60884 260788
rect 61108 260840 61160 260846
rect 61108 260782 61160 260788
rect 60844 251258 60872 260782
rect 60832 251252 60884 251258
rect 60832 251194 60884 251200
rect 61016 251252 61068 251258
rect 61016 251194 61068 251200
rect 61028 244202 61056 251194
rect 60844 244174 61056 244202
rect 60844 234682 60872 244174
rect 60752 234654 60872 234682
rect 60752 225010 60780 234654
rect 60740 225004 60792 225010
rect 60740 224946 60792 224952
rect 60924 224868 60976 224874
rect 60924 224810 60976 224816
rect 60936 215354 60964 224810
rect 60740 215348 60792 215354
rect 60740 215290 60792 215296
rect 60924 215348 60976 215354
rect 60924 215290 60976 215296
rect 60752 207754 60780 215290
rect 60660 207726 60780 207754
rect 60660 205562 60688 207726
rect 60648 205556 60700 205562
rect 60648 205498 60700 205504
rect 60924 205556 60976 205562
rect 60924 205498 60976 205504
rect 60936 196042 60964 205498
rect 60924 196036 60976 196042
rect 60924 195978 60976 195984
rect 61016 195968 61068 195974
rect 61016 195910 61068 195916
rect 61028 186266 61056 195910
rect 60936 186238 61056 186266
rect 60936 181558 60964 186238
rect 60924 181552 60976 181558
rect 60924 181494 60976 181500
rect 61108 181552 61160 181558
rect 61108 181494 61160 181500
rect 61120 173913 61148 181494
rect 60922 173904 60978 173913
rect 60922 173839 60978 173848
rect 61106 173904 61162 173913
rect 61106 173839 61162 173848
rect 60936 167006 60964 173839
rect 60924 167000 60976 167006
rect 60924 166942 60976 166948
rect 61108 167000 61160 167006
rect 61108 166942 61160 166948
rect 61120 164234 61148 166942
rect 61120 164206 61240 164234
rect 59360 158704 59412 158710
rect 59360 158646 59412 158652
rect 61212 157486 61240 164206
rect 61200 157480 61252 157486
rect 61200 157422 61252 157428
rect 61016 157276 61068 157282
rect 61016 157218 61068 157224
rect 61028 153202 61056 157218
rect 61016 153196 61068 153202
rect 61016 153138 61068 153144
rect 61200 153196 61252 153202
rect 61200 153138 61252 153144
rect 61212 143585 61240 153138
rect 60922 143576 60978 143585
rect 60922 143511 60978 143520
rect 61198 143576 61254 143585
rect 61198 143511 61254 143520
rect 60936 138038 60964 143511
rect 60924 138032 60976 138038
rect 60924 137974 60976 137980
rect 61016 137964 61068 137970
rect 61016 137906 61068 137912
rect 61028 135232 61056 137906
rect 60844 135204 61056 135232
rect 60844 125610 60872 135204
rect 60844 125582 60964 125610
rect 60936 118726 60964 125582
rect 60924 118720 60976 118726
rect 60924 118662 60976 118668
rect 61016 118652 61068 118658
rect 61016 118594 61068 118600
rect 61028 106321 61056 118594
rect 60738 106312 60794 106321
rect 60738 106247 60794 106256
rect 61014 106312 61070 106321
rect 61014 106247 61070 106256
rect 60752 99414 60780 106247
rect 60740 99408 60792 99414
rect 60740 99350 60792 99356
rect 61108 99272 61160 99278
rect 61108 99214 61160 99220
rect 61120 89706 61148 99214
rect 61028 89678 61148 89706
rect 61028 86970 61056 89678
rect 60740 86964 60792 86970
rect 60740 86906 60792 86912
rect 61016 86964 61068 86970
rect 61016 86906 61068 86912
rect 60752 77314 60780 86906
rect 60740 77308 60792 77314
rect 60740 77250 60792 77256
rect 60924 77308 60976 77314
rect 60924 77250 60976 77256
rect 60936 75886 60964 77250
rect 60648 75880 60700 75886
rect 60648 75822 60700 75828
rect 60924 75880 60976 75886
rect 60924 75822 60976 75828
rect 60660 70258 60688 75822
rect 60660 70230 60872 70258
rect 60844 60738 60872 70230
rect 60844 60722 60964 60738
rect 60844 60716 60976 60722
rect 60844 60710 60924 60716
rect 60924 60658 60976 60664
rect 61108 60716 61160 60722
rect 61108 60658 61160 60664
rect 61120 57934 61148 60658
rect 60832 57928 60884 57934
rect 60832 57870 60884 57876
rect 61108 57928 61160 57934
rect 61108 57870 61160 57876
rect 60844 48346 60872 57870
rect 60832 48340 60884 48346
rect 60832 48282 60884 48288
rect 61016 48340 61068 48346
rect 61016 48282 61068 48288
rect 61028 41426 61056 48282
rect 60936 41398 61056 41426
rect 60936 31890 60964 41398
rect 60924 31884 60976 31890
rect 60924 31826 60976 31832
rect 60924 31748 60976 31754
rect 60924 31690 60976 31696
rect 60936 22114 60964 31690
rect 60752 22086 60964 22114
rect 59268 17944 59320 17950
rect 59268 17886 59320 17892
rect 60752 12510 60780 22086
rect 60740 12504 60792 12510
rect 60740 12446 60792 12452
rect 60832 12368 60884 12374
rect 60832 12310 60884 12316
rect 60844 9654 60872 12310
rect 59176 9648 59228 9654
rect 59176 9590 59228 9596
rect 60832 9648 60884 9654
rect 60832 9590 60884 9596
rect 52828 4752 52880 4758
rect 52828 4694 52880 4700
rect 51816 3052 51868 3058
rect 51816 2994 51868 3000
rect 52840 480 52868 4694
rect 58808 4412 58860 4418
rect 58808 4354 58860 4360
rect 55220 4344 55272 4350
rect 55220 4286 55272 4292
rect 54024 3052 54076 3058
rect 54024 2994 54076 3000
rect 54036 480 54064 2994
rect 55232 480 55260 4286
rect 57612 3188 57664 3194
rect 57612 3130 57664 3136
rect 56416 3120 56468 3126
rect 56416 3062 56468 3068
rect 56428 480 56456 3062
rect 57624 480 57652 3130
rect 58820 480 58848 4354
rect 59188 3398 59216 9590
rect 60004 6452 60056 6458
rect 60004 6394 60056 6400
rect 59176 3392 59228 3398
rect 59176 3334 59228 3340
rect 60016 480 60044 6394
rect 62040 4146 62068 296958
rect 61108 4140 61160 4146
rect 61108 4082 61160 4088
rect 61200 4140 61252 4146
rect 61200 4082 61252 4088
rect 62028 4140 62080 4146
rect 62028 4082 62080 4088
rect 61120 3466 61148 4082
rect 61108 3460 61160 3466
rect 61108 3402 61160 3408
rect 61212 480 61240 4082
rect 62224 3330 62252 300070
rect 64800 297974 64828 300084
rect 66272 300070 66746 300098
rect 64788 297968 64840 297974
rect 64788 297910 64840 297916
rect 64788 297084 64840 297090
rect 64788 297026 64840 297032
rect 62396 4480 62448 4486
rect 62396 4422 62448 4428
rect 62212 3324 62264 3330
rect 62212 3266 62264 3272
rect 62408 480 62436 4422
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64144 3392 64196 3398
rect 64144 3334 64196 3340
rect 63604 480 63632 3334
rect 64156 3262 64184 3334
rect 64144 3256 64196 3262
rect 64144 3198 64196 3204
rect 64800 480 64828 297026
rect 65524 5296 65576 5302
rect 65524 5238 65576 5244
rect 65536 4758 65564 5238
rect 65524 4752 65576 4758
rect 65524 4694 65576 4700
rect 65984 4548 66036 4554
rect 65984 4490 66036 4496
rect 65996 480 66024 4490
rect 66272 3466 66300 300070
rect 68664 298110 68692 300084
rect 68652 298104 68704 298110
rect 68652 298046 68704 298052
rect 70596 297362 70624 300084
rect 71792 300070 72542 300098
rect 70584 297356 70636 297362
rect 70584 297298 70636 297304
rect 67548 297152 67600 297158
rect 67548 297094 67600 297100
rect 67560 280430 67588 297094
rect 67548 280424 67600 280430
rect 67548 280366 67600 280372
rect 67548 280288 67600 280294
rect 67548 280230 67600 280236
rect 67560 240145 67588 280230
rect 67362 240136 67418 240145
rect 67362 240071 67418 240080
rect 67546 240136 67602 240145
rect 67546 240071 67602 240080
rect 67376 231878 67404 240071
rect 67364 231872 67416 231878
rect 67364 231814 67416 231820
rect 67364 231736 67416 231742
rect 67364 231678 67416 231684
rect 67376 230450 67404 231678
rect 67272 230444 67324 230450
rect 67272 230386 67324 230392
rect 67364 230444 67416 230450
rect 67364 230386 67416 230392
rect 67284 220862 67312 230386
rect 67272 220856 67324 220862
rect 67272 220798 67324 220804
rect 67548 220856 67600 220862
rect 67548 220798 67600 220804
rect 67560 212566 67588 220798
rect 67548 212560 67600 212566
rect 67548 212502 67600 212508
rect 67456 212492 67508 212498
rect 67456 212434 67508 212440
rect 67468 211138 67496 212434
rect 67456 211132 67508 211138
rect 67456 211074 67508 211080
rect 67548 211132 67600 211138
rect 67548 211074 67600 211080
rect 67560 202910 67588 211074
rect 67548 202904 67600 202910
rect 67548 202846 67600 202852
rect 67456 202836 67508 202842
rect 67456 202778 67508 202784
rect 67468 201498 67496 202778
rect 67468 201470 67588 201498
rect 67560 177313 67588 201470
rect 67546 177304 67602 177313
rect 67546 177239 67602 177248
rect 67546 164248 67602 164257
rect 67546 164183 67602 164192
rect 67560 126041 67588 164183
rect 67546 126032 67602 126041
rect 67546 125967 67602 125976
rect 67546 125624 67602 125633
rect 67546 125559 67602 125568
rect 67560 115938 67588 125559
rect 67456 115932 67508 115938
rect 67456 115874 67508 115880
rect 67548 115932 67600 115938
rect 67548 115874 67600 115880
rect 67468 114510 67496 115874
rect 67272 114504 67324 114510
rect 67272 114446 67324 114452
rect 67456 114504 67508 114510
rect 67456 114446 67508 114452
rect 67284 104922 67312 114446
rect 67272 104916 67324 104922
rect 67272 104858 67324 104864
rect 67548 104916 67600 104922
rect 67548 104858 67600 104864
rect 67560 57934 67588 104858
rect 67456 57928 67508 57934
rect 67456 57870 67508 57876
rect 67548 57928 67600 57934
rect 67548 57870 67600 57876
rect 67468 56574 67496 57870
rect 67272 56568 67324 56574
rect 67272 56510 67324 56516
rect 67456 56568 67508 56574
rect 67456 56510 67508 56516
rect 67284 46986 67312 56510
rect 67272 46980 67324 46986
rect 67272 46922 67324 46928
rect 67548 46980 67600 46986
rect 67548 46922 67600 46928
rect 67560 37330 67588 46922
rect 67456 37324 67508 37330
rect 67456 37266 67508 37272
rect 67548 37324 67600 37330
rect 67548 37266 67600 37272
rect 67468 37233 67496 37266
rect 67454 37224 67510 37233
rect 67454 37159 67510 37168
rect 67730 37224 67786 37233
rect 67730 37159 67786 37168
rect 67744 27674 67772 37159
rect 67548 27668 67600 27674
rect 67548 27610 67600 27616
rect 67732 27668 67784 27674
rect 67732 27610 67784 27616
rect 67560 19310 67588 27610
rect 67548 19304 67600 19310
rect 67548 19246 67600 19252
rect 66996 19236 67048 19242
rect 66996 19178 67048 19184
rect 67008 4842 67036 19178
rect 71792 5506 71820 300070
rect 74448 297288 74500 297294
rect 74448 297230 74500 297236
rect 72976 297220 73028 297226
rect 72976 297162 73028 297168
rect 71780 5500 71832 5506
rect 71780 5442 71832 5448
rect 71872 5500 71924 5506
rect 71872 5442 71924 5448
rect 71884 5302 71912 5442
rect 71872 5296 71924 5302
rect 71872 5238 71924 5244
rect 67008 4814 67220 4842
rect 66260 3460 66312 3466
rect 66260 3402 66312 3408
rect 67192 480 67220 4814
rect 69480 4616 69532 4622
rect 69480 4558 69532 4564
rect 68284 4140 68336 4146
rect 68284 4082 68336 4088
rect 68296 480 68324 4082
rect 68650 3496 68706 3505
rect 68650 3431 68706 3440
rect 68664 3330 68692 3431
rect 68652 3324 68704 3330
rect 68652 3266 68704 3272
rect 69492 480 69520 4558
rect 72988 3466 73016 297162
rect 73068 4684 73120 4690
rect 73068 4626 73120 4632
rect 71872 3460 71924 3466
rect 71872 3402 71924 3408
rect 72976 3460 73028 3466
rect 72976 3402 73028 3408
rect 70676 1148 70728 1154
rect 70676 1090 70728 1096
rect 70688 480 70716 1090
rect 71884 480 71912 3402
rect 73080 480 73108 4626
rect 73344 4140 73396 4146
rect 73344 4082 73396 4088
rect 73252 3392 73304 3398
rect 73252 3334 73304 3340
rect 73264 1154 73292 3334
rect 73356 3330 73384 4082
rect 74460 3448 74488 297230
rect 74552 4078 74580 300084
rect 76484 297906 76512 300084
rect 78416 298042 78444 300084
rect 80072 300070 80362 300098
rect 81452 300070 82294 300098
rect 78404 298036 78456 298042
rect 78404 297978 78456 297984
rect 76472 297900 76524 297906
rect 76472 297842 76524 297848
rect 79968 297356 80020 297362
rect 79968 297298 80020 297304
rect 77206 76256 77262 76265
rect 77206 76191 77262 76200
rect 77220 75857 77248 76191
rect 77206 75848 77262 75857
rect 77206 75783 77262 75792
rect 77206 40352 77262 40361
rect 77206 40287 77262 40296
rect 77220 39953 77248 40287
rect 77206 39944 77262 39953
rect 77206 39879 77262 39888
rect 76656 4752 76708 4758
rect 76656 4694 76708 4700
rect 74540 4072 74592 4078
rect 74540 4014 74592 4020
rect 75460 4004 75512 4010
rect 75460 3946 75512 3952
rect 74630 3632 74686 3641
rect 74630 3567 74686 3576
rect 74644 3534 74672 3567
rect 74632 3528 74684 3534
rect 74632 3470 74684 3476
rect 74276 3420 74488 3448
rect 73344 3324 73396 3330
rect 73344 3266 73396 3272
rect 73252 1148 73304 1154
rect 73252 1090 73304 1096
rect 74276 480 74304 3420
rect 75472 480 75500 3946
rect 76668 480 76696 4694
rect 77852 4072 77904 4078
rect 77852 4014 77904 4020
rect 78954 4040 79010 4049
rect 77864 480 77892 4014
rect 79980 4010 80008 297298
rect 80072 5438 80100 300070
rect 80244 5500 80296 5506
rect 80244 5442 80296 5448
rect 80060 5432 80112 5438
rect 80060 5374 80112 5380
rect 78954 3975 78956 3984
rect 79008 3975 79010 3984
rect 79048 4004 79100 4010
rect 78956 3946 79008 3952
rect 79048 3946 79100 3952
rect 79968 4004 80020 4010
rect 79968 3946 80020 3952
rect 79060 480 79088 3946
rect 80256 480 80284 5442
rect 81452 4146 81480 300070
rect 82728 298104 82780 298110
rect 82728 298046 82780 298052
rect 81440 4140 81492 4146
rect 81440 4082 81492 4088
rect 82636 4072 82688 4078
rect 82636 4014 82688 4020
rect 81440 4004 81492 4010
rect 81440 3946 81492 3952
rect 81452 480 81480 3946
rect 82648 480 82676 4014
rect 82740 4010 82768 298046
rect 84212 297702 84240 300084
rect 86236 297838 86264 300084
rect 86972 300070 88182 300098
rect 89732 300070 90114 300098
rect 86868 298036 86920 298042
rect 86868 297978 86920 297984
rect 86224 297832 86276 297838
rect 86224 297774 86276 297780
rect 84200 297696 84252 297702
rect 84200 297638 84252 297644
rect 86880 29306 86908 297978
rect 86868 29300 86920 29306
rect 86868 29242 86920 29248
rect 86868 29164 86920 29170
rect 86868 29106 86920 29112
rect 83752 5494 83964 5522
rect 83752 5438 83780 5494
rect 83740 5432 83792 5438
rect 83740 5374 83792 5380
rect 83832 5432 83884 5438
rect 83832 5374 83884 5380
rect 83936 5386 83964 5494
rect 83004 4140 83056 4146
rect 83004 4082 83056 4088
rect 83016 4049 83044 4082
rect 83002 4040 83058 4049
rect 82728 4004 82780 4010
rect 83002 3975 83058 3984
rect 82728 3946 82780 3952
rect 83844 480 83872 5374
rect 83936 5358 84148 5386
rect 84120 5302 84148 5358
rect 84108 5296 84160 5302
rect 84108 5238 84160 5244
rect 86038 4040 86094 4049
rect 86038 3975 86094 3984
rect 86052 3942 86080 3975
rect 86880 3942 86908 29106
rect 86972 5370 87000 300070
rect 89628 297968 89680 297974
rect 89628 297910 89680 297916
rect 89536 76152 89588 76158
rect 89534 76120 89536 76129
rect 89588 76120 89590 76129
rect 89534 76055 89590 76064
rect 89534 40216 89590 40225
rect 89534 40151 89536 40160
rect 89588 40151 89590 40160
rect 89536 40122 89588 40128
rect 86960 5364 87012 5370
rect 86960 5306 87012 5312
rect 87328 5364 87380 5370
rect 87328 5306 87380 5312
rect 86040 3936 86092 3942
rect 86040 3878 86092 3884
rect 86132 3936 86184 3942
rect 86132 3878 86184 3884
rect 86868 3936 86920 3942
rect 86868 3878 86920 3884
rect 84934 3768 84990 3777
rect 84934 3703 84990 3712
rect 84014 3632 84070 3641
rect 84014 3567 84070 3576
rect 84028 3534 84056 3567
rect 84016 3528 84068 3534
rect 84016 3470 84068 3476
rect 84106 3496 84162 3505
rect 84106 3431 84108 3440
rect 84160 3431 84162 3440
rect 84108 3402 84160 3408
rect 84948 480 84976 3703
rect 86144 480 86172 3878
rect 87340 480 87368 5306
rect 89640 3942 89668 297910
rect 89732 4049 89760 300070
rect 92032 297634 92060 300084
rect 93768 297832 93820 297838
rect 93768 297774 93820 297780
rect 92020 297628 92072 297634
rect 92020 297570 92072 297576
rect 89812 76152 89864 76158
rect 89810 76120 89812 76129
rect 89864 76120 89866 76129
rect 89810 76055 89866 76064
rect 91742 40216 91798 40225
rect 91742 40151 91744 40160
rect 91796 40151 91798 40160
rect 91744 40122 91796 40128
rect 91742 29608 91798 29617
rect 91742 29543 91798 29552
rect 91756 29209 91784 29543
rect 91742 29200 91798 29209
rect 91742 29135 91798 29144
rect 90914 5264 90970 5273
rect 90914 5199 90970 5208
rect 89718 4040 89774 4049
rect 89718 3975 89774 3984
rect 88524 3936 88576 3942
rect 88524 3878 88576 3884
rect 89628 3936 89680 3942
rect 89628 3878 89680 3884
rect 89720 3936 89772 3942
rect 89720 3878 89772 3884
rect 88536 480 88564 3878
rect 89732 480 89760 3878
rect 90928 480 90956 5199
rect 93780 3942 93808 297774
rect 93964 297566 93992 300084
rect 95252 300070 95910 300098
rect 96632 300070 97934 300098
rect 93952 297560 94004 297566
rect 93952 297502 94004 297508
rect 93860 5568 93912 5574
rect 93860 5510 93912 5516
rect 93872 5302 93900 5510
rect 93860 5296 93912 5302
rect 93860 5238 93912 5244
rect 95252 5234 95280 300070
rect 96528 297900 96580 297906
rect 96528 297842 96580 297848
rect 95240 5228 95292 5234
rect 95240 5170 95292 5176
rect 94502 5128 94558 5137
rect 94502 5063 94558 5072
rect 93216 3936 93268 3942
rect 93214 3904 93216 3913
rect 93308 3936 93360 3942
rect 93268 3904 93270 3913
rect 93308 3878 93360 3884
rect 93768 3936 93820 3942
rect 93860 3936 93912 3942
rect 93768 3878 93820 3884
rect 93858 3904 93860 3913
rect 93912 3904 93914 3913
rect 93214 3839 93270 3848
rect 92110 3632 92166 3641
rect 92110 3567 92166 3576
rect 92124 480 92152 3567
rect 93320 480 93348 3878
rect 93858 3839 93914 3848
rect 93952 3528 94004 3534
rect 93952 3470 94004 3476
rect 93860 3460 93912 3466
rect 93860 3402 93912 3408
rect 93872 3369 93900 3402
rect 93858 3360 93914 3369
rect 93858 3295 93914 3304
rect 93964 3233 93992 3470
rect 93950 3224 94006 3233
rect 93950 3159 94006 3168
rect 94516 480 94544 5063
rect 95514 3904 95570 3913
rect 95514 3839 95516 3848
rect 95568 3839 95570 3848
rect 95516 3810 95568 3816
rect 96540 3806 96568 297842
rect 96632 3913 96660 300070
rect 99852 297498 99880 300084
rect 100668 297696 100720 297702
rect 100668 297638 100720 297644
rect 99840 297492 99892 297498
rect 99840 297434 99892 297440
rect 99472 5568 99524 5574
rect 99472 5510 99524 5516
rect 99484 5234 99512 5510
rect 98092 5228 98144 5234
rect 98092 5170 98144 5176
rect 99472 5228 99524 5234
rect 99472 5170 99524 5176
rect 96618 3904 96674 3913
rect 96618 3839 96674 3848
rect 96896 3868 96948 3874
rect 96896 3810 96948 3816
rect 95700 3800 95752 3806
rect 95700 3742 95752 3748
rect 96528 3800 96580 3806
rect 96528 3742 96580 3748
rect 95712 480 95740 3742
rect 96908 480 96936 3810
rect 98104 480 98132 5170
rect 99472 3528 99524 3534
rect 99286 3496 99342 3505
rect 99472 3470 99524 3476
rect 99286 3431 99342 3440
rect 99380 3460 99432 3466
rect 99300 480 99328 3431
rect 99380 3402 99432 3408
rect 99392 3369 99420 3402
rect 99378 3360 99434 3369
rect 99378 3295 99434 3304
rect 99484 3233 99512 3470
rect 99470 3224 99526 3233
rect 99470 3159 99526 3168
rect 100680 626 100708 297638
rect 101784 297430 101812 300084
rect 103532 300070 103730 300098
rect 104912 300070 105662 300098
rect 107304 300070 107594 300098
rect 109052 300070 109526 300098
rect 110432 300070 111550 300098
rect 113192 300070 113482 300098
rect 114572 300070 115414 300098
rect 103428 297628 103480 297634
rect 103428 297570 103480 297576
rect 101772 297424 101824 297430
rect 101772 297366 101824 297372
rect 101586 4992 101642 5001
rect 101586 4927 101642 4936
rect 100496 598 100708 626
rect 100496 480 100524 598
rect 101600 480 101628 4927
rect 102690 3904 102746 3913
rect 102690 3839 102746 3848
rect 102704 3806 102732 3839
rect 103440 3806 103468 297570
rect 103532 5166 103560 300070
rect 103520 5160 103572 5166
rect 103520 5102 103572 5108
rect 104912 3913 104940 300070
rect 107304 296750 107332 300070
rect 107568 297560 107620 297566
rect 107568 297502 107620 297508
rect 107476 297492 107528 297498
rect 107476 297434 107528 297440
rect 107292 296744 107344 296750
rect 107292 296686 107344 296692
rect 105176 5228 105228 5234
rect 105176 5170 105228 5176
rect 104898 3904 104954 3913
rect 104898 3839 104954 3848
rect 102692 3800 102744 3806
rect 102692 3742 102744 3748
rect 102784 3800 102836 3806
rect 102784 3742 102836 3748
rect 103428 3800 103480 3806
rect 103428 3742 103480 3748
rect 102796 480 102824 3742
rect 103978 3360 104034 3369
rect 103978 3295 104034 3304
rect 103992 480 104020 3295
rect 105188 480 105216 5170
rect 106372 3800 106424 3806
rect 106372 3742 106424 3748
rect 106384 480 106412 3742
rect 107488 3618 107516 297434
rect 107580 3806 107608 297502
rect 108764 6384 108816 6390
rect 108764 6326 108816 6332
rect 107568 3800 107620 3806
rect 107568 3742 107620 3748
rect 107660 3800 107712 3806
rect 107660 3742 107712 3748
rect 107488 3590 107608 3618
rect 107672 3602 107700 3742
rect 107580 480 107608 3590
rect 107660 3596 107712 3602
rect 107660 3538 107712 3544
rect 108776 480 108804 6326
rect 109052 5658 109080 300070
rect 109052 5630 109172 5658
rect 108948 5568 109000 5574
rect 108948 5510 109000 5516
rect 109040 5568 109092 5574
rect 109040 5510 109092 5516
rect 108960 5302 108988 5510
rect 109052 5302 109080 5510
rect 108948 5296 109000 5302
rect 108948 5238 109000 5244
rect 109040 5296 109092 5302
rect 109040 5238 109092 5244
rect 109144 5098 109172 5630
rect 109132 5092 109184 5098
rect 109132 5034 109184 5040
rect 109866 3904 109922 3913
rect 109866 3839 109922 3848
rect 109880 3670 109908 3839
rect 110432 3738 110460 300070
rect 112352 6316 112404 6322
rect 112352 6258 112404 6264
rect 110420 3732 110472 3738
rect 110420 3674 110472 3680
rect 109868 3664 109920 3670
rect 109868 3606 109920 3612
rect 109960 3664 110012 3670
rect 109960 3606 110012 3612
rect 109972 480 110000 3606
rect 111156 3596 111208 3602
rect 111156 3538 111208 3544
rect 111168 480 111196 3538
rect 112364 480 112392 6258
rect 113192 3806 113220 300070
rect 114468 297424 114520 297430
rect 114468 297366 114520 297372
rect 114480 3806 114508 297366
rect 114572 5030 114600 300070
rect 115846 297664 115902 297673
rect 115846 297599 115902 297608
rect 114560 5024 114612 5030
rect 114560 4966 114612 4972
rect 115860 3806 115888 297599
rect 115940 76016 115992 76022
rect 115938 75984 115940 75993
rect 115992 75984 115994 75993
rect 115938 75919 115994 75928
rect 115940 40112 115992 40118
rect 115938 40080 115940 40089
rect 115992 40080 115994 40089
rect 115938 40015 115994 40024
rect 115940 29096 115992 29102
rect 115938 29064 115940 29073
rect 115992 29064 115994 29073
rect 115938 28999 115994 29008
rect 115940 6248 115992 6254
rect 115940 6190 115992 6196
rect 113180 3800 113232 3806
rect 113180 3742 113232 3748
rect 113548 3800 113600 3806
rect 113548 3742 113600 3748
rect 114468 3800 114520 3806
rect 114468 3742 114520 3748
rect 114744 3800 114796 3806
rect 114744 3742 114796 3748
rect 115848 3800 115900 3806
rect 115848 3742 115900 3748
rect 113560 480 113588 3742
rect 114756 480 114784 3742
rect 115952 480 115980 6190
rect 117332 3913 117360 300084
rect 118804 300070 119278 300098
rect 120092 300070 121210 300098
rect 122944 300070 123234 300098
rect 124784 300070 125166 300098
rect 126992 300070 127098 300098
rect 117318 3904 117374 3913
rect 117318 3839 117374 3848
rect 117136 3664 117188 3670
rect 117136 3606 117188 3612
rect 117148 480 117176 3606
rect 118240 3596 118292 3602
rect 118240 3538 118292 3544
rect 118252 480 118280 3538
rect 118804 3534 118832 300070
rect 118882 76256 118938 76265
rect 118882 76191 118938 76200
rect 118896 76022 118924 76191
rect 118884 76016 118936 76022
rect 118884 75958 118936 75964
rect 118882 40352 118938 40361
rect 118882 40287 118938 40296
rect 118896 40118 118924 40287
rect 118884 40112 118936 40118
rect 118884 40054 118936 40060
rect 119436 5092 119488 5098
rect 119436 5034 119488 5040
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 119448 480 119476 5034
rect 120092 4962 120120 300070
rect 121366 297528 121422 297537
rect 121366 297463 121422 297472
rect 120814 29336 120870 29345
rect 120814 29271 120870 29280
rect 120828 29102 120856 29271
rect 120816 29096 120868 29102
rect 120816 29038 120868 29044
rect 120080 4956 120132 4962
rect 120080 4898 120132 4904
rect 121380 3670 121408 297463
rect 122746 297392 122802 297401
rect 122746 297327 122802 297336
rect 122760 3670 122788 297327
rect 120632 3664 120684 3670
rect 120632 3606 120684 3612
rect 121368 3664 121420 3670
rect 121368 3606 121420 3612
rect 121828 3664 121880 3670
rect 121828 3606 121880 3612
rect 122748 3664 122800 3670
rect 122748 3606 122800 3612
rect 122840 3664 122892 3670
rect 122840 3606 122892 3612
rect 120644 480 120672 3606
rect 121840 480 121868 3606
rect 122656 3528 122708 3534
rect 122852 3482 122880 3606
rect 122708 3476 122880 3482
rect 122656 3470 122880 3476
rect 122668 3454 122880 3470
rect 122944 3466 122972 300070
rect 124784 296818 124812 300070
rect 124772 296812 124824 296818
rect 124772 296754 124824 296760
rect 124864 296812 124916 296818
rect 124864 296754 124916 296760
rect 123024 6180 123076 6186
rect 123024 6122 123076 6128
rect 122932 3460 122984 3466
rect 122932 3402 122984 3408
rect 123036 480 123064 6122
rect 124876 5166 124904 296754
rect 124864 5160 124916 5166
rect 124864 5102 124916 5108
rect 126612 4956 126664 4962
rect 126612 4898 126664 4904
rect 124220 3528 124272 3534
rect 124220 3470 124272 3476
rect 124232 480 124260 3470
rect 125416 3460 125468 3466
rect 125416 3402 125468 3408
rect 125428 480 125456 3402
rect 126624 480 126652 4898
rect 126992 4894 127020 300070
rect 129016 297770 129044 300084
rect 129844 300070 130962 300098
rect 132512 300070 132894 300098
rect 133984 300070 134918 300098
rect 129004 297764 129056 297770
rect 129004 297706 129056 297712
rect 128266 29336 128322 29345
rect 128266 29271 128322 29280
rect 128280 29186 128308 29271
rect 128450 29200 128506 29209
rect 128280 29158 128450 29186
rect 128450 29135 128506 29144
rect 127808 5160 127860 5166
rect 127808 5102 127860 5108
rect 126980 4888 127032 4894
rect 126980 4830 127032 4836
rect 127820 480 127848 5102
rect 129004 4956 129056 4962
rect 129004 4898 129056 4904
rect 129016 480 129044 4898
rect 129844 2854 129872 300070
rect 130200 5024 130252 5030
rect 130200 4966 130252 4972
rect 129832 2848 129884 2854
rect 129832 2790 129884 2796
rect 130212 480 130240 4966
rect 131394 4856 131450 4865
rect 132512 4826 132540 300070
rect 131394 4791 131450 4800
rect 132500 4820 132552 4826
rect 131408 480 131436 4791
rect 132500 4762 132552 4768
rect 132592 4820 132644 4826
rect 132592 4762 132644 4768
rect 132604 480 132632 4762
rect 133984 2922 134012 300070
rect 134524 297764 134576 297770
rect 134524 297706 134576 297712
rect 134536 5098 134564 297706
rect 136836 296886 136864 300084
rect 138032 300070 138782 300098
rect 139412 300070 140714 300098
rect 136824 296880 136876 296886
rect 136824 296822 136876 296828
rect 135166 76528 135222 76537
rect 135166 76463 135222 76472
rect 135180 76129 135208 76463
rect 135166 76120 135222 76129
rect 135166 76055 135222 76064
rect 135166 40624 135222 40633
rect 135166 40559 135222 40568
rect 135180 40225 135208 40559
rect 135166 40216 135222 40225
rect 135166 40151 135222 40160
rect 137204 5222 137600 5250
rect 137204 5098 137232 5222
rect 137376 5160 137428 5166
rect 137428 5108 137508 5114
rect 137376 5102 137508 5108
rect 134524 5092 134576 5098
rect 134524 5034 134576 5040
rect 134616 5092 134668 5098
rect 134616 5034 134668 5040
rect 137192 5092 137244 5098
rect 137388 5086 137508 5102
rect 137192 5034 137244 5040
rect 134628 4826 134656 5034
rect 137480 5030 137508 5086
rect 137468 5024 137520 5030
rect 137468 4966 137520 4972
rect 137572 4894 137600 5222
rect 137652 5160 137704 5166
rect 137652 5102 137704 5108
rect 137468 4888 137520 4894
rect 137468 4830 137520 4836
rect 137560 4888 137612 4894
rect 137560 4830 137612 4836
rect 134616 4820 134668 4826
rect 134616 4762 134668 4768
rect 134892 4820 134944 4826
rect 134892 4762 134944 4768
rect 133972 2916 134024 2922
rect 133972 2858 134024 2864
rect 134904 480 134932 4762
rect 137480 4706 137508 4830
rect 137664 4706 137692 5102
rect 137480 4678 137692 4706
rect 138032 4214 138060 300070
rect 138020 4208 138072 4214
rect 138020 4150 138072 4156
rect 139412 2990 139440 300070
rect 142632 296954 142660 300084
rect 143552 300070 144578 300098
rect 142620 296948 142672 296954
rect 142620 296890 142672 296896
rect 140042 76392 140098 76401
rect 140042 76327 140098 76336
rect 140056 75993 140084 76327
rect 140042 75984 140098 75993
rect 140042 75919 140098 75928
rect 140042 40488 140098 40497
rect 140042 40423 140098 40432
rect 140056 40089 140084 40423
rect 140042 40080 140098 40089
rect 140042 40015 140098 40024
rect 143446 29472 143502 29481
rect 143446 29407 143502 29416
rect 143460 29073 143488 29407
rect 143446 29064 143502 29073
rect 143446 28999 143502 29008
rect 143552 4282 143580 300070
rect 146588 296818 146616 300084
rect 147692 300070 148534 300098
rect 146576 296812 146628 296818
rect 146576 296754 146628 296760
rect 147588 76152 147640 76158
rect 147586 76120 147588 76129
rect 147640 76120 147642 76129
rect 147586 76055 147642 76064
rect 147588 40248 147640 40254
rect 147586 40216 147588 40225
rect 147640 40216 147642 40225
rect 147586 40151 147642 40160
rect 147588 29232 147640 29238
rect 147586 29200 147588 29209
rect 147640 29200 147642 29209
rect 147586 29135 147642 29144
rect 143540 4276 143592 4282
rect 143540 4218 143592 4224
rect 147692 3058 147720 300070
rect 150452 4350 150480 300084
rect 151832 300070 152398 300098
rect 153212 300070 154330 300098
rect 155972 300070 156262 300098
rect 157352 300070 158194 300098
rect 150440 4344 150492 4350
rect 150440 4286 150492 4292
rect 151832 3126 151860 300070
rect 153212 3194 153240 300070
rect 154486 76256 154542 76265
rect 154486 76191 154542 76200
rect 154500 76158 154528 76191
rect 154488 76152 154540 76158
rect 154488 76094 154540 76100
rect 154486 40352 154542 40361
rect 154486 40287 154542 40296
rect 154500 40254 154528 40287
rect 154488 40248 154540 40254
rect 154488 40190 154540 40196
rect 154486 29336 154542 29345
rect 154486 29271 154542 29280
rect 154500 29238 154528 29271
rect 154488 29232 154540 29238
rect 154488 29174 154540 29180
rect 155972 4418 156000 300070
rect 157352 6458 157380 300070
rect 160204 297022 160232 300084
rect 161492 300070 162150 300098
rect 162872 300070 164082 300098
rect 160192 297016 160244 297022
rect 160192 296958 160244 296964
rect 157340 6452 157392 6458
rect 157340 6394 157392 6400
rect 161492 4486 161520 300070
rect 161480 4480 161532 4486
rect 161480 4422 161532 4428
rect 155960 4412 156012 4418
rect 155960 4354 156012 4360
rect 162872 3262 162900 300070
rect 166000 297090 166028 300084
rect 167012 300070 167946 300098
rect 165988 297084 166040 297090
rect 165988 297026 166040 297032
rect 167012 4554 167040 300070
rect 169864 297158 169892 300084
rect 171152 300070 171902 300098
rect 172532 300070 173834 300098
rect 175292 300070 175766 300098
rect 169852 297152 169904 297158
rect 169852 297094 169904 297100
rect 167000 4548 167052 4554
rect 167000 4490 167052 4496
rect 171152 3330 171180 300070
rect 172532 4622 172560 300070
rect 172520 4616 172572 4622
rect 172520 4558 172572 4564
rect 175292 3398 175320 300070
rect 177684 297226 177712 300084
rect 179432 300070 179630 300098
rect 177672 297220 177724 297226
rect 177672 297162 177724 297168
rect 179432 4690 179460 300070
rect 181548 297294 181576 300084
rect 181536 297288 181588 297294
rect 181536 297230 181588 297236
rect 179420 4684 179472 4690
rect 179420 4626 179472 4632
rect 183572 4146 183600 300084
rect 184952 300070 185518 300098
rect 186332 300070 187450 300098
rect 184952 4758 184980 300070
rect 184940 4752 184992 4758
rect 184940 4694 184992 4700
rect 183560 4140 183612 4146
rect 183560 4082 183612 4088
rect 186332 4078 186360 300070
rect 189368 297362 189396 300084
rect 190472 300070 191314 300098
rect 189356 297356 189408 297362
rect 189356 297298 189408 297304
rect 190472 5506 190500 300070
rect 193232 298110 193260 300084
rect 194612 300070 195178 300098
rect 195992 300070 197202 300098
rect 198752 300070 199134 300098
rect 193220 298104 193272 298110
rect 193220 298046 193272 298052
rect 190460 5500 190512 5506
rect 190460 5442 190512 5448
rect 186320 4072 186372 4078
rect 186320 4014 186372 4020
rect 194612 4010 194640 300070
rect 195992 5438 196020 300070
rect 195980 5432 196032 5438
rect 195980 5374 196032 5380
rect 194600 4004 194652 4010
rect 194600 3946 194652 3952
rect 198752 3777 198780 300070
rect 201052 298042 201080 300084
rect 202892 300070 202998 300098
rect 201040 298036 201092 298042
rect 201040 297978 201092 297984
rect 202892 5370 202920 300070
rect 204916 297974 204944 300084
rect 205652 300070 206862 300098
rect 208412 300070 208886 300098
rect 209792 300070 210818 300098
rect 204904 297968 204956 297974
rect 204904 297910 204956 297916
rect 202880 5364 202932 5370
rect 202880 5306 202932 5312
rect 205652 3942 205680 300070
rect 208412 5273 208440 300070
rect 208398 5264 208454 5273
rect 208398 5199 208454 5208
rect 205640 3936 205692 3942
rect 205640 3878 205692 3884
rect 198738 3768 198794 3777
rect 198738 3703 198794 3712
rect 209792 3641 209820 300070
rect 212736 297838 212764 300084
rect 213932 300070 214682 300098
rect 212724 297832 212776 297838
rect 212724 297774 212776 297780
rect 213932 5137 213960 300070
rect 216600 297906 216628 300084
rect 218072 300070 218546 300098
rect 219452 300070 220570 300098
rect 222212 300070 222502 300098
rect 216588 297900 216640 297906
rect 216588 297842 216640 297848
rect 213918 5128 213974 5137
rect 213918 5063 213974 5072
rect 218072 3874 218100 300070
rect 219452 5302 219480 300070
rect 219440 5296 219492 5302
rect 219440 5238 219492 5244
rect 218060 3868 218112 3874
rect 218060 3810 218112 3816
rect 209778 3632 209834 3641
rect 209778 3567 209834 3576
rect 222212 3505 222240 300070
rect 224420 297702 224448 300084
rect 224408 297696 224460 297702
rect 224408 297638 224460 297644
rect 226352 5001 226380 300084
rect 228284 297634 228312 300084
rect 229112 300070 230230 300098
rect 231872 300070 232254 300098
rect 228272 297628 228324 297634
rect 228272 297570 228324 297576
rect 226338 4992 226394 5001
rect 226338 4927 226394 4936
rect 222198 3496 222254 3505
rect 222198 3431 222254 3440
rect 175280 3392 175332 3398
rect 229112 3369 229140 300070
rect 231872 5234 231900 300070
rect 234172 297566 234200 300084
rect 234160 297560 234212 297566
rect 234160 297502 234212 297508
rect 236104 297498 236132 300084
rect 237392 300070 238050 300098
rect 238772 300070 239982 300098
rect 241532 300070 241914 300098
rect 242912 300070 243846 300098
rect 236092 297492 236144 297498
rect 236092 297434 236144 297440
rect 237392 6390 237420 300070
rect 237380 6384 237432 6390
rect 237380 6326 237432 6332
rect 231860 5228 231912 5234
rect 231860 5170 231912 5176
rect 238772 3806 238800 300070
rect 238760 3800 238812 3806
rect 238760 3742 238812 3748
rect 241532 3738 241560 300070
rect 242912 6322 242940 300070
rect 245856 297430 245884 300084
rect 247788 297673 247816 300084
rect 248432 300070 249734 300098
rect 251192 300070 251666 300098
rect 252572 300070 253598 300098
rect 247774 297664 247830 297673
rect 247774 297599 247830 297608
rect 245844 297424 245896 297430
rect 245844 297366 245896 297372
rect 242900 6316 242952 6322
rect 242900 6258 242952 6264
rect 248432 6254 248460 300070
rect 248420 6248 248472 6254
rect 248420 6190 248472 6196
rect 241520 3732 241572 3738
rect 241520 3674 241572 3680
rect 251192 3602 251220 300070
rect 252572 3670 252600 300070
rect 255516 297770 255544 300084
rect 255504 297764 255556 297770
rect 255504 297706 255556 297712
rect 257540 297537 257568 300084
rect 257526 297528 257582 297537
rect 257526 297463 257582 297472
rect 259472 297401 259500 300084
rect 260852 300070 261418 300098
rect 262232 300070 263350 300098
rect 264992 300070 265282 300098
rect 266372 300070 267214 300098
rect 269132 300070 269238 300098
rect 270512 300070 271170 300098
rect 271892 300070 273102 300098
rect 274652 300070 275034 300098
rect 276032 300070 276966 300098
rect 278792 300070 278898 300098
rect 514760 300086 514812 300092
rect 259458 297392 259514 297401
rect 259458 297327 259514 297336
rect 260852 6186 260880 300070
rect 260840 6180 260892 6186
rect 260840 6122 260892 6128
rect 252560 3664 252612 3670
rect 252560 3606 252612 3612
rect 251180 3596 251232 3602
rect 251180 3538 251232 3544
rect 262232 3534 262260 300070
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 264992 3466 265020 300070
rect 266372 5166 266400 300070
rect 266360 5160 266412 5166
rect 266360 5102 266412 5108
rect 269132 5030 269160 300070
rect 269120 5024 269172 5030
rect 269120 4966 269172 4972
rect 270512 4962 270540 300070
rect 271892 5098 271920 300070
rect 271880 5092 271932 5098
rect 271880 5034 271932 5040
rect 270500 4956 270552 4962
rect 270500 4898 270552 4904
rect 274652 4865 274680 300070
rect 276032 4894 276060 300070
rect 276020 4888 276072 4894
rect 274638 4856 274694 4865
rect 276020 4830 276072 4836
rect 278792 4826 278820 300070
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 580172 229084 580224 229090
rect 580172 229026 580224 229032
rect 580184 228857 580212 229026
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 274638 4791 274694 4800
rect 278780 4820 278832 4826
rect 278780 4762 278832 4768
rect 264980 3460 265032 3466
rect 264980 3402 265032 3408
rect 175280 3334 175332 3340
rect 229098 3360 229154 3369
rect 171140 3324 171192 3330
rect 229098 3295 229154 3304
rect 171140 3266 171192 3272
rect 162860 3256 162912 3262
rect 162860 3198 162912 3204
rect 153200 3188 153252 3194
rect 153200 3130 153252 3136
rect 151820 3120 151872 3126
rect 151820 3062 151872 3068
rect 147680 3052 147732 3058
rect 147680 2994 147732 3000
rect 139400 2984 139452 2990
rect 139400 2926 139452 2932
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 682216 2834 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3882 624824 3938 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3974 567296 4030 567352
rect 3882 553016 3938 553072
rect 2962 538600 3018 538656
rect 2778 509904 2834 509960
rect 3330 495488 3386 495544
rect 3238 481072 3294 481128
rect 3330 452396 3386 452432
rect 3330 452376 3332 452396
rect 3332 452376 3384 452396
rect 3384 452376 3386 452396
rect 2962 366152 3018 366208
rect 3330 337456 3386 337512
rect 3054 323040 3110 323096
rect 3330 308760 3386 308816
rect 2962 294344 3018 294400
rect 3330 280100 3332 280120
rect 3332 280100 3384 280120
rect 3384 280100 3386 280120
rect 3330 280064 3386 280100
rect 3146 265648 3202 265704
rect 3238 236952 3294 237008
rect 3330 222536 3386 222592
rect 3238 179424 3294 179480
rect 4066 437960 4122 438016
rect 3974 423680 4030 423736
rect 3790 394984 3846 395040
rect 3698 380568 3754 380624
rect 3606 251232 3662 251288
rect 3514 208120 3570 208176
rect 3514 193840 3570 193896
rect 3422 165008 3478 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 2778 122032 2834 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 2778 78920 2834 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 2778 35844 2780 35864
rect 2780 35844 2832 35864
rect 2832 35844 2834 35864
rect 2778 35808 2834 35844
rect 2870 21392 2926 21448
rect 3422 7112 3478 7168
rect 56598 646040 56654 646096
rect 57242 644952 57298 645008
rect 57150 643184 57206 643240
rect 57058 641960 57114 642016
rect 56966 640328 57022 640384
rect 56874 639240 56930 639296
rect 56782 637608 56838 637664
rect 56690 579672 56746 579728
rect 56598 542952 56654 543008
rect 56598 488280 56654 488336
rect 56598 486240 56654 486296
rect 56598 484064 56654 484120
rect 56598 482024 56654 482080
rect 56598 479984 56654 480040
rect 56598 477808 56654 477864
rect 56598 475768 56654 475824
rect 56598 473592 56654 473648
rect 56598 471552 56654 471608
rect 56506 469920 56562 469976
rect 56506 467780 56508 467800
rect 56508 467780 56560 467800
rect 56560 467780 56562 467800
rect 56506 467744 56562 467780
rect 56506 465704 56562 465760
rect 56506 463528 56562 463584
rect 56506 461488 56562 461544
rect 56598 458904 56654 458960
rect 56598 456748 56654 456784
rect 56598 456728 56600 456748
rect 56600 456728 56652 456748
rect 56652 456728 56654 456748
rect 56598 454688 56654 454744
rect 56598 452532 56654 452568
rect 56598 452512 56600 452532
rect 56600 452512 56652 452532
rect 56652 452512 56654 452532
rect 56598 450472 56654 450528
rect 56598 444080 56654 444136
rect 56690 433608 56746 433664
rect 56782 427216 56838 427272
rect 57242 538872 57298 538928
rect 56966 496712 57022 496768
rect 56966 490456 57022 490512
rect 56874 420960 56930 421016
rect 56598 353640 56654 353696
rect 56690 343032 56746 343088
rect 56598 309304 56654 309360
rect 56782 338816 56838 338872
rect 57058 380976 57114 381032
rect 57242 536852 57298 536888
rect 57242 536832 57244 536852
rect 57244 536832 57296 536852
rect 57296 536832 57298 536852
rect 57242 534656 57298 534712
rect 57242 532616 57298 532672
rect 57242 530440 57298 530496
rect 57242 528400 57298 528456
rect 57242 526224 57298 526280
rect 57242 524184 57298 524240
rect 57242 522008 57298 522064
rect 57242 519968 57298 520024
rect 57242 517792 57298 517848
rect 57242 515752 57298 515808
rect 57242 513576 57298 513632
rect 57242 511536 57298 511592
rect 57242 509360 57298 509416
rect 57242 507320 57298 507376
rect 57242 505164 57298 505200
rect 57242 505144 57244 505164
rect 57244 505144 57296 505164
rect 57296 505144 57298 505164
rect 57242 503104 57298 503160
rect 57242 500964 57244 500984
rect 57244 500964 57296 500984
rect 57296 500964 57298 500984
rect 57242 500928 57298 500964
rect 57242 498888 57298 498944
rect 57242 494672 57298 494728
rect 57242 492496 57298 492552
rect 57150 366152 57206 366208
rect 57058 361936 57114 361992
rect 57150 355680 57206 355736
rect 56966 336776 57022 336832
rect 56874 334600 56930 334656
rect 56782 296656 56838 296712
rect 56782 277344 56838 277400
rect 57058 332560 57114 332616
rect 57150 328344 57206 328400
rect 57518 448296 57574 448352
rect 57518 446256 57574 446312
rect 57426 439864 57482 439920
rect 57610 437824 57666 437880
rect 57334 374584 57390 374640
rect 57702 418920 57758 418976
rect 57610 368328 57666 368384
rect 57794 412528 57850 412584
rect 57886 406272 57942 406328
rect 57978 383016 58034 383072
rect 58070 376760 58126 376816
rect 58438 442040 58494 442096
rect 58530 435648 58586 435704
rect 58346 404096 58402 404152
rect 58714 431432 58770 431488
rect 58806 429392 58862 429448
rect 58898 425176 58954 425232
rect 58990 423000 59046 423056
rect 59082 416744 59138 416800
rect 59174 410488 59230 410544
rect 77206 697176 77262 697232
rect 96526 697176 96582 697232
rect 70306 697076 70308 697096
rect 70308 697076 70360 697096
rect 70360 697076 70362 697096
rect 70306 697040 70362 697076
rect 89626 697076 89628 697096
rect 89628 697076 89680 697096
rect 89680 697076 89682 697096
rect 89626 697040 89682 697076
rect 115846 697176 115902 697232
rect 135166 697176 135222 697232
rect 108946 697076 108948 697096
rect 108948 697076 109000 697096
rect 109000 697076 109002 697096
rect 108946 697040 109002 697076
rect 128266 697076 128268 697096
rect 128268 697076 128320 697096
rect 128320 697076 128322 697096
rect 128266 697040 128322 697076
rect 129278 652840 129334 652896
rect 133602 652840 133658 652896
rect 59634 578527 59690 578583
rect 67546 558864 67602 558920
rect 70122 558864 70178 558920
rect 72422 558864 72478 558920
rect 73710 558864 73766 558920
rect 75734 558864 75790 558920
rect 76010 558864 76066 558920
rect 77390 558864 77446 558920
rect 78494 558864 78550 558920
rect 64326 558728 64382 558784
rect 68926 558048 68982 558104
rect 70214 558728 70270 558784
rect 77298 558320 77354 558376
rect 73158 558184 73214 558240
rect 71594 557504 71650 557560
rect 71778 557640 71834 557696
rect 74538 557796 74594 557832
rect 74538 557776 74540 557796
rect 74540 557776 74592 557796
rect 74592 557776 74594 557796
rect 79506 558864 79562 558920
rect 80702 558864 80758 558920
rect 81438 558884 81494 558920
rect 81438 558864 81440 558884
rect 81440 558864 81492 558884
rect 81492 558864 81494 558884
rect 78678 557932 78734 557968
rect 78678 557912 78680 557932
rect 78680 557912 78732 557932
rect 78732 557912 78734 557932
rect 75918 557776 75974 557832
rect 78678 557640 78734 557696
rect 82910 558864 82966 558920
rect 84198 558864 84254 558920
rect 85394 558864 85450 558920
rect 85670 558864 85726 558920
rect 86222 558864 86278 558920
rect 80058 558728 80114 558784
rect 81622 558728 81678 558784
rect 82818 558320 82874 558376
rect 84290 558728 84346 558784
rect 87602 558864 87658 558920
rect 88982 558864 89038 558920
rect 89626 558864 89682 558920
rect 90086 558884 90142 558920
rect 90086 558864 90088 558884
rect 90088 558864 90140 558884
rect 90140 558864 90142 558884
rect 86866 558728 86922 558784
rect 87878 558764 87880 558784
rect 87880 558764 87932 558784
rect 87932 558764 87934 558784
rect 87878 558728 87934 558764
rect 91374 558864 91430 558920
rect 92478 558864 92534 558920
rect 93582 558864 93638 558920
rect 94594 558864 94650 558920
rect 95330 558864 95386 558920
rect 96618 558864 96674 558920
rect 98274 558864 98330 558920
rect 99562 558864 99618 558920
rect 100666 558864 100722 558920
rect 101954 558864 102010 558920
rect 102690 558864 102746 558920
rect 103426 558864 103482 558920
rect 103978 558864 104034 558920
rect 104806 558864 104862 558920
rect 105358 558864 105414 558920
rect 106186 558864 106242 558920
rect 107566 558864 107622 558920
rect 107842 558864 107898 558920
rect 108946 558864 109002 558920
rect 110326 558864 110382 558920
rect 100298 558748 100354 558784
rect 100298 558728 100300 558748
rect 100300 558728 100352 558748
rect 100352 558728 100354 558748
rect 93674 557640 93730 557696
rect 91006 557504 91062 557560
rect 92386 557504 92442 557560
rect 93766 557504 93822 557560
rect 95146 557504 95202 557560
rect 96526 557504 96582 557560
rect 97906 557504 97962 557560
rect 99286 557504 99342 557560
rect 101862 558592 101918 558648
rect 102046 558728 102102 558784
rect 106278 558728 106334 558784
rect 108578 558728 108634 558784
rect 154486 697176 154542 697232
rect 147586 697076 147588 697096
rect 147588 697076 147640 697096
rect 147640 697076 147642 697096
rect 147586 697040 147642 697076
rect 166906 697040 166962 697096
rect 172426 697196 172482 697232
rect 172426 697176 172428 697196
rect 172428 697176 172480 697196
rect 172480 697176 172482 697196
rect 193126 697176 193182 697232
rect 212446 697176 212502 697232
rect 231766 697176 231822 697232
rect 251086 697176 251142 697232
rect 270406 697176 270462 697232
rect 289726 697176 289782 697232
rect 186226 697076 186228 697096
rect 186228 697076 186280 697096
rect 186280 697076 186282 697096
rect 186226 697040 186282 697076
rect 205546 697076 205548 697096
rect 205548 697076 205600 697096
rect 205600 697076 205602 697096
rect 205546 697040 205602 697076
rect 224866 697076 224868 697096
rect 224868 697076 224920 697096
rect 224920 697076 224922 697096
rect 224866 697040 224922 697076
rect 244186 697076 244188 697096
rect 244188 697076 244240 697096
rect 244240 697076 244242 697096
rect 244186 697040 244242 697076
rect 263506 697076 263508 697096
rect 263508 697076 263560 697096
rect 263560 697076 263562 697096
rect 263506 697040 263562 697076
rect 282826 697076 282828 697096
rect 282828 697076 282880 697096
rect 282880 697076 282882 697096
rect 282826 697040 282882 697076
rect 166906 686296 166962 686352
rect 167090 686296 167146 686352
rect 154578 686180 154634 686216
rect 154578 686160 154580 686180
rect 154580 686160 154632 686180
rect 154632 686160 154634 686180
rect 162214 685888 162270 685944
rect 188342 686432 188398 686488
rect 173898 686316 173954 686352
rect 173898 686296 173900 686316
rect 173900 686296 173952 686316
rect 173952 686296 173954 686316
rect 178774 686160 178830 686216
rect 188342 686160 188398 686216
rect 289818 686180 289874 686216
rect 289818 686160 289820 686180
rect 289820 686160 289872 686180
rect 289872 686160 289874 686180
rect 294510 685888 294566 685944
rect 309046 697176 309102 697232
rect 328366 697176 328422 697232
rect 302146 697076 302148 697096
rect 302148 697076 302200 697096
rect 302200 697076 302202 697096
rect 302146 697040 302202 697076
rect 321466 697076 321468 697096
rect 321468 697076 321520 697096
rect 321520 697076 321522 697096
rect 321466 697040 321522 697076
rect 360106 686296 360162 686352
rect 360290 686296 360346 686352
rect 347778 686180 347834 686216
rect 347778 686160 347780 686180
rect 347780 686160 347832 686180
rect 347832 686160 347834 686180
rect 355414 685888 355470 685944
rect 166998 673920 167054 673976
rect 154578 673804 154634 673840
rect 154578 673784 154580 673804
rect 154580 673784 154632 673804
rect 154632 673784 154634 673804
rect 162214 673512 162270 673568
rect 166906 673512 166962 673568
rect 188342 674056 188398 674112
rect 173898 673940 173954 673976
rect 173898 673920 173900 673940
rect 173900 673920 173952 673940
rect 173952 673920 173954 673940
rect 178774 673784 178830 673840
rect 188342 673784 188398 673840
rect 289818 673804 289874 673840
rect 289818 673784 289820 673804
rect 289820 673784 289872 673804
rect 289872 673784 289874 673804
rect 292670 673512 292726 673568
rect 169850 666576 169906 666632
rect 170034 666576 170090 666632
rect 360106 673920 360162 673976
rect 360290 673920 360346 673976
rect 347778 673804 347834 673840
rect 347778 673784 347780 673804
rect 347780 673784 347832 673804
rect 347832 673784 347834 673804
rect 355414 673512 355470 673568
rect 379518 686432 379574 686488
rect 367098 686316 367154 686352
rect 367098 686296 367100 686316
rect 367100 686296 367152 686316
rect 367152 686296 367154 686316
rect 371974 686160 372030 686216
rect 379518 686160 379574 686216
rect 427542 686160 427598 686216
rect 427726 686160 427782 686216
rect 441526 686432 441582 686488
rect 441526 686160 441582 686216
rect 379518 674056 379574 674112
rect 367098 673940 367154 673976
rect 367098 673920 367100 673940
rect 367100 673920 367152 673940
rect 367152 673920 367154 673940
rect 371974 673784 372030 673840
rect 379518 673784 379574 673840
rect 139398 649848 139454 649904
rect 259182 652840 259238 652896
rect 263782 652840 263838 652896
rect 266450 649848 266506 649904
rect 187698 646176 187754 646232
rect 169758 645904 169814 645960
rect 170034 645904 170090 645960
rect 139398 589600 139454 589656
rect 158534 542952 158590 543008
rect 187698 644816 187754 644872
rect 187698 643184 187754 643240
rect 187698 641960 187754 642016
rect 187698 640348 187754 640384
rect 187698 640328 187700 640348
rect 187700 640328 187752 640348
rect 187752 640328 187754 640348
rect 188342 639240 188398 639296
rect 170034 587832 170090 587888
rect 170310 587832 170366 587888
rect 187698 579692 187754 579728
rect 187698 579672 187700 579692
rect 187700 579672 187752 579692
rect 187752 579672 187754 579692
rect 188434 637608 188490 637664
rect 269118 589328 269174 589384
rect 269118 587696 269174 587752
rect 270038 580896 270094 580952
rect 188986 578312 189042 578368
rect 211066 559952 211122 560008
rect 210422 559816 210478 559872
rect 193770 558864 193826 558920
rect 202786 558864 202842 558920
rect 204166 558864 204222 558920
rect 205546 558864 205602 558920
rect 195978 558728 196034 558784
rect 201498 558728 201554 558784
rect 202142 558728 202198 558784
rect 197358 558592 197414 558648
rect 198738 558456 198794 558512
rect 200210 558456 200266 558512
rect 203522 558592 203578 558648
rect 204902 558728 204958 558784
rect 209042 558592 209098 558648
rect 206282 558068 206338 558104
rect 206282 558048 206284 558068
rect 206284 558048 206336 558068
rect 206336 558048 206338 558068
rect 207662 557676 207664 557696
rect 207664 557676 207716 557696
rect 207716 557676 207718 557696
rect 206926 557504 206982 557560
rect 207662 557640 207718 557676
rect 209226 557640 209282 557696
rect 208306 557504 208362 557560
rect 209686 557504 209742 557560
rect 210974 557640 211030 557696
rect 211894 558864 211950 558920
rect 213182 558864 213238 558920
rect 213918 558864 213974 558920
rect 216586 558864 216642 558920
rect 217598 558864 217654 558920
rect 217874 558864 217930 558920
rect 218886 558864 218942 558920
rect 219346 558864 219402 558920
rect 220082 558864 220138 558920
rect 220726 558864 220782 558920
rect 221094 558864 221150 558920
rect 222106 558864 222162 558920
rect 222290 558864 222346 558920
rect 223486 558864 223542 558920
rect 224866 558864 224922 558920
rect 225786 558864 225842 558920
rect 226246 558864 226302 558920
rect 227166 558864 227222 558920
rect 227626 558864 227682 558920
rect 229006 558864 229062 558920
rect 229466 558864 229522 558920
rect 230386 558864 230442 558920
rect 231766 558864 231822 558920
rect 231950 558864 232006 558920
rect 233146 558864 233202 558920
rect 234526 558864 234582 558920
rect 235906 558864 235962 558920
rect 237286 558864 237342 558920
rect 240046 558864 240102 558920
rect 215298 558728 215354 558784
rect 212446 557504 212502 557560
rect 213826 557504 213882 557560
rect 215206 557504 215262 557560
rect 211250 550568 211306 550624
rect 211434 550568 211490 550624
rect 216770 558748 216826 558784
rect 216770 558728 216772 558748
rect 216772 558728 216824 558748
rect 216824 558728 216826 558748
rect 217966 558728 218022 558784
rect 223578 558764 223580 558784
rect 223580 558764 223632 558784
rect 223632 558764 223634 558784
rect 223578 558728 223634 558764
rect 224406 558728 224462 558784
rect 226154 558728 226210 558784
rect 227718 558728 227774 558784
rect 230478 558592 230534 558648
rect 233054 558728 233110 558784
rect 231858 558612 231914 558648
rect 231858 558592 231860 558612
rect 231860 558592 231912 558612
rect 231912 558592 231914 558612
rect 233238 558728 233294 558784
rect 234618 558592 234674 558648
rect 235998 558748 236054 558784
rect 235998 558728 236000 558748
rect 236000 558728 236052 558748
rect 236052 558728 236054 558748
rect 237378 558456 237434 558512
rect 238758 558456 238814 558512
rect 238666 558048 238722 558104
rect 59542 414704 59598 414760
rect 59450 402056 59506 402112
rect 59358 399880 59414 399936
rect 59266 397840 59322 397896
rect 59726 408312 59782 408368
rect 59634 395664 59690 395720
rect 58622 385192 58678 385248
rect 58254 372544 58310 372600
rect 58162 370368 58218 370424
rect 57702 364112 57758 364168
rect 57702 359896 57758 359952
rect 57426 357856 57482 357912
rect 57334 349424 57390 349480
rect 57334 330384 57390 330440
rect 57518 351464 57574 351520
rect 57426 326168 57482 326224
rect 57334 315968 57390 316024
rect 57334 306448 57390 306504
rect 57334 277344 57390 277400
rect 57610 345208 57666 345264
rect 57794 347248 57850 347304
rect 57702 324128 57758 324184
rect 57886 340992 57942 341048
rect 57794 321952 57850 322008
rect 57794 317736 57850 317792
rect 57702 315696 57758 315752
rect 57610 296656 57666 296712
rect 59082 313520 59138 313576
rect 59174 307264 59230 307320
rect 59358 319912 59414 319968
rect 59266 301008 59322 301064
rect 378506 652840 378562 652896
rect 383474 652840 383530 652896
rect 281538 303320 281594 303376
rect 281722 538872 281778 538928
rect 282826 536732 282828 536752
rect 282828 536732 282880 536752
rect 282880 536732 282882 536752
rect 282826 536696 282882 536732
rect 282826 534520 282882 534576
rect 282826 532344 282882 532400
rect 282826 530168 282882 530224
rect 282826 527856 282882 527912
rect 282826 525716 282828 525736
rect 282828 525716 282880 525736
rect 282880 525716 282882 525736
rect 282826 525680 282882 525716
rect 282826 523504 282882 523560
rect 282826 521328 282882 521384
rect 282826 519152 282882 519208
rect 281906 516840 281962 516896
rect 282826 514700 282828 514720
rect 282828 514700 282880 514720
rect 282880 514700 282882 514720
rect 282826 514664 282882 514700
rect 282090 512488 282146 512544
rect 282826 510312 282882 510368
rect 282274 508136 282330 508192
rect 281906 505824 281962 505880
rect 282826 503668 282882 503704
rect 282826 503648 282828 503668
rect 282828 503648 282880 503668
rect 282880 503648 282882 503668
rect 282090 501472 282146 501528
rect 282826 499296 282882 499352
rect 282274 497120 282330 497176
rect 281906 494808 281962 494864
rect 282458 492632 282514 492688
rect 282090 490456 282146 490512
rect 282826 488280 282882 488336
rect 282826 486104 282882 486160
rect 282826 483792 282882 483848
rect 282458 481616 282514 481672
rect 282090 479440 282146 479496
rect 282826 477264 282882 477320
rect 282550 475088 282606 475144
rect 282090 472912 282146 472968
rect 282458 470600 282514 470656
rect 282090 468424 282146 468480
rect 282826 466248 282882 466304
rect 282274 464072 282330 464128
rect 282826 461896 282882 461952
rect 282458 459584 282514 459640
rect 282090 457408 282146 457464
rect 282826 455232 282882 455288
rect 282826 453056 282882 453112
rect 282826 450880 282882 450936
rect 282458 448568 282514 448624
rect 282826 446392 282882 446448
rect 282826 444216 282882 444272
rect 282826 442040 282882 442096
rect 282826 439864 282882 439920
rect 282458 437552 282514 437608
rect 282826 435376 282882 435432
rect 282826 433236 282828 433256
rect 282828 433236 282880 433256
rect 282880 433236 282882 433256
rect 282826 433200 282882 433236
rect 282826 431024 282882 431080
rect 282826 428848 282882 428904
rect 282826 426572 282828 426592
rect 282828 426572 282880 426592
rect 282880 426572 282882 426592
rect 282826 426536 282882 426572
rect 282458 424360 282514 424416
rect 282090 422220 282092 422240
rect 282092 422220 282144 422240
rect 282144 422220 282146 422240
rect 282090 422184 282146 422220
rect 281722 420008 281778 420064
rect 282826 417832 282882 417888
rect 282826 415656 282882 415712
rect 281906 413344 281962 413400
rect 282826 411204 282828 411224
rect 282828 411204 282880 411224
rect 282880 411204 282882 411224
rect 282826 411168 282882 411204
rect 282090 408992 282146 409048
rect 282826 406816 282882 406872
rect 282826 404640 282882 404696
rect 281906 402328 281962 402384
rect 282826 400172 282882 400208
rect 282826 400152 282828 400172
rect 282828 400152 282880 400172
rect 282880 400152 282882 400172
rect 282090 397976 282146 398032
rect 282090 395836 282092 395856
rect 282092 395836 282144 395856
rect 282144 395836 282146 395856
rect 282090 395800 282146 395836
rect 282274 393624 282330 393680
rect 281906 391312 281962 391368
rect 282458 389136 282514 389192
rect 282090 386960 282146 387016
rect 282826 384784 282882 384840
rect 282826 382608 282882 382664
rect 282826 380296 282882 380352
rect 282458 378120 282514 378176
rect 282090 375944 282146 376000
rect 282826 373768 282882 373824
rect 282550 371592 282606 371648
rect 282826 369280 282882 369336
rect 282458 367104 282514 367160
rect 282090 364928 282146 364984
rect 282826 362752 282882 362808
rect 282550 360576 282606 360632
rect 282826 358400 282882 358456
rect 282458 356088 282514 356144
rect 282090 353912 282146 353968
rect 282826 351736 282882 351792
rect 282550 349560 282606 349616
rect 282826 347384 282882 347440
rect 282458 345072 282514 345128
rect 282826 342896 282882 342952
rect 282826 340720 282882 340776
rect 282826 338544 282882 338600
rect 282826 336368 282882 336424
rect 282366 334056 282422 334112
rect 282826 331880 282882 331936
rect 282826 329740 282828 329760
rect 282828 329740 282880 329760
rect 282880 329740 282882 329760
rect 282826 329704 282882 329740
rect 282826 327528 282882 327584
rect 282826 325352 282882 325408
rect 282366 323040 282422 323096
rect 282826 320864 282882 320920
rect 389178 649848 389234 649904
rect 553306 697312 553362 697368
rect 553490 697312 553546 697368
rect 540978 697196 541034 697232
rect 540978 697176 540980 697196
rect 540980 697176 541032 697196
rect 541032 697176 541034 697196
rect 548614 696904 548670 696960
rect 553306 686296 553362 686352
rect 553490 686296 553546 686352
rect 540978 686180 541034 686216
rect 540978 686160 540980 686180
rect 540980 686160 541032 686180
rect 541032 686160 541034 686180
rect 548614 685888 548670 685944
rect 560298 697332 560354 697368
rect 560298 697312 560300 697332
rect 560300 697312 560352 697332
rect 560352 697312 560354 697332
rect 565174 697176 565230 697232
rect 572718 697176 572774 697232
rect 572626 697040 572682 697096
rect 560298 686316 560354 686352
rect 560298 686296 560300 686316
rect 560300 686296 560352 686316
rect 560352 686296 560354 686316
rect 565174 686160 565230 686216
rect 572718 686160 572774 686216
rect 572626 686024 572682 686080
rect 559010 684392 559066 684448
rect 559010 684256 559066 684312
rect 553398 673920 553454 673976
rect 540978 673804 541034 673840
rect 540978 673784 540980 673804
rect 540980 673784 541032 673804
rect 541032 673784 541034 673804
rect 548614 673512 548670 673568
rect 553306 673512 553362 673568
rect 560298 673940 560354 673976
rect 560298 673920 560300 673940
rect 560300 673920 560352 673940
rect 560352 673920 560354 673940
rect 565174 673784 565230 673840
rect 572718 673784 572774 673840
rect 572626 673648 572682 673704
rect 507858 652840 507914 652896
rect 513378 652860 513434 652896
rect 513378 652840 513380 652860
rect 513380 652840 513432 652860
rect 513432 652840 513434 652860
rect 307390 646040 307446 646096
rect 307114 644952 307170 645008
rect 307114 643456 307170 643512
rect 307666 642096 307722 642152
rect 307666 640464 307722 640520
rect 306654 639376 306710 639432
rect 299570 637880 299626 637936
rect 299662 637472 299718 637528
rect 300030 637472 300086 637528
rect 306930 579944 306986 580000
rect 306378 578312 306434 578368
rect 347962 559272 348018 559328
rect 357714 559272 357770 559328
rect 313738 558864 313794 558920
rect 316038 558864 316094 558920
rect 318798 558864 318854 558920
rect 320270 558864 320326 558920
rect 321558 558864 321614 558920
rect 323582 558864 323638 558920
rect 325698 558864 325754 558920
rect 327078 558864 327134 558920
rect 329930 558864 329986 558920
rect 331770 558864 331826 558920
rect 332598 558864 332654 558920
rect 333978 558864 334034 558920
rect 335358 558864 335414 558920
rect 282826 318724 282828 318744
rect 282828 318724 282880 318744
rect 282880 318724 282882 318744
rect 282826 318688 282882 318724
rect 282826 316512 282882 316568
rect 282826 314336 282882 314392
rect 282366 312024 282422 312080
rect 281906 309848 281962 309904
rect 317418 558456 317474 558512
rect 320178 557776 320234 557832
rect 282826 307708 282828 307728
rect 282828 307708 282880 307728
rect 282880 307708 282882 307728
rect 282826 307672 282882 307708
rect 322294 558728 322350 558784
rect 322938 557912 322994 557968
rect 323674 558592 323730 558648
rect 324962 558592 325018 558648
rect 326342 558592 326398 558648
rect 327722 558728 327778 558784
rect 329102 558728 329158 558784
rect 328458 558184 328514 558240
rect 329286 558592 329342 558648
rect 329838 558320 329894 558376
rect 330482 558592 330538 558648
rect 331218 558184 331274 558240
rect 332690 558728 332746 558784
rect 334070 558728 334126 558784
rect 336738 558864 336794 558920
rect 337382 558864 337438 558920
rect 338118 558864 338174 558920
rect 339498 558864 339554 558920
rect 340878 558864 340934 558920
rect 342258 558864 342314 558920
rect 343638 558864 343694 558920
rect 344282 558884 344338 558920
rect 344282 558864 344284 558884
rect 344284 558864 344336 558884
rect 344336 558864 344338 558884
rect 335450 558728 335506 558784
rect 336646 558728 336702 558784
rect 336830 558456 336886 558512
rect 338946 558728 339002 558784
rect 339866 558728 339922 558784
rect 340970 558728 341026 558784
rect 342534 558728 342590 558784
rect 345018 558864 345074 558920
rect 346398 558864 346454 558920
rect 347778 558864 347834 558920
rect 343730 558764 343732 558784
rect 343732 558764 343784 558784
rect 343784 558764 343786 558784
rect 343730 558728 343786 558764
rect 343730 557640 343786 557696
rect 346306 558728 346362 558784
rect 346950 558728 347006 558784
rect 349158 558864 349214 558920
rect 351918 558864 351974 558920
rect 348330 558728 348386 558784
rect 349526 558728 349582 558784
rect 353298 558748 353354 558784
rect 353298 558728 353300 558748
rect 353300 558728 353352 558748
rect 353352 558728 353354 558748
rect 350538 558476 350594 558512
rect 350538 558456 350540 558476
rect 350540 558456 350592 558476
rect 350592 558456 350594 558476
rect 354678 558320 354734 558376
rect 352010 557640 352066 557696
rect 350538 557504 350594 557560
rect 352194 555464 352250 555520
rect 353298 557504 353354 557560
rect 354770 557504 354826 557560
rect 357438 558728 357494 558784
rect 356058 558612 356114 558648
rect 356058 558592 356060 558612
rect 356060 558592 356112 558612
rect 356112 558592 356114 558612
rect 356058 557504 356114 557560
rect 357438 557504 357494 557560
rect 358818 555464 358874 555520
rect 389178 589600 389234 589656
rect 516414 649848 516470 649904
rect 437478 646176 437534 646232
rect 437478 644816 437534 644872
rect 437478 643184 437534 643240
rect 437478 641960 437534 642016
rect 437478 640348 437534 640384
rect 437478 640328 437480 640348
rect 437480 640328 437532 640348
rect 437532 640328 437534 640348
rect 437478 639240 437534 639296
rect 437478 637628 437534 637664
rect 437478 637608 437480 637628
rect 437480 637608 437532 637628
rect 437532 637608 437534 637628
rect 580170 651072 580226 651128
rect 580262 639376 580318 639432
rect 518898 589328 518954 589384
rect 518898 587696 518954 587752
rect 437478 579692 437534 579728
rect 437478 579672 437480 579692
rect 437480 579672 437532 579692
rect 437532 579672 437534 579692
rect 438122 578312 438178 578368
rect 443090 558864 443146 558920
rect 445758 558864 445814 558920
rect 446402 558864 446458 558920
rect 447782 558864 447838 558920
rect 449162 558864 449218 558920
rect 452750 558864 452806 558920
rect 453486 558864 453542 558920
rect 454682 558864 454738 558920
rect 458822 558864 458878 558920
rect 460938 558864 460994 558920
rect 461766 558864 461822 558920
rect 462318 558864 462374 558920
rect 463698 558864 463754 558920
rect 465078 558864 465134 558920
rect 466458 558864 466514 558920
rect 467838 558864 467894 558920
rect 468574 558864 468630 558920
rect 469218 558864 469274 558920
rect 470598 558864 470654 558920
rect 471978 558864 472034 558920
rect 473358 558864 473414 558920
rect 474738 558864 474794 558920
rect 476210 558864 476266 558920
rect 477130 558864 477186 558920
rect 478326 558864 478382 558920
rect 479430 558864 479486 558920
rect 480534 558864 480590 558920
rect 483018 558884 483074 558920
rect 483018 558864 483020 558884
rect 483020 558864 483072 558884
rect 483072 558864 483074 558884
rect 452658 558184 452714 558240
rect 451370 557640 451426 557696
rect 453302 558728 453358 558784
rect 454038 558320 454094 558376
rect 456062 558592 456118 558648
rect 457442 558592 457498 558648
rect 455418 558456 455474 558512
rect 456798 558340 456854 558376
rect 456798 558320 456800 558340
rect 456800 558320 456852 558340
rect 456852 558320 456854 558340
rect 458178 558320 458234 558376
rect 460202 558728 460258 558784
rect 460662 558748 460718 558784
rect 460662 558728 460664 558748
rect 460664 558728 460716 558748
rect 460716 558728 460718 558748
rect 459558 558204 459614 558240
rect 459558 558184 459560 558204
rect 459560 558184 459612 558204
rect 459612 558184 459614 558204
rect 460846 558592 460902 558648
rect 461030 558728 461086 558784
rect 462962 558728 463018 558784
rect 464342 558728 464398 558784
rect 465170 558728 465226 558784
rect 466550 558592 466606 558648
rect 467930 558728 467986 558784
rect 468022 558592 468078 558648
rect 470046 558728 470102 558784
rect 471242 558728 471298 558784
rect 472254 558728 472310 558784
rect 473542 558728 473598 558784
rect 474646 557640 474702 557696
rect 474830 558728 474886 558784
rect 475566 558748 475622 558784
rect 475566 558728 475568 558748
rect 475568 558728 475620 558748
rect 475620 558728 475622 558748
rect 476118 558068 476174 558104
rect 476118 558048 476120 558068
rect 476120 558048 476172 558068
rect 476172 558048 476174 558068
rect 480442 558728 480498 558784
rect 477498 558048 477554 558104
rect 478878 557932 478934 557968
rect 478878 557912 478880 557932
rect 478880 557912 478932 557932
rect 478932 557912 478934 557932
rect 484490 558864 484546 558920
rect 485778 558864 485834 558920
rect 484398 558748 484454 558784
rect 484398 558728 484400 558748
rect 484400 558728 484452 558748
rect 484452 558728 484454 558748
rect 483018 558612 483074 558648
rect 483018 558592 483020 558612
rect 483020 558592 483072 558612
rect 483072 558592 483074 558612
rect 488538 558592 488594 558648
rect 481638 558456 481694 558512
rect 487158 558456 487214 558512
rect 488538 558320 488594 558376
rect 483018 558184 483074 558240
rect 485778 558184 485834 558240
rect 487158 558204 487214 558240
rect 487158 558184 487160 558204
rect 487160 558184 487212 558204
rect 487212 558184 487214 558204
rect 481638 557776 481694 557832
rect 483018 557640 483074 557696
rect 579618 557232 579674 557288
rect 580170 545536 580226 545592
rect 580354 627680 580410 627736
rect 580262 539144 580318 539200
rect 580446 604152 580502 604208
rect 580538 592456 580594 592512
rect 580446 539008 580502 539064
rect 580630 580760 580686 580816
rect 579802 533840 579858 533896
rect 580262 510312 580318 510368
rect 580262 498616 580318 498672
rect 578882 486784 578938 486840
rect 579986 463392 580042 463448
rect 580262 451696 580318 451752
rect 579618 439864 579674 439920
rect 580262 416472 580318 416528
rect 580906 404776 580962 404832
rect 282090 305496 282146 305552
rect 281630 301144 281686 301200
rect 60830 300600 60886 300656
rect 579618 392944 579674 393000
rect 579526 369552 579582 369608
rect 579526 357856 579582 357912
rect 580170 346024 580226 346080
rect 580262 322632 580318 322688
rect 580354 310800 580410 310856
rect 61106 299512 61162 299568
rect 60922 173848 60978 173904
rect 61106 173848 61162 173904
rect 60922 143520 60978 143576
rect 61198 143520 61254 143576
rect 60738 106256 60794 106312
rect 61014 106256 61070 106312
rect 67362 240080 67418 240136
rect 67546 240080 67602 240136
rect 67546 177248 67602 177304
rect 67546 164192 67602 164248
rect 67546 125976 67602 126032
rect 67546 125568 67602 125624
rect 67454 37168 67510 37224
rect 67730 37168 67786 37224
rect 68650 3440 68706 3496
rect 77206 76200 77262 76256
rect 77206 75792 77262 75848
rect 77206 40296 77262 40352
rect 77206 39888 77262 39944
rect 74630 3576 74686 3632
rect 78954 4004 79010 4040
rect 78954 3984 78956 4004
rect 78956 3984 79008 4004
rect 79008 3984 79010 4004
rect 83002 3984 83058 4040
rect 86038 3984 86094 4040
rect 89534 76100 89536 76120
rect 89536 76100 89588 76120
rect 89588 76100 89590 76120
rect 89534 76064 89590 76100
rect 89534 40180 89590 40216
rect 89534 40160 89536 40180
rect 89536 40160 89588 40180
rect 89588 40160 89590 40180
rect 84934 3712 84990 3768
rect 84014 3576 84070 3632
rect 84106 3460 84162 3496
rect 84106 3440 84108 3460
rect 84108 3440 84160 3460
rect 84160 3440 84162 3460
rect 89810 76100 89812 76120
rect 89812 76100 89864 76120
rect 89864 76100 89866 76120
rect 89810 76064 89866 76100
rect 91742 40180 91798 40216
rect 91742 40160 91744 40180
rect 91744 40160 91796 40180
rect 91796 40160 91798 40180
rect 91742 29552 91798 29608
rect 91742 29144 91798 29200
rect 90914 5208 90970 5264
rect 89718 3984 89774 4040
rect 94502 5072 94558 5128
rect 93214 3884 93216 3904
rect 93216 3884 93268 3904
rect 93268 3884 93270 3904
rect 93214 3848 93270 3884
rect 93858 3884 93860 3904
rect 93860 3884 93912 3904
rect 93912 3884 93914 3904
rect 92110 3576 92166 3632
rect 93858 3848 93914 3884
rect 93858 3304 93914 3360
rect 93950 3168 94006 3224
rect 95514 3868 95570 3904
rect 95514 3848 95516 3868
rect 95516 3848 95568 3868
rect 95568 3848 95570 3868
rect 96618 3848 96674 3904
rect 99286 3440 99342 3496
rect 99378 3304 99434 3360
rect 99470 3168 99526 3224
rect 101586 4936 101642 4992
rect 102690 3848 102746 3904
rect 104898 3848 104954 3904
rect 103978 3304 104034 3360
rect 109866 3848 109922 3904
rect 115846 297608 115902 297664
rect 115938 75964 115940 75984
rect 115940 75964 115992 75984
rect 115992 75964 115994 75984
rect 115938 75928 115994 75964
rect 115938 40060 115940 40080
rect 115940 40060 115992 40080
rect 115992 40060 115994 40080
rect 115938 40024 115994 40060
rect 115938 29044 115940 29064
rect 115940 29044 115992 29064
rect 115992 29044 115994 29064
rect 115938 29008 115994 29044
rect 117318 3848 117374 3904
rect 118882 76200 118938 76256
rect 118882 40296 118938 40352
rect 121366 297472 121422 297528
rect 120814 29280 120870 29336
rect 122746 297336 122802 297392
rect 128266 29280 128322 29336
rect 128450 29144 128506 29200
rect 131394 4800 131450 4856
rect 135166 76472 135222 76528
rect 135166 76064 135222 76120
rect 135166 40568 135222 40624
rect 135166 40160 135222 40216
rect 140042 76336 140098 76392
rect 140042 75928 140098 75984
rect 140042 40432 140098 40488
rect 140042 40024 140098 40080
rect 143446 29416 143502 29472
rect 143446 29008 143502 29064
rect 147586 76100 147588 76120
rect 147588 76100 147640 76120
rect 147640 76100 147642 76120
rect 147586 76064 147642 76100
rect 147586 40196 147588 40216
rect 147588 40196 147640 40216
rect 147640 40196 147642 40216
rect 147586 40160 147642 40196
rect 147586 29180 147588 29200
rect 147588 29180 147640 29200
rect 147640 29180 147642 29200
rect 147586 29144 147642 29180
rect 154486 76200 154542 76256
rect 154486 40296 154542 40352
rect 154486 29280 154542 29336
rect 208398 5208 208454 5264
rect 198738 3712 198794 3768
rect 213918 5072 213974 5128
rect 209778 3576 209834 3632
rect 226338 4936 226394 4992
rect 222198 3440 222254 3496
rect 247774 297608 247830 297664
rect 257526 297472 257582 297528
rect 259458 297336 259514 297392
rect 274638 4800 274694 4856
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 580170 228792 580226 228848
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 579802 64504 579858 64560
rect 579802 17584 579858 17640
rect 229098 3304 229154 3360
<< metal3 >>
rect 583520 698050 584960 698140
rect 583342 697990 584960 698050
rect 550582 697308 550588 697372
rect 550652 697370 550658 697372
rect 553301 697370 553367 697373
rect 550652 697368 553367 697370
rect 550652 697312 553306 697368
rect 553362 697312 553367 697368
rect 550652 697310 553367 697312
rect 550652 697308 550658 697310
rect 553301 697307 553367 697310
rect 553485 697370 553551 697373
rect 560293 697370 560359 697373
rect 553485 697368 560359 697370
rect 553485 697312 553490 697368
rect 553546 697312 560298 697368
rect 560354 697312 560359 697368
rect 553485 697310 560359 697312
rect 553485 697307 553551 697310
rect 560293 697307 560359 697310
rect 59118 697172 59124 697236
rect 59188 697234 59194 697236
rect 77201 697234 77267 697237
rect 96521 697234 96587 697237
rect 115841 697234 115907 697237
rect 135161 697234 135227 697237
rect 154481 697234 154547 697237
rect 172421 697234 172487 697237
rect 193121 697234 193187 697237
rect 212441 697234 212507 697237
rect 231761 697234 231827 697237
rect 251081 697234 251147 697237
rect 270401 697234 270467 697237
rect 289721 697234 289787 697237
rect 309041 697234 309107 697237
rect 328361 697234 328427 697237
rect 540973 697234 541039 697237
rect 59188 697174 60842 697234
rect 59188 697172 59194 697174
rect 60782 697098 60842 697174
rect 77201 697232 80162 697234
rect 77201 697176 77206 697232
rect 77262 697176 80162 697232
rect 77201 697174 80162 697176
rect 77201 697171 77267 697174
rect 70301 697098 70367 697101
rect 60782 697096 70367 697098
rect 60782 697040 70306 697096
rect 70362 697040 70367 697096
rect 60782 697038 70367 697040
rect 80102 697098 80162 697174
rect 96521 697232 99482 697234
rect 96521 697176 96526 697232
rect 96582 697176 99482 697232
rect 96521 697174 99482 697176
rect 96521 697171 96587 697174
rect 89621 697098 89687 697101
rect 80102 697096 89687 697098
rect 80102 697040 89626 697096
rect 89682 697040 89687 697096
rect 80102 697038 89687 697040
rect 99422 697098 99482 697174
rect 115841 697232 118802 697234
rect 115841 697176 115846 697232
rect 115902 697176 118802 697232
rect 115841 697174 118802 697176
rect 115841 697171 115907 697174
rect 108941 697098 109007 697101
rect 99422 697096 109007 697098
rect 99422 697040 108946 697096
rect 109002 697040 109007 697096
rect 99422 697038 109007 697040
rect 118742 697098 118802 697174
rect 135161 697232 138122 697234
rect 135161 697176 135166 697232
rect 135222 697176 138122 697232
rect 135161 697174 138122 697176
rect 135161 697171 135227 697174
rect 128261 697098 128327 697101
rect 118742 697096 128327 697098
rect 118742 697040 128266 697096
rect 128322 697040 128327 697096
rect 118742 697038 128327 697040
rect 138062 697098 138122 697174
rect 154481 697232 157442 697234
rect 154481 697176 154486 697232
rect 154542 697176 157442 697232
rect 154481 697174 157442 697176
rect 154481 697171 154547 697174
rect 147581 697098 147647 697101
rect 138062 697096 147647 697098
rect 138062 697040 147586 697096
rect 147642 697040 147647 697096
rect 138062 697038 147647 697040
rect 157382 697098 157442 697174
rect 172421 697232 176762 697234
rect 172421 697176 172426 697232
rect 172482 697176 176762 697232
rect 172421 697174 176762 697176
rect 172421 697171 172487 697174
rect 166901 697098 166967 697101
rect 157382 697096 166967 697098
rect 157382 697040 166906 697096
rect 166962 697040 166967 697096
rect 157382 697038 166967 697040
rect 176702 697098 176762 697174
rect 193121 697232 196082 697234
rect 193121 697176 193126 697232
rect 193182 697176 196082 697232
rect 193121 697174 196082 697176
rect 193121 697171 193187 697174
rect 186221 697098 186287 697101
rect 176702 697096 186287 697098
rect 176702 697040 186226 697096
rect 186282 697040 186287 697096
rect 176702 697038 186287 697040
rect 196022 697098 196082 697174
rect 212441 697232 215402 697234
rect 212441 697176 212446 697232
rect 212502 697176 215402 697232
rect 212441 697174 215402 697176
rect 212441 697171 212507 697174
rect 205541 697098 205607 697101
rect 196022 697096 205607 697098
rect 196022 697040 205546 697096
rect 205602 697040 205607 697096
rect 196022 697038 205607 697040
rect 215342 697098 215402 697174
rect 231761 697232 234722 697234
rect 231761 697176 231766 697232
rect 231822 697176 234722 697232
rect 231761 697174 234722 697176
rect 231761 697171 231827 697174
rect 224861 697098 224927 697101
rect 215342 697096 224927 697098
rect 215342 697040 224866 697096
rect 224922 697040 224927 697096
rect 215342 697038 224927 697040
rect 234662 697098 234722 697174
rect 251081 697232 254042 697234
rect 251081 697176 251086 697232
rect 251142 697176 254042 697232
rect 251081 697174 254042 697176
rect 251081 697171 251147 697174
rect 244181 697098 244247 697101
rect 234662 697096 244247 697098
rect 234662 697040 244186 697096
rect 244242 697040 244247 697096
rect 234662 697038 244247 697040
rect 253982 697098 254042 697174
rect 270401 697232 273362 697234
rect 270401 697176 270406 697232
rect 270462 697176 273362 697232
rect 270401 697174 273362 697176
rect 270401 697171 270467 697174
rect 263501 697098 263567 697101
rect 253982 697096 263567 697098
rect 253982 697040 263506 697096
rect 263562 697040 263567 697096
rect 253982 697038 263567 697040
rect 273302 697098 273362 697174
rect 289721 697232 292682 697234
rect 289721 697176 289726 697232
rect 289782 697176 292682 697232
rect 289721 697174 292682 697176
rect 289721 697171 289787 697174
rect 282821 697098 282887 697101
rect 273302 697096 282887 697098
rect 273302 697040 282826 697096
rect 282882 697040 282887 697096
rect 273302 697038 282887 697040
rect 292622 697098 292682 697174
rect 309041 697232 312002 697234
rect 309041 697176 309046 697232
rect 309102 697176 312002 697232
rect 309041 697174 312002 697176
rect 309041 697171 309107 697174
rect 302141 697098 302207 697101
rect 292622 697096 302207 697098
rect 292622 697040 302146 697096
rect 302202 697040 302207 697096
rect 292622 697038 302207 697040
rect 311942 697098 312002 697174
rect 328361 697232 340890 697234
rect 328361 697176 328366 697232
rect 328422 697176 340890 697232
rect 328361 697174 340890 697176
rect 328361 697171 328427 697174
rect 321461 697098 321527 697101
rect 311942 697096 321527 697098
rect 311942 697040 321466 697096
rect 321522 697040 321527 697096
rect 311942 697038 321527 697040
rect 340830 697098 340890 697174
rect 373950 697174 383578 697234
rect 340830 697038 350458 697098
rect 70301 697035 70367 697038
rect 89621 697035 89687 697038
rect 108941 697035 109007 697038
rect 128261 697035 128327 697038
rect 147581 697035 147647 697038
rect 166901 697035 166967 697038
rect 186221 697035 186287 697038
rect 205541 697035 205607 697038
rect 224861 697035 224927 697038
rect 244181 697035 244247 697038
rect 263501 697035 263567 697038
rect 282821 697035 282887 697038
rect 302141 697035 302207 697038
rect 321461 697035 321527 697038
rect 350398 696962 350458 697038
rect 373950 696962 374010 697174
rect 350398 696902 374010 696962
rect 383518 696962 383578 697174
rect 383702 697174 393330 697234
rect 383702 696962 383762 697174
rect 393270 697098 393330 697174
rect 403022 697174 412650 697234
rect 393270 697038 402898 697098
rect 383518 696902 383762 696962
rect 402838 696962 402898 697038
rect 403022 696962 403082 697174
rect 412590 697098 412650 697174
rect 422342 697174 431970 697234
rect 412590 697038 422218 697098
rect 402838 696902 403082 696962
rect 422158 696962 422218 697038
rect 422342 696962 422402 697174
rect 431910 697098 431970 697174
rect 441662 697174 451290 697234
rect 431910 697038 441538 697098
rect 422158 696902 422402 696962
rect 441478 696962 441538 697038
rect 441662 696962 441722 697174
rect 451230 697098 451290 697174
rect 460982 697174 470610 697234
rect 451230 697038 460858 697098
rect 441478 696902 441722 696962
rect 460798 696962 460858 697038
rect 460982 696962 461042 697174
rect 470550 697098 470610 697174
rect 480302 697174 489930 697234
rect 470550 697038 480178 697098
rect 460798 696902 461042 696962
rect 480118 696962 480178 697038
rect 480302 696962 480362 697174
rect 489870 697098 489930 697174
rect 499622 697174 509250 697234
rect 489870 697038 499498 697098
rect 480118 696902 480362 696962
rect 499438 696962 499498 697038
rect 499622 696962 499682 697174
rect 509190 697098 509250 697174
rect 518942 697174 528570 697234
rect 509190 697038 518818 697098
rect 499438 696902 499682 696962
rect 518758 696962 518818 697038
rect 518942 696962 519002 697174
rect 528510 697098 528570 697174
rect 538262 697232 541039 697234
rect 538262 697176 540978 697232
rect 541034 697176 541039 697232
rect 538262 697174 541039 697176
rect 528510 697038 538138 697098
rect 518758 696902 519002 696962
rect 538078 696962 538138 697038
rect 538262 696962 538322 697174
rect 540973 697171 541039 697174
rect 565169 697234 565235 697237
rect 572713 697234 572779 697237
rect 565169 697232 569970 697234
rect 565169 697176 565174 697232
rect 565230 697176 569970 697232
rect 565169 697174 569970 697176
rect 565169 697171 565235 697174
rect 569910 697098 569970 697174
rect 572713 697232 576962 697234
rect 572713 697176 572718 697232
rect 572774 697176 576962 697232
rect 572713 697174 576962 697176
rect 572713 697171 572779 697174
rect 572621 697098 572687 697101
rect 569910 697096 572687 697098
rect 569910 697040 572626 697096
rect 572682 697040 572687 697096
rect 569910 697038 572687 697040
rect 576902 697098 576962 697174
rect 583342 697098 583402 697990
rect 583520 697900 584960 697990
rect 576902 697038 583402 697098
rect 572621 697035 572687 697038
rect 538078 696902 538322 696962
rect 548609 696962 548675 696965
rect 550582 696962 550588 696964
rect 548609 696960 550588 696962
rect 548609 696904 548614 696960
rect 548670 696904 550588 696960
rect 548609 696902 550588 696904
rect 548609 696899 548675 696902
rect 550582 696900 550588 696902
rect 550652 696900 550658 696964
rect -960 696540 480 696780
rect 183502 686428 183508 686492
rect 183572 686490 183578 686492
rect 188337 686490 188403 686493
rect 183572 686488 188403 686490
rect 183572 686432 188342 686488
rect 188398 686432 188403 686488
rect 183572 686430 188403 686432
rect 183572 686428 183578 686430
rect 188337 686427 188403 686430
rect 376702 686428 376708 686492
rect 376772 686490 376778 686492
rect 379513 686490 379579 686493
rect 376772 686488 379579 686490
rect 376772 686432 379518 686488
rect 379574 686432 379579 686488
rect 376772 686430 379579 686432
rect 376772 686428 376778 686430
rect 379513 686427 379579 686430
rect 434662 686428 434668 686492
rect 434732 686490 434738 686492
rect 441521 686490 441587 686493
rect 434732 686488 441587 686490
rect 434732 686432 441526 686488
rect 441582 686432 441587 686488
rect 434732 686430 441587 686432
rect 434732 686428 434738 686430
rect 441521 686427 441587 686430
rect 164182 686292 164188 686356
rect 164252 686354 164258 686356
rect 166901 686354 166967 686357
rect 164252 686352 166967 686354
rect 164252 686296 166906 686352
rect 166962 686296 166967 686352
rect 164252 686294 166967 686296
rect 164252 686292 164258 686294
rect 166901 686291 166967 686294
rect 167085 686354 167151 686357
rect 173893 686354 173959 686357
rect 167085 686352 173959 686354
rect 167085 686296 167090 686352
rect 167146 686296 173898 686352
rect 173954 686296 173959 686352
rect 167085 686294 173959 686296
rect 167085 686291 167151 686294
rect 173893 686291 173959 686294
rect 357382 686292 357388 686356
rect 357452 686354 357458 686356
rect 360101 686354 360167 686357
rect 357452 686352 360167 686354
rect 357452 686296 360106 686352
rect 360162 686296 360167 686352
rect 357452 686294 360167 686296
rect 357452 686292 357458 686294
rect 360101 686291 360167 686294
rect 360285 686354 360351 686357
rect 367093 686354 367159 686357
rect 360285 686352 367159 686354
rect 360285 686296 360290 686352
rect 360346 686296 367098 686352
rect 367154 686296 367159 686352
rect 360285 686294 367159 686296
rect 360285 686291 360351 686294
rect 367093 686291 367159 686294
rect 550582 686292 550588 686356
rect 550652 686354 550658 686356
rect 553301 686354 553367 686357
rect 550652 686352 553367 686354
rect 550652 686296 553306 686352
rect 553362 686296 553367 686352
rect 550652 686294 553367 686296
rect 550652 686292 550658 686294
rect 553301 686291 553367 686294
rect 553485 686354 553551 686357
rect 560293 686354 560359 686357
rect 583520 686354 584960 686444
rect 553485 686352 560359 686354
rect 553485 686296 553490 686352
rect 553546 686296 560298 686352
rect 560354 686296 560359 686352
rect 553485 686294 560359 686296
rect 553485 686291 553551 686294
rect 560293 686291 560359 686294
rect 583342 686294 584960 686354
rect 57830 686156 57836 686220
rect 57900 686218 57906 686220
rect 154573 686218 154639 686221
rect 57900 686158 64890 686218
rect 57900 686156 57906 686158
rect 64830 686082 64890 686158
rect 74582 686158 84210 686218
rect 64830 686022 74458 686082
rect 74398 685946 74458 686022
rect 74582 685946 74642 686158
rect 84150 686082 84210 686158
rect 93902 686158 103530 686218
rect 84150 686022 93778 686082
rect 74398 685886 74642 685946
rect 93718 685946 93778 686022
rect 93902 685946 93962 686158
rect 103470 686082 103530 686158
rect 113222 686158 122850 686218
rect 103470 686022 113098 686082
rect 93718 685886 93962 685946
rect 113038 685946 113098 686022
rect 113222 685946 113282 686158
rect 122790 686082 122850 686158
rect 132542 686158 142170 686218
rect 122790 686022 132418 686082
rect 113038 685886 113282 685946
rect 132358 685946 132418 686022
rect 132542 685946 132602 686158
rect 142110 686082 142170 686158
rect 151862 686216 154639 686218
rect 151862 686160 154578 686216
rect 154634 686160 154639 686216
rect 151862 686158 154639 686160
rect 142110 686022 151738 686082
rect 132358 685886 132602 685946
rect 151678 685946 151738 686022
rect 151862 685946 151922 686158
rect 154573 686155 154639 686158
rect 178769 686218 178835 686221
rect 183502 686218 183508 686220
rect 178769 686216 183508 686218
rect 178769 686160 178774 686216
rect 178830 686160 183508 686216
rect 178769 686158 183508 686160
rect 178769 686155 178835 686158
rect 183502 686156 183508 686158
rect 183572 686156 183578 686220
rect 188337 686218 188403 686221
rect 289813 686218 289879 686221
rect 188337 686216 200130 686218
rect 188337 686160 188342 686216
rect 188398 686160 200130 686216
rect 188337 686158 200130 686160
rect 188337 686155 188403 686158
rect 200070 686082 200130 686158
rect 209822 686158 219450 686218
rect 200070 686022 209698 686082
rect 151678 685886 151922 685946
rect 162209 685946 162275 685949
rect 164182 685946 164188 685948
rect 162209 685944 164188 685946
rect 162209 685888 162214 685944
rect 162270 685888 164188 685944
rect 162209 685886 164188 685888
rect 162209 685883 162275 685886
rect 164182 685884 164188 685886
rect 164252 685884 164258 685948
rect 209638 685946 209698 686022
rect 209822 685946 209882 686158
rect 219390 686082 219450 686158
rect 229142 686158 238770 686218
rect 219390 686022 229018 686082
rect 209638 685886 209882 685946
rect 228958 685946 229018 686022
rect 229142 685946 229202 686158
rect 238710 686082 238770 686158
rect 248462 686158 258090 686218
rect 238710 686022 248338 686082
rect 228958 685886 229202 685946
rect 248278 685946 248338 686022
rect 248462 685946 248522 686158
rect 258030 686082 258090 686158
rect 267782 686158 277410 686218
rect 258030 686022 267658 686082
rect 248278 685886 248522 685946
rect 267598 685946 267658 686022
rect 267782 685946 267842 686158
rect 277350 686082 277410 686158
rect 287102 686216 289879 686218
rect 287102 686160 289818 686216
rect 289874 686160 289879 686216
rect 287102 686158 289879 686160
rect 277350 686022 286978 686082
rect 267598 685886 267842 685946
rect 286918 685946 286978 686022
rect 287102 685946 287162 686158
rect 289813 686155 289879 686158
rect 299422 686156 299428 686220
rect 299492 686218 299498 686220
rect 347773 686218 347839 686221
rect 299492 686158 316050 686218
rect 299492 686156 299498 686158
rect 315990 686082 316050 686158
rect 325742 686158 335370 686218
rect 315990 686022 325618 686082
rect 286918 685886 287162 685946
rect 294505 685946 294571 685949
rect 299422 685946 299428 685948
rect 294505 685944 299428 685946
rect 294505 685888 294510 685944
rect 294566 685888 299428 685944
rect 294505 685886 299428 685888
rect 294505 685883 294571 685886
rect 299422 685884 299428 685886
rect 299492 685884 299498 685948
rect 325558 685946 325618 686022
rect 325742 685946 325802 686158
rect 335310 686082 335370 686158
rect 345062 686216 347839 686218
rect 345062 686160 347778 686216
rect 347834 686160 347839 686216
rect 345062 686158 347839 686160
rect 335310 686022 344938 686082
rect 325558 685886 325802 685946
rect 344878 685946 344938 686022
rect 345062 685946 345122 686158
rect 347773 686155 347839 686158
rect 371969 686218 372035 686221
rect 376702 686218 376708 686220
rect 371969 686216 376708 686218
rect 371969 686160 371974 686216
rect 372030 686160 376708 686216
rect 371969 686158 376708 686160
rect 371969 686155 372035 686158
rect 376702 686156 376708 686158
rect 376772 686156 376778 686220
rect 379513 686218 379579 686221
rect 427537 686218 427603 686221
rect 379513 686216 393330 686218
rect 379513 686160 379518 686216
rect 379574 686160 393330 686216
rect 379513 686158 393330 686160
rect 379513 686155 379579 686158
rect 393270 686082 393330 686158
rect 403022 686216 427603 686218
rect 403022 686160 427542 686216
rect 427598 686160 427603 686216
rect 403022 686158 427603 686160
rect 393270 686022 402898 686082
rect 344878 685886 345122 685946
rect 355409 685946 355475 685949
rect 357382 685946 357388 685948
rect 355409 685944 357388 685946
rect 355409 685888 355414 685944
rect 355470 685888 357388 685944
rect 355409 685886 357388 685888
rect 355409 685883 355475 685886
rect 357382 685884 357388 685886
rect 357452 685884 357458 685948
rect 402838 685946 402898 686022
rect 403022 685946 403082 686158
rect 427537 686155 427603 686158
rect 427721 686218 427787 686221
rect 441521 686218 441587 686221
rect 540973 686218 541039 686221
rect 427721 686216 429762 686218
rect 427721 686160 427726 686216
rect 427782 686160 429762 686216
rect 427721 686158 429762 686160
rect 427721 686155 427787 686158
rect 429702 686082 429762 686158
rect 441521 686216 451290 686218
rect 441521 686160 441526 686216
rect 441582 686160 451290 686216
rect 441521 686158 451290 686160
rect 441521 686155 441587 686158
rect 434662 686082 434668 686084
rect 429702 686022 434668 686082
rect 434662 686020 434668 686022
rect 434732 686020 434738 686084
rect 451230 686082 451290 686158
rect 460982 686158 470610 686218
rect 451230 686022 460858 686082
rect 402838 685886 403082 685946
rect 460798 685946 460858 686022
rect 460982 685946 461042 686158
rect 470550 686082 470610 686158
rect 480302 686158 489930 686218
rect 470550 686022 480178 686082
rect 460798 685886 461042 685946
rect 480118 685946 480178 686022
rect 480302 685946 480362 686158
rect 489870 686082 489930 686158
rect 499622 686158 509250 686218
rect 489870 686022 499498 686082
rect 480118 685886 480362 685946
rect 499438 685946 499498 686022
rect 499622 685946 499682 686158
rect 509190 686082 509250 686158
rect 518942 686158 528570 686218
rect 509190 686022 518818 686082
rect 499438 685886 499682 685946
rect 518758 685946 518818 686022
rect 518942 685946 519002 686158
rect 528510 686082 528570 686158
rect 538262 686216 541039 686218
rect 538262 686160 540978 686216
rect 541034 686160 541039 686216
rect 538262 686158 541039 686160
rect 528510 686022 538138 686082
rect 518758 685886 519002 685946
rect 538078 685946 538138 686022
rect 538262 685946 538322 686158
rect 540973 686155 541039 686158
rect 565169 686218 565235 686221
rect 572713 686218 572779 686221
rect 565169 686216 569970 686218
rect 565169 686160 565174 686216
rect 565230 686160 569970 686216
rect 565169 686158 569970 686160
rect 565169 686155 565235 686158
rect 569910 686082 569970 686158
rect 572713 686216 576962 686218
rect 572713 686160 572718 686216
rect 572774 686160 576962 686216
rect 572713 686158 576962 686160
rect 572713 686155 572779 686158
rect 572621 686082 572687 686085
rect 569910 686080 572687 686082
rect 569910 686024 572626 686080
rect 572682 686024 572687 686080
rect 569910 686022 572687 686024
rect 576902 686082 576962 686158
rect 583342 686082 583402 686294
rect 583520 686204 584960 686294
rect 576902 686022 583402 686082
rect 572621 686019 572687 686022
rect 538078 685886 538322 685946
rect 548609 685946 548675 685949
rect 550582 685946 550588 685948
rect 548609 685944 550588 685946
rect 548609 685888 548614 685944
rect 548670 685888 550588 685944
rect 548609 685886 550588 685888
rect 548609 685883 548675 685886
rect 550582 685884 550588 685886
rect 550652 685884 550658 685948
rect 559005 684448 559071 684453
rect 559005 684392 559010 684448
rect 559066 684392 559071 684448
rect 559005 684387 559071 684392
rect 559008 684317 559068 684387
rect 559005 684312 559071 684317
rect 559005 684256 559010 684312
rect 559066 684256 559071 684312
rect 559005 684251 559071 684256
rect -960 682274 480 682364
rect 2773 682274 2839 682277
rect -960 682272 2839 682274
rect -960 682216 2778 682272
rect 2834 682216 2839 682272
rect -960 682214 2839 682216
rect -960 682124 480 682214
rect 2773 682211 2839 682214
rect 583520 674658 584960 674748
rect 583342 674598 584960 674658
rect 183502 674052 183508 674116
rect 183572 674114 183578 674116
rect 188337 674114 188403 674117
rect 183572 674112 188403 674114
rect 183572 674056 188342 674112
rect 188398 674056 188403 674112
rect 183572 674054 188403 674056
rect 183572 674052 183578 674054
rect 188337 674051 188403 674054
rect 376702 674052 376708 674116
rect 376772 674114 376778 674116
rect 379513 674114 379579 674117
rect 376772 674112 379579 674114
rect 376772 674056 379518 674112
rect 379574 674056 379579 674112
rect 376772 674054 379579 674056
rect 376772 674052 376778 674054
rect 379513 674051 379579 674054
rect 166993 673978 167059 673981
rect 173893 673978 173959 673981
rect 166993 673976 173959 673978
rect 166993 673920 166998 673976
rect 167054 673920 173898 673976
rect 173954 673920 173959 673976
rect 166993 673918 173959 673920
rect 166993 673915 167059 673918
rect 173893 673915 173959 673918
rect 357382 673916 357388 673980
rect 357452 673978 357458 673980
rect 360101 673978 360167 673981
rect 357452 673976 360167 673978
rect 357452 673920 360106 673976
rect 360162 673920 360167 673976
rect 357452 673918 360167 673920
rect 357452 673916 357458 673918
rect 360101 673915 360167 673918
rect 360285 673978 360351 673981
rect 367093 673978 367159 673981
rect 360285 673976 367159 673978
rect 360285 673920 360290 673976
rect 360346 673920 367098 673976
rect 367154 673920 367159 673976
rect 360285 673918 367159 673920
rect 360285 673915 360351 673918
rect 367093 673915 367159 673918
rect 553393 673978 553459 673981
rect 560293 673978 560359 673981
rect 553393 673976 560359 673978
rect 553393 673920 553398 673976
rect 553454 673920 560298 673976
rect 560354 673920 560359 673976
rect 553393 673918 560359 673920
rect 553393 673915 553459 673918
rect 560293 673915 560359 673918
rect 58198 673780 58204 673844
rect 58268 673842 58274 673844
rect 154573 673842 154639 673845
rect 58268 673782 64890 673842
rect 58268 673780 58274 673782
rect 64830 673706 64890 673782
rect 74582 673782 84210 673842
rect 64830 673646 74458 673706
rect 74398 673570 74458 673646
rect 74582 673570 74642 673782
rect 84150 673706 84210 673782
rect 93902 673782 103530 673842
rect 84150 673646 93778 673706
rect 74398 673510 74642 673570
rect 93718 673570 93778 673646
rect 93902 673570 93962 673782
rect 103470 673706 103530 673782
rect 113222 673782 122850 673842
rect 103470 673646 113098 673706
rect 93718 673510 93962 673570
rect 113038 673570 113098 673646
rect 113222 673570 113282 673782
rect 122790 673706 122850 673782
rect 132542 673782 142170 673842
rect 122790 673646 132418 673706
rect 113038 673510 113282 673570
rect 132358 673570 132418 673646
rect 132542 673570 132602 673782
rect 142110 673706 142170 673782
rect 151862 673840 154639 673842
rect 151862 673784 154578 673840
rect 154634 673784 154639 673840
rect 151862 673782 154639 673784
rect 142110 673646 151738 673706
rect 132358 673510 132602 673570
rect 151678 673570 151738 673646
rect 151862 673570 151922 673782
rect 154573 673779 154639 673782
rect 178769 673842 178835 673845
rect 183502 673842 183508 673844
rect 178769 673840 183508 673842
rect 178769 673784 178774 673840
rect 178830 673784 183508 673840
rect 178769 673782 183508 673784
rect 178769 673779 178835 673782
rect 183502 673780 183508 673782
rect 183572 673780 183578 673844
rect 188337 673842 188403 673845
rect 289813 673842 289879 673845
rect 188337 673840 200130 673842
rect 188337 673784 188342 673840
rect 188398 673784 200130 673840
rect 188337 673782 200130 673784
rect 188337 673779 188403 673782
rect 200070 673706 200130 673782
rect 209822 673782 219450 673842
rect 200070 673646 209698 673706
rect 151678 673510 151922 673570
rect 162209 673570 162275 673573
rect 166901 673570 166967 673573
rect 162209 673568 166967 673570
rect 162209 673512 162214 673568
rect 162270 673512 166906 673568
rect 166962 673512 166967 673568
rect 162209 673510 166967 673512
rect 209638 673570 209698 673646
rect 209822 673570 209882 673782
rect 219390 673706 219450 673782
rect 229142 673782 238770 673842
rect 219390 673646 229018 673706
rect 209638 673510 209882 673570
rect 228958 673570 229018 673646
rect 229142 673570 229202 673782
rect 238710 673706 238770 673782
rect 248462 673782 258090 673842
rect 238710 673646 248338 673706
rect 228958 673510 229202 673570
rect 248278 673570 248338 673646
rect 248462 673570 248522 673782
rect 258030 673706 258090 673782
rect 267782 673782 277410 673842
rect 258030 673646 267658 673706
rect 248278 673510 248522 673570
rect 267598 673570 267658 673646
rect 267782 673570 267842 673782
rect 277350 673706 277410 673782
rect 287102 673840 289879 673842
rect 287102 673784 289818 673840
rect 289874 673784 289879 673840
rect 287102 673782 289879 673784
rect 277350 673646 286978 673706
rect 267598 673510 267842 673570
rect 286918 673570 286978 673646
rect 287102 673570 287162 673782
rect 289813 673779 289879 673782
rect 299422 673780 299428 673844
rect 299492 673842 299498 673844
rect 347773 673842 347839 673845
rect 299492 673782 316050 673842
rect 299492 673780 299498 673782
rect 315990 673706 316050 673782
rect 325742 673782 335370 673842
rect 315990 673646 325618 673706
rect 286918 673510 287162 673570
rect 292665 673570 292731 673573
rect 299422 673570 299428 673572
rect 292665 673568 299428 673570
rect 292665 673512 292670 673568
rect 292726 673512 299428 673568
rect 292665 673510 299428 673512
rect 162209 673507 162275 673510
rect 166901 673507 166967 673510
rect 292665 673507 292731 673510
rect 299422 673508 299428 673510
rect 299492 673508 299498 673572
rect 325558 673570 325618 673646
rect 325742 673570 325802 673782
rect 335310 673706 335370 673782
rect 345062 673840 347839 673842
rect 345062 673784 347778 673840
rect 347834 673784 347839 673840
rect 345062 673782 347839 673784
rect 335310 673646 344938 673706
rect 325558 673510 325802 673570
rect 344878 673570 344938 673646
rect 345062 673570 345122 673782
rect 347773 673779 347839 673782
rect 371969 673842 372035 673845
rect 376702 673842 376708 673844
rect 371969 673840 376708 673842
rect 371969 673784 371974 673840
rect 372030 673784 376708 673840
rect 371969 673782 376708 673784
rect 371969 673779 372035 673782
rect 376702 673780 376708 673782
rect 376772 673780 376778 673844
rect 379513 673842 379579 673845
rect 540973 673842 541039 673845
rect 379513 673840 393330 673842
rect 379513 673784 379518 673840
rect 379574 673784 393330 673840
rect 379513 673782 393330 673784
rect 379513 673779 379579 673782
rect 393270 673706 393330 673782
rect 403022 673782 412650 673842
rect 393270 673646 402898 673706
rect 344878 673510 345122 673570
rect 355409 673570 355475 673573
rect 357382 673570 357388 673572
rect 355409 673568 357388 673570
rect 355409 673512 355414 673568
rect 355470 673512 357388 673568
rect 355409 673510 357388 673512
rect 355409 673507 355475 673510
rect 357382 673508 357388 673510
rect 357452 673508 357458 673572
rect 402838 673570 402898 673646
rect 403022 673570 403082 673782
rect 412590 673706 412650 673782
rect 431910 673782 441538 673842
rect 412590 673646 422218 673706
rect 402838 673510 403082 673570
rect 422158 673570 422218 673646
rect 431910 673570 431970 673782
rect 422158 673510 431970 673570
rect 441478 673570 441538 673782
rect 441662 673782 451290 673842
rect 441662 673570 441722 673782
rect 451230 673706 451290 673782
rect 460982 673782 470610 673842
rect 451230 673646 460858 673706
rect 441478 673510 441722 673570
rect 460798 673570 460858 673646
rect 460982 673570 461042 673782
rect 470550 673706 470610 673782
rect 480302 673782 489930 673842
rect 470550 673646 480178 673706
rect 460798 673510 461042 673570
rect 480118 673570 480178 673646
rect 480302 673570 480362 673782
rect 489870 673706 489930 673782
rect 499622 673782 509250 673842
rect 489870 673646 499498 673706
rect 480118 673510 480362 673570
rect 499438 673570 499498 673646
rect 499622 673570 499682 673782
rect 509190 673706 509250 673782
rect 518942 673782 528570 673842
rect 509190 673646 518818 673706
rect 499438 673510 499682 673570
rect 518758 673570 518818 673646
rect 518942 673570 519002 673782
rect 528510 673706 528570 673782
rect 538262 673840 541039 673842
rect 538262 673784 540978 673840
rect 541034 673784 541039 673840
rect 538262 673782 541039 673784
rect 528510 673646 538138 673706
rect 518758 673510 519002 673570
rect 538078 673570 538138 673646
rect 538262 673570 538322 673782
rect 540973 673779 541039 673782
rect 565169 673842 565235 673845
rect 572713 673842 572779 673845
rect 565169 673840 569970 673842
rect 565169 673784 565174 673840
rect 565230 673784 569970 673840
rect 565169 673782 569970 673784
rect 565169 673779 565235 673782
rect 569910 673706 569970 673782
rect 572713 673840 576962 673842
rect 572713 673784 572718 673840
rect 572774 673784 576962 673840
rect 572713 673782 576962 673784
rect 572713 673779 572779 673782
rect 572621 673706 572687 673709
rect 569910 673704 572687 673706
rect 569910 673648 572626 673704
rect 572682 673648 572687 673704
rect 569910 673646 572687 673648
rect 576902 673706 576962 673782
rect 583342 673706 583402 674598
rect 583520 674508 584960 674598
rect 576902 673646 583402 673706
rect 572621 673643 572687 673646
rect 538078 673510 538322 673570
rect 548609 673570 548675 673573
rect 553301 673570 553367 673573
rect 548609 673568 553367 673570
rect 548609 673512 548614 673568
rect 548670 673512 553306 673568
rect 553362 673512 553367 673568
rect 548609 673510 553367 673512
rect 548609 673507 548675 673510
rect 553301 673507 553367 673510
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 169845 666634 169911 666637
rect 170029 666634 170095 666637
rect 169845 666632 170095 666634
rect 169845 666576 169850 666632
rect 169906 666576 170034 666632
rect 170090 666576 170095 666632
rect 169845 666574 170095 666576
rect 169845 666571 169911 666574
rect 170029 666571 170095 666574
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 129273 652900 129339 652901
rect 129222 652898 129228 652900
rect 129182 652838 129228 652898
rect 129292 652896 129339 652900
rect 129334 652840 129339 652896
rect 129222 652836 129228 652838
rect 129292 652836 129339 652840
rect 129273 652835 129339 652836
rect 133597 652900 133663 652901
rect 259177 652900 259243 652901
rect 263777 652900 263843 652901
rect 133597 652896 133644 652900
rect 133708 652898 133714 652900
rect 259126 652898 259132 652900
rect 133597 652840 133602 652896
rect 133597 652836 133644 652840
rect 133708 652838 133754 652898
rect 259086 652838 259132 652898
rect 259196 652896 259243 652900
rect 263726 652898 263732 652900
rect 259238 652840 259243 652896
rect 133708 652836 133714 652838
rect 259126 652836 259132 652838
rect 259196 652836 259243 652840
rect 263686 652838 263732 652898
rect 263796 652896 263843 652900
rect 263838 652840 263843 652896
rect 263726 652836 263732 652838
rect 263796 652836 263843 652840
rect 133597 652835 133663 652836
rect 259177 652835 259243 652836
rect 263777 652835 263843 652836
rect 378501 652900 378567 652901
rect 383469 652900 383535 652901
rect 507853 652900 507919 652901
rect 513373 652900 513439 652901
rect 378501 652896 378548 652900
rect 378612 652898 378618 652900
rect 378501 652840 378506 652896
rect 378501 652836 378548 652840
rect 378612 652838 378658 652898
rect 383469 652896 383516 652900
rect 383580 652898 383586 652900
rect 383469 652840 383474 652896
rect 378612 652836 378618 652838
rect 383469 652836 383516 652840
rect 383580 652838 383626 652898
rect 507853 652896 507900 652900
rect 507964 652898 507970 652900
rect 507853 652840 507858 652896
rect 383580 652836 383586 652838
rect 507853 652836 507900 652840
rect 507964 652838 508010 652898
rect 513373 652896 513420 652900
rect 513484 652898 513490 652900
rect 513373 652840 513378 652896
rect 507964 652836 507970 652838
rect 513373 652836 513420 652840
rect 513484 652838 513530 652898
rect 513484 652836 513490 652838
rect 378501 652835 378567 652836
rect 383469 652835 383535 652836
rect 507853 652835 507919 652836
rect 513373 652835 513439 652836
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 139393 649906 139459 649909
rect 137142 649904 139459 649906
rect 137142 649848 139398 649904
rect 139454 649848 139459 649904
rect 137142 649846 139459 649848
rect 137142 649683 137202 649846
rect 139393 649843 139459 649846
rect 266445 649906 266511 649909
rect 389173 649906 389239 649909
rect 266445 649904 266554 649906
rect 266445 649848 266450 649904
rect 266506 649848 266554 649904
rect 266445 649843 266554 649848
rect 266494 649683 266554 649843
rect 387198 649904 389239 649906
rect 387198 649848 389178 649904
rect 389234 649848 389239 649904
rect 387198 649846 389239 649848
rect 387198 649683 387258 649846
rect 389173 649843 389239 649846
rect 516409 649906 516475 649909
rect 516409 649904 516610 649906
rect 516409 649848 516414 649904
rect 516470 649848 516610 649904
rect 516409 649846 516610 649848
rect 516409 649843 516475 649846
rect 516550 649683 516610 649846
rect 56593 646098 56659 646101
rect 60046 646098 60106 646587
rect 187693 646234 187759 646237
rect 190134 646234 190194 646587
rect 187693 646232 190194 646234
rect 187693 646176 187698 646232
rect 187754 646176 190194 646232
rect 187693 646174 190194 646176
rect 187693 646171 187759 646174
rect 56593 646096 60106 646098
rect 56593 646040 56598 646096
rect 56654 646040 60106 646096
rect 56593 646038 60106 646040
rect 307385 646098 307451 646101
rect 310102 646098 310162 646587
rect 437473 646234 437539 646237
rect 440006 646234 440066 646587
rect 437473 646232 440066 646234
rect 437473 646176 437478 646232
rect 437534 646176 440066 646232
rect 437473 646174 440066 646176
rect 437473 646171 437539 646174
rect 307385 646096 310162 646098
rect 307385 646040 307390 646096
rect 307446 646040 310162 646096
rect 307385 646038 310162 646040
rect 56593 646035 56659 646038
rect 307385 646035 307451 646038
rect 169753 645962 169819 645965
rect 170029 645962 170095 645965
rect 169753 645960 170095 645962
rect 169753 645904 169758 645960
rect 169814 645904 170034 645960
rect 170090 645904 170095 645960
rect 169753 645902 170095 645904
rect 169753 645899 169819 645902
rect 170029 645899 170095 645902
rect 57237 645010 57303 645013
rect 60046 645010 60106 645459
rect 57237 645008 60106 645010
rect 57237 644952 57242 645008
rect 57298 644952 60106 645008
rect 57237 644950 60106 644952
rect 57237 644947 57303 644950
rect 187693 644874 187759 644877
rect 190134 644874 190194 645459
rect 307109 645010 307175 645013
rect 310102 645010 310162 645459
rect 307109 645008 310162 645010
rect 307109 644952 307114 645008
rect 307170 644952 310162 645008
rect 307109 644950 310162 644952
rect 307109 644947 307175 644950
rect 187693 644872 190194 644874
rect 187693 644816 187698 644872
rect 187754 644816 190194 644872
rect 187693 644814 190194 644816
rect 437473 644874 437539 644877
rect 440006 644874 440066 645459
rect 437473 644872 440066 644874
rect 437473 644816 437478 644872
rect 437534 644816 440066 644872
rect 437473 644814 440066 644816
rect 187693 644811 187759 644814
rect 437473 644811 437539 644814
rect 57145 643242 57211 643245
rect 60046 643242 60106 643759
rect 57145 643240 60106 643242
rect 57145 643184 57150 643240
rect 57206 643184 60106 643240
rect 57145 643182 60106 643184
rect 187693 643242 187759 643245
rect 190134 643242 190194 643759
rect 307109 643514 307175 643517
rect 310102 643514 310162 643759
rect 307109 643512 310162 643514
rect 307109 643456 307114 643512
rect 307170 643456 310162 643512
rect 307109 643454 310162 643456
rect 307109 643451 307175 643454
rect 187693 643240 190194 643242
rect 187693 643184 187698 643240
rect 187754 643184 190194 643240
rect 187693 643182 190194 643184
rect 437473 643242 437539 643245
rect 440006 643242 440066 643759
rect 437473 643240 440066 643242
rect 437473 643184 437478 643240
rect 437534 643184 440066 643240
rect 437473 643182 440066 643184
rect 57145 643179 57211 643182
rect 187693 643179 187759 643182
rect 437473 643179 437539 643182
rect 57053 642018 57119 642021
rect 60046 642018 60106 642631
rect 57053 642016 60106 642018
rect 57053 641960 57058 642016
rect 57114 641960 60106 642016
rect 57053 641958 60106 641960
rect 187693 642018 187759 642021
rect 190134 642018 190194 642631
rect 307661 642154 307727 642157
rect 310102 642154 310162 642631
rect 307661 642152 310162 642154
rect 307661 642096 307666 642152
rect 307722 642096 310162 642152
rect 307661 642094 310162 642096
rect 307661 642091 307727 642094
rect 187693 642016 190194 642018
rect 187693 641960 187698 642016
rect 187754 641960 190194 642016
rect 187693 641958 190194 641960
rect 437473 642018 437539 642021
rect 440006 642018 440066 642631
rect 437473 642016 440066 642018
rect 437473 641960 437478 642016
rect 437534 641960 440066 642016
rect 437473 641958 440066 641960
rect 57053 641955 57119 641958
rect 187693 641955 187759 641958
rect 437473 641955 437539 641958
rect 56961 640386 57027 640389
rect 60046 640386 60106 640931
rect 56961 640384 60106 640386
rect 56961 640328 56966 640384
rect 57022 640328 60106 640384
rect 56961 640326 60106 640328
rect 187693 640386 187759 640389
rect 190134 640386 190194 640931
rect 307661 640522 307727 640525
rect 310102 640522 310162 640931
rect 307661 640520 310162 640522
rect 307661 640464 307666 640520
rect 307722 640464 310162 640520
rect 307661 640462 310162 640464
rect 307661 640459 307727 640462
rect 187693 640384 190194 640386
rect 187693 640328 187698 640384
rect 187754 640328 190194 640384
rect 187693 640326 190194 640328
rect 437473 640386 437539 640389
rect 440006 640386 440066 640931
rect 437473 640384 440066 640386
rect 437473 640328 437478 640384
rect 437534 640328 440066 640384
rect 437473 640326 440066 640328
rect 56961 640323 57027 640326
rect 187693 640323 187759 640326
rect 437473 640323 437539 640326
rect 56869 639298 56935 639301
rect 60046 639298 60106 639803
rect 56869 639296 60106 639298
rect -960 639012 480 639252
rect 56869 639240 56874 639296
rect 56930 639240 60106 639296
rect 56869 639238 60106 639240
rect 188337 639298 188403 639301
rect 190134 639298 190194 639803
rect 306649 639434 306715 639437
rect 310102 639434 310162 639803
rect 306649 639432 310162 639434
rect 306649 639376 306654 639432
rect 306710 639376 310162 639432
rect 306649 639374 310162 639376
rect 306649 639371 306715 639374
rect 188337 639296 190194 639298
rect 188337 639240 188342 639296
rect 188398 639240 190194 639296
rect 188337 639238 190194 639240
rect 437473 639298 437539 639301
rect 440006 639298 440066 639803
rect 580257 639434 580323 639437
rect 583520 639434 584960 639524
rect 580257 639432 584960 639434
rect 580257 639376 580262 639432
rect 580318 639376 584960 639432
rect 580257 639374 584960 639376
rect 580257 639371 580323 639374
rect 437473 639296 440066 639298
rect 437473 639240 437478 639296
rect 437534 639240 440066 639296
rect 583520 639284 584960 639374
rect 437473 639238 440066 639240
rect 56869 639235 56935 639238
rect 188337 639235 188403 639238
rect 437473 639235 437539 639238
rect 56777 637666 56843 637669
rect 60046 637666 60106 638103
rect 56777 637664 60106 637666
rect 56777 637608 56782 637664
rect 56838 637608 60106 637664
rect 56777 637606 60106 637608
rect 188429 637666 188495 637669
rect 190134 637666 190194 638103
rect 299565 637938 299631 637941
rect 310102 637938 310162 638103
rect 299565 637936 310162 637938
rect 299565 637880 299570 637936
rect 299626 637880 310162 637936
rect 299565 637878 310162 637880
rect 299565 637875 299631 637878
rect 188429 637664 190194 637666
rect 188429 637608 188434 637664
rect 188490 637608 190194 637664
rect 188429 637606 190194 637608
rect 437473 637666 437539 637669
rect 440006 637666 440066 638103
rect 437473 637664 440066 637666
rect 437473 637608 437478 637664
rect 437534 637608 440066 637664
rect 437473 637606 440066 637608
rect 56777 637603 56843 637606
rect 188429 637603 188495 637606
rect 437473 637603 437539 637606
rect 299657 637530 299723 637533
rect 300025 637530 300091 637533
rect 299657 637528 300091 637530
rect 299657 637472 299662 637528
rect 299718 637472 300030 637528
rect 300086 637472 300091 637528
rect 299657 637470 300091 637472
rect 299657 637467 299723 637470
rect 300025 637467 300091 637470
rect 580349 627738 580415 627741
rect 583520 627738 584960 627828
rect 580349 627736 584960 627738
rect 580349 627680 580354 627736
rect 580410 627680 584960 627736
rect 580349 627678 584960 627680
rect 580349 627675 580415 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3877 624882 3943 624885
rect -960 624880 3943 624882
rect -960 624824 3882 624880
rect 3938 624824 3943 624880
rect -960 624822 3943 624824
rect -960 624732 480 624822
rect 3877 624819 3943 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580441 604210 580507 604213
rect 583520 604210 584960 604300
rect 580441 604208 584960 604210
rect 580441 604152 580446 604208
rect 580502 604152 584960 604208
rect 580441 604150 584960 604152
rect 580441 604147 580507 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580533 592514 580599 592517
rect 583520 592514 584960 592604
rect 580533 592512 584960 592514
rect 580533 592456 580538 592512
rect 580594 592456 584960 592512
rect 580533 592454 584960 592456
rect 580533 592451 580599 592454
rect 583520 592364 584960 592454
rect 139393 589658 139459 589661
rect 389173 589658 389239 589661
rect 136958 589656 139459 589658
rect 136958 589600 139398 589656
rect 139454 589600 139459 589656
rect 136958 589598 139459 589600
rect 136958 586614 137018 589598
rect 139393 589595 139459 589598
rect 387014 589656 389239 589658
rect 387014 589600 389178 589656
rect 389234 589600 389239 589656
rect 387014 589598 389239 589600
rect 267230 589386 267290 589412
rect 269113 589386 269179 589389
rect 267230 589384 269179 589386
rect 267230 589328 269118 589384
rect 269174 589328 269179 589384
rect 267230 589326 269179 589328
rect 269113 589323 269179 589326
rect 170029 587890 170095 587893
rect 170305 587890 170371 587893
rect 170029 587888 170371 587890
rect 170029 587832 170034 587888
rect 170090 587832 170310 587888
rect 170366 587832 170371 587888
rect 170029 587830 170371 587832
rect 170029 587827 170095 587830
rect 170305 587827 170371 587830
rect 269113 587754 269179 587757
rect 267230 587752 269179 587754
rect 267230 587696 269118 587752
rect 269174 587696 269179 587752
rect 267230 587694 269179 587696
rect 136958 586584 137172 586614
rect 136988 586554 137202 586584
rect -960 581620 480 581860
rect 137142 580928 137202 586554
rect 267230 580954 267290 587694
rect 269113 587691 269179 587694
rect 387014 586614 387074 589598
rect 389173 589595 389239 589598
rect 517102 589386 517162 589412
rect 518893 589386 518959 589389
rect 517102 589384 518959 589386
rect 517102 589328 518898 589384
rect 518954 589328 518959 589384
rect 517102 589326 518959 589328
rect 518893 589323 518959 589326
rect 518893 587754 518959 587757
rect 517102 587752 518959 587754
rect 517102 587696 518898 587752
rect 518954 587696 518959 587752
rect 517102 587694 518959 587696
rect 387014 586584 387228 586614
rect 387044 586554 387258 586584
rect 270033 580954 270099 580957
rect 267230 580952 270099 580954
rect 267230 580896 270038 580952
rect 270094 580896 270099 580952
rect 387198 580928 387258 586554
rect 517102 580928 517162 587694
rect 518893 587691 518959 587694
rect 267230 580894 270099 580896
rect 270033 580891 270099 580894
rect 580625 580818 580691 580821
rect 583520 580818 584960 580908
rect 580625 580816 584960 580818
rect 580625 580760 580630 580816
rect 580686 580760 584960 580816
rect 580625 580758 584960 580760
rect 580625 580755 580691 580758
rect 583520 580668 584960 580758
rect 56685 579730 56751 579733
rect 60046 579730 60106 580255
rect 56685 579728 60106 579730
rect 56685 579672 56690 579728
rect 56746 579672 60106 579728
rect 56685 579670 60106 579672
rect 187693 579730 187759 579733
rect 190134 579730 190194 580255
rect 306925 580002 306991 580005
rect 310102 580002 310162 580255
rect 306925 580000 310162 580002
rect 306925 579944 306930 580000
rect 306986 579944 310162 580000
rect 306925 579942 310162 579944
rect 306925 579939 306991 579942
rect 187693 579728 190194 579730
rect 187693 579672 187698 579728
rect 187754 579672 190194 579728
rect 187693 579670 190194 579672
rect 437473 579730 437539 579733
rect 440006 579730 440066 580255
rect 437473 579728 440066 579730
rect 437473 579672 437478 579728
rect 437534 579672 440066 579728
rect 437473 579670 440066 579672
rect 56685 579667 56751 579670
rect 187693 579667 187759 579670
rect 437473 579667 437539 579670
rect 59629 578585 59695 578588
rect 59629 578583 60076 578585
rect 59629 578527 59634 578583
rect 59690 578527 60076 578583
rect 59629 578525 60076 578527
rect 59629 578522 59695 578525
rect 188981 578370 189047 578373
rect 190134 578370 190194 578555
rect 188981 578368 190194 578370
rect 188981 578312 188986 578368
rect 189042 578312 190194 578368
rect 188981 578310 190194 578312
rect 306373 578370 306439 578373
rect 310102 578370 310162 578555
rect 306373 578368 310162 578370
rect 306373 578312 306378 578368
rect 306434 578312 310162 578368
rect 306373 578310 310162 578312
rect 438117 578370 438183 578373
rect 440006 578370 440066 578555
rect 438117 578368 440066 578370
rect 438117 578312 438122 578368
rect 438178 578312 440066 578368
rect 438117 578310 440066 578312
rect 188981 578307 189047 578310
rect 306373 578307 306439 578310
rect 438117 578307 438183 578310
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3969 567354 4035 567357
rect -960 567352 4035 567354
rect -960 567296 3974 567352
rect 4030 567296 4035 567352
rect -960 567294 4035 567296
rect -960 567204 480 567294
rect 3969 567291 4035 567294
rect 211061 560012 211127 560013
rect 211061 560008 211108 560012
rect 211172 560010 211178 560012
rect 211061 559952 211066 560008
rect 211061 559948 211108 559952
rect 211172 559950 211218 560010
rect 211172 559948 211178 559950
rect 211061 559947 211127 559948
rect 210417 559874 210483 559877
rect 210550 559874 210556 559876
rect 210417 559872 210556 559874
rect 210417 559816 210422 559872
rect 210478 559816 210556 559872
rect 210417 559814 210556 559816
rect 210417 559811 210483 559814
rect 210550 559812 210556 559814
rect 210620 559812 210626 559876
rect 347957 559330 348023 559333
rect 351862 559330 351868 559332
rect 347957 559328 351868 559330
rect 347957 559272 347962 559328
rect 348018 559272 351868 559328
rect 347957 559270 351868 559272
rect 347957 559267 348023 559270
rect 351862 559268 351868 559270
rect 351932 559268 351938 559332
rect 357709 559330 357775 559333
rect 358854 559330 358860 559332
rect 357709 559328 358860 559330
rect 357709 559272 357714 559328
rect 357770 559272 358860 559328
rect 357709 559270 358860 559272
rect 357709 559267 357775 559270
rect 358854 559268 358860 559270
rect 358924 559268 358930 559332
rect 67398 558860 67404 558924
rect 67468 558922 67474 558924
rect 67541 558922 67607 558925
rect 67468 558920 67607 558922
rect 67468 558864 67546 558920
rect 67602 558864 67607 558920
rect 67468 558862 67607 558864
rect 67468 558860 67474 558862
rect 67541 558859 67607 558862
rect 69790 558860 69796 558924
rect 69860 558922 69866 558924
rect 70117 558922 70183 558925
rect 72417 558924 72483 558925
rect 73705 558924 73771 558925
rect 72366 558922 72372 558924
rect 69860 558920 70183 558922
rect 69860 558864 70122 558920
rect 70178 558864 70183 558920
rect 69860 558862 70183 558864
rect 72326 558862 72372 558922
rect 72436 558920 72483 558924
rect 73654 558922 73660 558924
rect 72478 558864 72483 558920
rect 69860 558860 69866 558862
rect 70117 558859 70183 558862
rect 72366 558860 72372 558862
rect 72436 558860 72483 558864
rect 73614 558862 73660 558922
rect 73724 558920 73771 558924
rect 73766 558864 73771 558920
rect 73654 558860 73660 558862
rect 73724 558860 73771 558864
rect 74942 558860 74948 558924
rect 75012 558922 75018 558924
rect 75729 558922 75795 558925
rect 75012 558920 75795 558922
rect 75012 558864 75734 558920
rect 75790 558864 75795 558920
rect 75012 558862 75795 558864
rect 75012 558860 75018 558862
rect 72417 558859 72483 558860
rect 73705 558859 73771 558860
rect 75729 558859 75795 558862
rect 75862 558860 75868 558924
rect 75932 558922 75938 558924
rect 76005 558922 76071 558925
rect 77385 558924 77451 558925
rect 78489 558924 78555 558925
rect 77334 558922 77340 558924
rect 75932 558920 76071 558922
rect 75932 558864 76010 558920
rect 76066 558864 76071 558920
rect 75932 558862 76071 558864
rect 77294 558862 77340 558922
rect 77404 558920 77451 558924
rect 78438 558922 78444 558924
rect 77446 558864 77451 558920
rect 75932 558860 75938 558862
rect 76005 558859 76071 558862
rect 77334 558860 77340 558862
rect 77404 558860 77451 558864
rect 78398 558862 78444 558922
rect 78508 558920 78555 558924
rect 78550 558864 78555 558920
rect 78438 558860 78444 558862
rect 78508 558860 78555 558864
rect 79358 558860 79364 558924
rect 79428 558922 79434 558924
rect 79501 558922 79567 558925
rect 80697 558924 80763 558925
rect 80646 558922 80652 558924
rect 79428 558920 79567 558922
rect 79428 558864 79506 558920
rect 79562 558864 79567 558920
rect 79428 558862 79567 558864
rect 80606 558862 80652 558922
rect 80716 558920 80763 558924
rect 80758 558864 80763 558920
rect 79428 558860 79434 558862
rect 77385 558859 77451 558860
rect 78489 558859 78555 558860
rect 79501 558859 79567 558862
rect 80646 558860 80652 558862
rect 80716 558860 80763 558864
rect 80697 558859 80763 558860
rect 81433 558922 81499 558925
rect 82905 558924 82971 558925
rect 82118 558922 82124 558924
rect 81433 558920 82124 558922
rect 81433 558864 81438 558920
rect 81494 558864 82124 558920
rect 81433 558862 82124 558864
rect 81433 558859 81499 558862
rect 82118 558860 82124 558862
rect 82188 558860 82194 558924
rect 82854 558922 82860 558924
rect 82814 558862 82860 558922
rect 82924 558920 82971 558924
rect 82966 558864 82971 558920
rect 82854 558860 82860 558862
rect 82924 558860 82971 558864
rect 82905 558859 82971 558860
rect 84193 558922 84259 558925
rect 85389 558924 85455 558925
rect 85665 558924 85731 558925
rect 84694 558922 84700 558924
rect 84193 558920 84700 558922
rect 84193 558864 84198 558920
rect 84254 558864 84700 558920
rect 84193 558862 84700 558864
rect 84193 558859 84259 558862
rect 84694 558860 84700 558862
rect 84764 558860 84770 558924
rect 85389 558920 85436 558924
rect 85500 558922 85506 558924
rect 85389 558864 85394 558920
rect 85389 558860 85436 558864
rect 85500 558862 85546 558922
rect 85500 558860 85506 558862
rect 85614 558860 85620 558924
rect 85684 558922 85731 558924
rect 86217 558922 86283 558925
rect 86718 558922 86724 558924
rect 85684 558920 85776 558922
rect 85726 558864 85776 558920
rect 85684 558862 85776 558864
rect 86217 558920 86724 558922
rect 86217 558864 86222 558920
rect 86278 558864 86724 558920
rect 86217 558862 86724 558864
rect 85684 558860 85731 558862
rect 85389 558859 85455 558860
rect 85665 558859 85731 558860
rect 86217 558859 86283 558862
rect 86718 558860 86724 558862
rect 86788 558860 86794 558924
rect 87597 558922 87663 558925
rect 88977 558924 89043 558925
rect 88190 558922 88196 558924
rect 87597 558920 88196 558922
rect 87597 558864 87602 558920
rect 87658 558864 88196 558920
rect 87597 558862 88196 558864
rect 87597 558859 87663 558862
rect 88190 558860 88196 558862
rect 88260 558860 88266 558924
rect 88926 558922 88932 558924
rect 88886 558862 88932 558922
rect 88996 558920 89043 558924
rect 89038 558864 89043 558920
rect 88926 558860 88932 558862
rect 88996 558860 89043 558864
rect 89110 558860 89116 558924
rect 89180 558922 89186 558924
rect 89621 558922 89687 558925
rect 90081 558924 90147 558925
rect 91369 558924 91435 558925
rect 92473 558924 92539 558925
rect 93577 558924 93643 558925
rect 90030 558922 90036 558924
rect 89180 558920 89687 558922
rect 89180 558864 89626 558920
rect 89682 558864 89687 558920
rect 89180 558862 89687 558864
rect 89990 558862 90036 558922
rect 90100 558920 90147 558924
rect 91318 558922 91324 558924
rect 90142 558864 90147 558920
rect 89180 558860 89186 558862
rect 88977 558859 89043 558860
rect 89621 558859 89687 558862
rect 90030 558860 90036 558862
rect 90100 558860 90147 558864
rect 91278 558862 91324 558922
rect 91388 558920 91435 558924
rect 92422 558922 92428 558924
rect 91430 558864 91435 558920
rect 91318 558860 91324 558862
rect 91388 558860 91435 558864
rect 92382 558862 92428 558922
rect 92492 558920 92539 558924
rect 93526 558922 93532 558924
rect 92534 558864 92539 558920
rect 92422 558860 92428 558862
rect 92492 558860 92539 558864
rect 93486 558862 93532 558922
rect 93596 558920 93643 558924
rect 93638 558864 93643 558920
rect 93526 558860 93532 558862
rect 93596 558860 93643 558864
rect 90081 558859 90147 558860
rect 91369 558859 91435 558860
rect 92473 558859 92539 558860
rect 93577 558859 93643 558860
rect 94589 558924 94655 558925
rect 95325 558924 95391 558925
rect 96613 558924 96679 558925
rect 98269 558924 98335 558925
rect 99557 558924 99623 558925
rect 94589 558920 94636 558924
rect 94700 558922 94706 558924
rect 94589 558864 94594 558920
rect 94589 558860 94636 558864
rect 94700 558862 94746 558922
rect 95325 558920 95372 558924
rect 95436 558922 95442 558924
rect 95325 558864 95330 558920
rect 94700 558860 94706 558862
rect 95325 558860 95372 558864
rect 95436 558862 95482 558922
rect 96613 558920 96660 558924
rect 96724 558922 96730 558924
rect 96613 558864 96618 558920
rect 95436 558860 95442 558862
rect 96613 558860 96660 558864
rect 96724 558862 96770 558922
rect 98269 558920 98316 558924
rect 98380 558922 98386 558924
rect 98269 558864 98274 558920
rect 96724 558860 96730 558862
rect 98269 558860 98316 558864
rect 98380 558862 98426 558922
rect 99557 558920 99604 558924
rect 99668 558922 99674 558924
rect 99557 558864 99562 558920
rect 98380 558860 98386 558862
rect 99557 558860 99604 558864
rect 99668 558862 99714 558922
rect 99668 558860 99674 558862
rect 100150 558860 100156 558924
rect 100220 558922 100226 558924
rect 100661 558922 100727 558925
rect 101949 558924 102015 558925
rect 102685 558924 102751 558925
rect 101949 558922 101996 558924
rect 100220 558920 100727 558922
rect 100220 558864 100666 558920
rect 100722 558864 100727 558920
rect 100220 558862 100727 558864
rect 101904 558920 101996 558922
rect 101904 558864 101954 558920
rect 101904 558862 101996 558864
rect 100220 558860 100226 558862
rect 94589 558859 94655 558860
rect 95325 558859 95391 558860
rect 96613 558859 96679 558860
rect 98269 558859 98335 558860
rect 99557 558859 99623 558860
rect 100661 558859 100727 558862
rect 101949 558860 101996 558862
rect 102060 558860 102066 558924
rect 102685 558920 102732 558924
rect 102796 558922 102802 558924
rect 102685 558864 102690 558920
rect 102685 558860 102732 558864
rect 102796 558862 102842 558922
rect 102796 558860 102802 558862
rect 103278 558860 103284 558924
rect 103348 558922 103354 558924
rect 103421 558922 103487 558925
rect 103348 558920 103487 558922
rect 103348 558864 103426 558920
rect 103482 558864 103487 558920
rect 103348 558862 103487 558864
rect 103348 558860 103354 558862
rect 101949 558859 102015 558860
rect 102685 558859 102751 558860
rect 103421 558859 103487 558862
rect 103973 558924 104039 558925
rect 104801 558924 104867 558925
rect 105353 558924 105419 558925
rect 103973 558920 104020 558924
rect 104084 558922 104090 558924
rect 103973 558864 103978 558920
rect 103973 558860 104020 558864
rect 104084 558862 104130 558922
rect 104084 558860 104090 558862
rect 104750 558860 104756 558924
rect 104820 558922 104867 558924
rect 105302 558922 105308 558924
rect 104820 558920 104912 558922
rect 104862 558864 104912 558920
rect 104820 558862 104912 558864
rect 105262 558862 105308 558922
rect 105372 558920 105419 558924
rect 105414 558864 105419 558920
rect 104820 558860 104867 558862
rect 105302 558860 105308 558862
rect 105372 558860 105419 558864
rect 106038 558860 106044 558924
rect 106108 558922 106114 558924
rect 106181 558922 106247 558925
rect 106108 558920 106247 558922
rect 106108 558864 106186 558920
rect 106242 558864 106247 558920
rect 106108 558862 106247 558864
rect 106108 558860 106114 558862
rect 103973 558859 104039 558860
rect 104801 558859 104867 558860
rect 105353 558859 105419 558860
rect 106181 558859 106247 558862
rect 107142 558860 107148 558924
rect 107212 558922 107218 558924
rect 107561 558922 107627 558925
rect 107212 558920 107627 558922
rect 107212 558864 107566 558920
rect 107622 558864 107627 558920
rect 107212 558862 107627 558864
rect 107212 558860 107218 558862
rect 107561 558859 107627 558862
rect 107694 558860 107700 558924
rect 107764 558922 107770 558924
rect 107837 558922 107903 558925
rect 107764 558920 107903 558922
rect 107764 558864 107842 558920
rect 107898 558864 107903 558920
rect 107764 558862 107903 558864
rect 107764 558860 107770 558862
rect 107837 558859 107903 558862
rect 108430 558860 108436 558924
rect 108500 558922 108506 558924
rect 108941 558922 109007 558925
rect 108500 558920 109007 558922
rect 108500 558864 108946 558920
rect 109002 558864 109007 558920
rect 108500 558862 109007 558864
rect 108500 558860 108506 558862
rect 108941 558859 109007 558862
rect 109534 558860 109540 558924
rect 109604 558922 109610 558924
rect 110321 558922 110387 558925
rect 109604 558920 110387 558922
rect 109604 558864 110326 558920
rect 110382 558864 110387 558920
rect 109604 558862 110387 558864
rect 109604 558860 109610 558862
rect 110321 558859 110387 558862
rect 193765 558924 193831 558925
rect 193765 558920 193812 558924
rect 193876 558922 193882 558924
rect 193765 558864 193770 558920
rect 193765 558860 193812 558864
rect 193876 558862 193922 558922
rect 193876 558860 193882 558862
rect 202638 558860 202644 558924
rect 202708 558922 202714 558924
rect 202781 558922 202847 558925
rect 202708 558920 202847 558922
rect 202708 558864 202786 558920
rect 202842 558864 202847 558920
rect 202708 558862 202847 558864
rect 202708 558860 202714 558862
rect 193765 558859 193831 558860
rect 202781 558859 202847 558862
rect 203926 558860 203932 558924
rect 203996 558922 204002 558924
rect 204161 558922 204227 558925
rect 203996 558920 204227 558922
rect 203996 558864 204166 558920
rect 204222 558864 204227 558920
rect 203996 558862 204227 558864
rect 203996 558860 204002 558862
rect 204161 558859 204227 558862
rect 205398 558860 205404 558924
rect 205468 558922 205474 558924
rect 205541 558922 205607 558925
rect 211889 558924 211955 558925
rect 213177 558924 213243 558925
rect 211838 558922 211844 558924
rect 205468 558920 205607 558922
rect 205468 558864 205546 558920
rect 205602 558864 205607 558920
rect 205468 558862 205607 558864
rect 211798 558862 211844 558922
rect 211908 558920 211955 558924
rect 213126 558922 213132 558924
rect 211950 558864 211955 558920
rect 205468 558860 205474 558862
rect 205541 558859 205607 558862
rect 211838 558860 211844 558862
rect 211908 558860 211955 558864
rect 213086 558862 213132 558922
rect 213196 558920 213243 558924
rect 213238 558864 213243 558920
rect 213126 558860 213132 558862
rect 213196 558860 213243 558864
rect 211889 558859 211955 558860
rect 213177 558859 213243 558860
rect 213913 558922 213979 558925
rect 214046 558922 214052 558924
rect 213913 558920 214052 558922
rect 213913 558864 213918 558920
rect 213974 558864 214052 558920
rect 213913 558862 214052 558864
rect 213913 558859 213979 558862
rect 214046 558860 214052 558862
rect 214116 558860 214122 558924
rect 216254 558860 216260 558924
rect 216324 558922 216330 558924
rect 216581 558922 216647 558925
rect 217593 558924 217659 558925
rect 217542 558922 217548 558924
rect 216324 558920 216647 558922
rect 216324 558864 216586 558920
rect 216642 558864 216647 558920
rect 216324 558862 216647 558864
rect 217502 558862 217548 558922
rect 217612 558920 217659 558924
rect 217869 558924 217935 558925
rect 218881 558924 218947 558925
rect 217869 558922 217916 558924
rect 217654 558864 217659 558920
rect 216324 558860 216330 558862
rect 216581 558859 216647 558862
rect 217542 558860 217548 558862
rect 217612 558860 217659 558864
rect 217824 558920 217916 558922
rect 217824 558864 217874 558920
rect 217824 558862 217916 558864
rect 217593 558859 217659 558860
rect 217869 558860 217916 558862
rect 217980 558860 217986 558924
rect 218830 558922 218836 558924
rect 218790 558862 218836 558922
rect 218900 558920 218947 558924
rect 218942 558864 218947 558920
rect 218830 558860 218836 558862
rect 218900 558860 218947 558864
rect 219198 558860 219204 558924
rect 219268 558922 219274 558924
rect 219341 558922 219407 558925
rect 219268 558920 219407 558922
rect 219268 558864 219346 558920
rect 219402 558864 219407 558920
rect 219268 558862 219407 558864
rect 219268 558860 219274 558862
rect 217869 558859 217935 558860
rect 218881 558859 218947 558860
rect 219341 558859 219407 558862
rect 220077 558924 220143 558925
rect 220721 558924 220787 558925
rect 221089 558924 221155 558925
rect 220077 558920 220124 558924
rect 220188 558922 220194 558924
rect 220077 558864 220082 558920
rect 220077 558860 220124 558864
rect 220188 558862 220234 558922
rect 220188 558860 220194 558862
rect 220670 558860 220676 558924
rect 220740 558922 220787 558924
rect 221038 558922 221044 558924
rect 220740 558920 220832 558922
rect 220782 558864 220832 558920
rect 220740 558862 220832 558864
rect 220998 558862 221044 558922
rect 221108 558920 221155 558924
rect 221150 558864 221155 558920
rect 220740 558860 220787 558862
rect 221038 558860 221044 558862
rect 221108 558860 221155 558864
rect 221958 558860 221964 558924
rect 222028 558922 222034 558924
rect 222101 558922 222167 558925
rect 222028 558920 222167 558922
rect 222028 558864 222106 558920
rect 222162 558864 222167 558920
rect 222028 558862 222167 558864
rect 222028 558860 222034 558862
rect 220077 558859 220143 558860
rect 220721 558859 220787 558860
rect 221089 558859 221155 558860
rect 222101 558859 222167 558862
rect 222285 558924 222351 558925
rect 222285 558920 222332 558924
rect 222396 558922 222402 558924
rect 222285 558864 222290 558920
rect 222285 558860 222332 558864
rect 222396 558862 222442 558922
rect 222396 558860 222402 558862
rect 223246 558860 223252 558924
rect 223316 558922 223322 558924
rect 223481 558922 223547 558925
rect 223316 558920 223547 558922
rect 223316 558864 223486 558920
rect 223542 558864 223547 558920
rect 223316 558862 223547 558864
rect 223316 558860 223322 558862
rect 222285 558859 222351 558860
rect 223481 558859 223547 558862
rect 224350 558860 224356 558924
rect 224420 558922 224426 558924
rect 224861 558922 224927 558925
rect 224420 558920 224927 558922
rect 224420 558864 224866 558920
rect 224922 558864 224927 558920
rect 224420 558862 224927 558864
rect 224420 558860 224426 558862
rect 224861 558859 224927 558862
rect 225781 558924 225847 558925
rect 226241 558924 226307 558925
rect 227161 558924 227227 558925
rect 225781 558920 225828 558924
rect 225892 558922 225898 558924
rect 225781 558864 225786 558920
rect 225781 558860 225828 558864
rect 225892 558862 225938 558922
rect 225892 558860 225898 558862
rect 226190 558860 226196 558924
rect 226260 558922 226307 558924
rect 227110 558922 227116 558924
rect 226260 558920 226352 558922
rect 226302 558864 226352 558920
rect 226260 558862 226352 558864
rect 227070 558862 227116 558922
rect 227180 558920 227227 558924
rect 227222 558864 227227 558920
rect 226260 558860 226307 558862
rect 227110 558860 227116 558862
rect 227180 558860 227227 558864
rect 227478 558860 227484 558924
rect 227548 558922 227554 558924
rect 227621 558922 227687 558925
rect 227548 558920 227687 558922
rect 227548 558864 227626 558920
rect 227682 558864 227687 558920
rect 227548 558862 227687 558864
rect 227548 558860 227554 558862
rect 225781 558859 225847 558860
rect 226241 558859 226307 558860
rect 227161 558859 227227 558860
rect 227621 558859 227687 558862
rect 228766 558860 228772 558924
rect 228836 558922 228842 558924
rect 229001 558922 229067 558925
rect 228836 558920 229067 558922
rect 228836 558864 229006 558920
rect 229062 558864 229067 558920
rect 228836 558862 229067 558864
rect 228836 558860 228842 558862
rect 229001 558859 229067 558862
rect 229461 558924 229527 558925
rect 229461 558920 229508 558924
rect 229572 558922 229578 558924
rect 229461 558864 229466 558920
rect 229461 558860 229508 558864
rect 229572 558862 229618 558922
rect 229572 558860 229578 558862
rect 230238 558860 230244 558924
rect 230308 558922 230314 558924
rect 230381 558922 230447 558925
rect 230308 558920 230447 558922
rect 230308 558864 230386 558920
rect 230442 558864 230447 558920
rect 230308 558862 230447 558864
rect 230308 558860 230314 558862
rect 229461 558859 229527 558860
rect 230381 558859 230447 558862
rect 230790 558860 230796 558924
rect 230860 558922 230866 558924
rect 231761 558922 231827 558925
rect 230860 558920 231827 558922
rect 230860 558864 231766 558920
rect 231822 558864 231827 558920
rect 230860 558862 231827 558864
rect 230860 558860 230866 558862
rect 231761 558859 231827 558862
rect 231945 558922 232011 558925
rect 232814 558922 232820 558924
rect 231945 558920 232820 558922
rect 231945 558864 231950 558920
rect 232006 558864 232820 558920
rect 231945 558862 232820 558864
rect 231945 558859 232011 558862
rect 232814 558860 232820 558862
rect 232884 558860 232890 558924
rect 232998 558860 233004 558924
rect 233068 558922 233074 558924
rect 233141 558922 233207 558925
rect 234521 558924 234587 558925
rect 233068 558920 233207 558922
rect 233068 558864 233146 558920
rect 233202 558864 233207 558920
rect 233068 558862 233207 558864
rect 233068 558860 233074 558862
rect 233141 558859 233207 558862
rect 234470 558860 234476 558924
rect 234540 558922 234587 558924
rect 234540 558920 234632 558922
rect 234582 558864 234632 558920
rect 234540 558862 234632 558864
rect 234540 558860 234587 558862
rect 235758 558860 235764 558924
rect 235828 558922 235834 558924
rect 235901 558922 235967 558925
rect 237281 558924 237347 558925
rect 235828 558920 235967 558922
rect 235828 558864 235906 558920
rect 235962 558864 235967 558920
rect 235828 558862 235967 558864
rect 235828 558860 235834 558862
rect 234521 558859 234587 558860
rect 235901 558859 235967 558862
rect 237230 558860 237236 558924
rect 237300 558922 237347 558924
rect 237300 558920 237392 558922
rect 237342 558864 237392 558920
rect 237300 558862 237392 558864
rect 237300 558860 237347 558862
rect 239622 558860 239628 558924
rect 239692 558922 239698 558924
rect 240041 558922 240107 558925
rect 239692 558920 240107 558922
rect 239692 558864 240046 558920
rect 240102 558864 240107 558920
rect 239692 558862 240107 558864
rect 239692 558860 239698 558862
rect 237281 558859 237347 558860
rect 240041 558859 240107 558862
rect 313733 558924 313799 558925
rect 313733 558920 313780 558924
rect 313844 558922 313850 558924
rect 316033 558922 316099 558925
rect 316166 558922 316172 558924
rect 313733 558864 313738 558920
rect 313733 558860 313780 558864
rect 313844 558862 313890 558922
rect 316033 558920 316172 558922
rect 316033 558864 316038 558920
rect 316094 558864 316172 558920
rect 316033 558862 316172 558864
rect 313844 558860 313850 558862
rect 313733 558859 313799 558860
rect 316033 558859 316099 558862
rect 316166 558860 316172 558862
rect 316236 558860 316242 558924
rect 318793 558922 318859 558925
rect 318926 558922 318932 558924
rect 318793 558920 318932 558922
rect 318793 558864 318798 558920
rect 318854 558864 318932 558920
rect 318793 558862 318932 558864
rect 318793 558859 318859 558862
rect 318926 558860 318932 558862
rect 318996 558860 319002 558924
rect 320265 558922 320331 558925
rect 320950 558922 320956 558924
rect 320265 558920 320956 558922
rect 320265 558864 320270 558920
rect 320326 558864 320956 558920
rect 320265 558862 320956 558864
rect 320265 558859 320331 558862
rect 320950 558860 320956 558862
rect 321020 558860 321026 558924
rect 321553 558922 321619 558925
rect 322790 558922 322796 558924
rect 321553 558920 322796 558922
rect 321553 558864 321558 558920
rect 321614 558864 322796 558920
rect 321553 558862 322796 558864
rect 321553 558859 321619 558862
rect 322790 558860 322796 558862
rect 322860 558860 322866 558924
rect 323577 558922 323643 558925
rect 325182 558922 325188 558924
rect 323577 558920 325188 558922
rect 323577 558864 323582 558920
rect 323638 558864 325188 558920
rect 323577 558862 325188 558864
rect 323577 558859 323643 558862
rect 325182 558860 325188 558862
rect 325252 558860 325258 558924
rect 325693 558922 325759 558925
rect 326286 558922 326292 558924
rect 325693 558920 326292 558922
rect 325693 558864 325698 558920
rect 325754 558864 326292 558920
rect 325693 558862 326292 558864
rect 325693 558859 325759 558862
rect 326286 558860 326292 558862
rect 326356 558860 326362 558924
rect 327073 558922 327139 558925
rect 327574 558922 327580 558924
rect 327073 558920 327580 558922
rect 327073 558864 327078 558920
rect 327134 558864 327580 558920
rect 327073 558862 327580 558864
rect 327073 558859 327139 558862
rect 327574 558860 327580 558862
rect 327644 558860 327650 558924
rect 329925 558922 329991 558925
rect 331765 558924 331831 558925
rect 331070 558922 331076 558924
rect 329925 558920 331076 558922
rect 329925 558864 329930 558920
rect 329986 558864 331076 558920
rect 329925 558862 331076 558864
rect 329925 558859 329991 558862
rect 331070 558860 331076 558862
rect 331140 558860 331146 558924
rect 331765 558920 331812 558924
rect 331876 558922 331882 558924
rect 332593 558922 332659 558925
rect 333278 558922 333284 558924
rect 331765 558864 331770 558920
rect 331765 558860 331812 558864
rect 331876 558862 331922 558922
rect 332593 558920 333284 558922
rect 332593 558864 332598 558920
rect 332654 558864 333284 558920
rect 332593 558862 333284 558864
rect 331876 558860 331882 558862
rect 331765 558859 331831 558860
rect 332593 558859 332659 558862
rect 333278 558860 333284 558862
rect 333348 558860 333354 558924
rect 333973 558922 334039 558925
rect 334566 558922 334572 558924
rect 333973 558920 334572 558922
rect 333973 558864 333978 558920
rect 334034 558864 334572 558920
rect 333973 558862 334572 558864
rect 333973 558859 334039 558862
rect 334566 558860 334572 558862
rect 334636 558860 334642 558924
rect 335353 558922 335419 558925
rect 336733 558924 336799 558925
rect 335854 558922 335860 558924
rect 335353 558920 335860 558922
rect 335353 558864 335358 558920
rect 335414 558864 335860 558920
rect 335353 558862 335860 558864
rect 335353 558859 335419 558862
rect 335854 558860 335860 558862
rect 335924 558860 335930 558924
rect 336733 558922 336780 558924
rect 336688 558920 336780 558922
rect 336688 558864 336738 558920
rect 336688 558862 336780 558864
rect 336733 558860 336780 558862
rect 336844 558860 336850 558924
rect 337377 558922 337443 558925
rect 337694 558922 337700 558924
rect 337377 558920 337700 558922
rect 337377 558864 337382 558920
rect 337438 558864 337700 558920
rect 337377 558862 337700 558864
rect 336733 558859 336799 558860
rect 337377 558859 337443 558862
rect 337694 558860 337700 558862
rect 337764 558860 337770 558924
rect 338113 558922 338179 558925
rect 339166 558922 339172 558924
rect 338113 558920 339172 558922
rect 338113 558864 338118 558920
rect 338174 558864 339172 558920
rect 338113 558862 339172 558864
rect 338113 558859 338179 558862
rect 339166 558860 339172 558862
rect 339236 558860 339242 558924
rect 339493 558922 339559 558925
rect 340454 558922 340460 558924
rect 339493 558920 340460 558922
rect 339493 558864 339498 558920
rect 339554 558864 340460 558920
rect 339493 558862 340460 558864
rect 339493 558859 339559 558862
rect 340454 558860 340460 558862
rect 340524 558860 340530 558924
rect 340873 558922 340939 558925
rect 341742 558922 341748 558924
rect 340873 558920 341748 558922
rect 340873 558864 340878 558920
rect 340934 558864 341748 558920
rect 340873 558862 341748 558864
rect 340873 558859 340939 558862
rect 341742 558860 341748 558862
rect 341812 558860 341818 558924
rect 342253 558922 342319 558925
rect 342662 558922 342668 558924
rect 342253 558920 342668 558922
rect 342253 558864 342258 558920
rect 342314 558864 342668 558920
rect 342253 558862 342668 558864
rect 342253 558859 342319 558862
rect 342662 558860 342668 558862
rect 342732 558860 342738 558924
rect 343633 558922 343699 558925
rect 344277 558924 344343 558925
rect 343950 558922 343956 558924
rect 343633 558920 343956 558922
rect 343633 558864 343638 558920
rect 343694 558864 343956 558920
rect 343633 558862 343956 558864
rect 343633 558859 343699 558862
rect 343950 558860 343956 558862
rect 344020 558860 344026 558924
rect 344277 558920 344324 558924
rect 344388 558922 344394 558924
rect 345013 558922 345079 558925
rect 346158 558922 346164 558924
rect 344277 558864 344282 558920
rect 344277 558860 344324 558864
rect 344388 558862 344434 558922
rect 345013 558920 346164 558922
rect 345013 558864 345018 558920
rect 345074 558864 346164 558920
rect 345013 558862 346164 558864
rect 344388 558860 344394 558862
rect 344277 558859 344343 558860
rect 345013 558859 345079 558862
rect 346158 558860 346164 558862
rect 346228 558860 346234 558924
rect 346393 558922 346459 558925
rect 347446 558922 347452 558924
rect 346393 558920 347452 558922
rect 346393 558864 346398 558920
rect 346454 558864 347452 558920
rect 346393 558862 347452 558864
rect 346393 558859 346459 558862
rect 347446 558860 347452 558862
rect 347516 558860 347522 558924
rect 347773 558922 347839 558925
rect 348734 558922 348740 558924
rect 347773 558920 348740 558922
rect 347773 558864 347778 558920
rect 347834 558864 348740 558920
rect 347773 558862 348740 558864
rect 347773 558859 347839 558862
rect 348734 558860 348740 558862
rect 348804 558860 348810 558924
rect 349153 558922 349219 558925
rect 349654 558922 349660 558924
rect 349153 558920 349660 558922
rect 349153 558864 349158 558920
rect 349214 558864 349660 558920
rect 349153 558862 349660 558864
rect 349153 558859 349219 558862
rect 349654 558860 349660 558862
rect 349724 558860 349730 558924
rect 351913 558922 351979 558925
rect 443085 558924 443151 558925
rect 352414 558922 352420 558924
rect 351913 558920 352420 558922
rect 351913 558864 351918 558920
rect 351974 558864 352420 558920
rect 351913 558862 352420 558864
rect 351913 558859 351979 558862
rect 352414 558860 352420 558862
rect 352484 558860 352490 558924
rect 443085 558920 443132 558924
rect 443196 558922 443202 558924
rect 445753 558922 445819 558925
rect 446254 558922 446260 558924
rect 443085 558864 443090 558920
rect 443085 558860 443132 558864
rect 443196 558862 443242 558922
rect 445753 558920 446260 558922
rect 445753 558864 445758 558920
rect 445814 558864 446260 558920
rect 445753 558862 446260 558864
rect 443196 558860 443202 558862
rect 443085 558859 443151 558860
rect 445753 558859 445819 558862
rect 446254 558860 446260 558862
rect 446324 558860 446330 558924
rect 446397 558922 446463 558925
rect 447358 558922 447364 558924
rect 446397 558920 447364 558922
rect 446397 558864 446402 558920
rect 446458 558864 447364 558920
rect 446397 558862 447364 558864
rect 446397 558859 446463 558862
rect 447358 558860 447364 558862
rect 447428 558860 447434 558924
rect 447777 558922 447843 558925
rect 448462 558922 448468 558924
rect 447777 558920 448468 558922
rect 447777 558864 447782 558920
rect 447838 558864 448468 558920
rect 447777 558862 448468 558864
rect 447777 558859 447843 558862
rect 448462 558860 448468 558862
rect 448532 558860 448538 558924
rect 449157 558922 449223 558925
rect 449934 558922 449940 558924
rect 449157 558920 449940 558922
rect 449157 558864 449162 558920
rect 449218 558864 449940 558920
rect 449157 558862 449940 558864
rect 449157 558859 449223 558862
rect 449934 558860 449940 558862
rect 450004 558860 450010 558924
rect 452745 558922 452811 558925
rect 452878 558922 452884 558924
rect 452745 558920 452884 558922
rect 452745 558864 452750 558920
rect 452806 558864 452884 558920
rect 452745 558862 452884 558864
rect 452745 558859 452811 558862
rect 452878 558860 452884 558862
rect 452948 558860 452954 558924
rect 453481 558922 453547 558925
rect 454677 558924 454743 558925
rect 453614 558922 453620 558924
rect 453481 558920 453620 558922
rect 453481 558864 453486 558920
rect 453542 558864 453620 558920
rect 453481 558862 453620 558864
rect 453481 558859 453547 558862
rect 453614 558860 453620 558862
rect 453684 558860 453690 558924
rect 454677 558920 454724 558924
rect 454788 558922 454794 558924
rect 454677 558864 454682 558920
rect 454677 558860 454724 558864
rect 454788 558862 454834 558922
rect 454788 558860 454794 558862
rect 458398 558860 458404 558924
rect 458468 558922 458474 558924
rect 458817 558922 458883 558925
rect 458468 558920 458883 558922
rect 458468 558864 458822 558920
rect 458878 558864 458883 558920
rect 458468 558862 458883 558864
rect 458468 558860 458474 558862
rect 454677 558859 454743 558860
rect 458817 558859 458883 558862
rect 460933 558924 460999 558925
rect 461761 558924 461827 558925
rect 460933 558920 460980 558924
rect 461044 558922 461050 558924
rect 461710 558922 461716 558924
rect 460933 558864 460938 558920
rect 460933 558860 460980 558864
rect 461044 558862 461090 558922
rect 461670 558862 461716 558922
rect 461780 558920 461827 558924
rect 461822 558864 461827 558920
rect 461044 558860 461050 558862
rect 461710 558860 461716 558862
rect 461780 558860 461827 558864
rect 460933 558859 460999 558860
rect 461761 558859 461827 558860
rect 462313 558922 462379 558925
rect 463366 558922 463372 558924
rect 462313 558920 463372 558922
rect 462313 558864 462318 558920
rect 462374 558864 463372 558920
rect 462313 558862 463372 558864
rect 462313 558859 462379 558862
rect 463366 558860 463372 558862
rect 463436 558860 463442 558924
rect 463693 558922 463759 558925
rect 464470 558922 464476 558924
rect 463693 558920 464476 558922
rect 463693 558864 463698 558920
rect 463754 558864 464476 558920
rect 463693 558862 464476 558864
rect 463693 558859 463759 558862
rect 464470 558860 464476 558862
rect 464540 558860 464546 558924
rect 465073 558922 465139 558925
rect 465758 558922 465764 558924
rect 465073 558920 465764 558922
rect 465073 558864 465078 558920
rect 465134 558864 465764 558920
rect 465073 558862 465764 558864
rect 465073 558859 465139 558862
rect 465758 558860 465764 558862
rect 465828 558860 465834 558924
rect 466453 558922 466519 558925
rect 466862 558922 466868 558924
rect 466453 558920 466868 558922
rect 466453 558864 466458 558920
rect 466514 558864 466868 558920
rect 466453 558862 466868 558864
rect 466453 558859 466519 558862
rect 466862 558860 466868 558862
rect 466932 558860 466938 558924
rect 467833 558922 467899 558925
rect 467966 558922 467972 558924
rect 467833 558920 467972 558922
rect 467833 558864 467838 558920
rect 467894 558864 467972 558920
rect 467833 558862 467972 558864
rect 467833 558859 467899 558862
rect 467966 558860 467972 558862
rect 468036 558860 468042 558924
rect 468569 558922 468635 558925
rect 468702 558922 468708 558924
rect 468569 558920 468708 558922
rect 468569 558864 468574 558920
rect 468630 558864 468708 558920
rect 468569 558862 468708 558864
rect 468569 558859 468635 558862
rect 468702 558860 468708 558862
rect 468772 558860 468778 558924
rect 469213 558922 469279 558925
rect 470358 558922 470364 558924
rect 469213 558920 470364 558922
rect 469213 558864 469218 558920
rect 469274 558864 470364 558920
rect 469213 558862 470364 558864
rect 469213 558859 469279 558862
rect 470358 558860 470364 558862
rect 470428 558860 470434 558924
rect 470593 558922 470659 558925
rect 471462 558922 471468 558924
rect 470593 558920 471468 558922
rect 470593 558864 470598 558920
rect 470654 558864 471468 558920
rect 470593 558862 471468 558864
rect 470593 558859 470659 558862
rect 471462 558860 471468 558862
rect 471532 558860 471538 558924
rect 471973 558922 472039 558925
rect 472750 558922 472756 558924
rect 471973 558920 472756 558922
rect 471973 558864 471978 558920
rect 472034 558864 472756 558920
rect 471973 558862 472756 558864
rect 471973 558859 472039 558862
rect 472750 558860 472756 558862
rect 472820 558860 472826 558924
rect 473353 558922 473419 558925
rect 474038 558922 474044 558924
rect 473353 558920 474044 558922
rect 473353 558864 473358 558920
rect 473414 558864 474044 558920
rect 473353 558862 474044 558864
rect 473353 558859 473419 558862
rect 474038 558860 474044 558862
rect 474108 558860 474114 558924
rect 474733 558922 474799 558925
rect 476205 558924 476271 558925
rect 477125 558924 477191 558925
rect 478321 558924 478387 558925
rect 479425 558924 479491 558925
rect 474958 558922 474964 558924
rect 474733 558920 474964 558922
rect 474733 558864 474738 558920
rect 474794 558864 474964 558920
rect 474733 558862 474964 558864
rect 474733 558859 474799 558862
rect 474958 558860 474964 558862
rect 475028 558860 475034 558924
rect 476205 558922 476252 558924
rect 476160 558920 476252 558922
rect 476160 558864 476210 558920
rect 476160 558862 476252 558864
rect 476205 558860 476252 558862
rect 476316 558860 476322 558924
rect 477125 558920 477172 558924
rect 477236 558922 477242 558924
rect 478270 558922 478276 558924
rect 477125 558864 477130 558920
rect 477125 558860 477172 558864
rect 477236 558862 477282 558922
rect 478230 558862 478276 558922
rect 478340 558920 478387 558924
rect 479374 558922 479380 558924
rect 478382 558864 478387 558920
rect 477236 558860 477242 558862
rect 478270 558860 478276 558862
rect 478340 558860 478387 558864
rect 479334 558862 479380 558922
rect 479444 558920 479491 558924
rect 479486 558864 479491 558920
rect 479374 558860 479380 558862
rect 479444 558860 479491 558864
rect 476205 558859 476271 558860
rect 477125 558859 477191 558860
rect 478321 558859 478387 558860
rect 479425 558859 479491 558860
rect 480529 558922 480595 558925
rect 480846 558922 480852 558924
rect 480529 558920 480852 558922
rect 480529 558864 480534 558920
rect 480590 558864 480852 558920
rect 480529 558862 480852 558864
rect 480529 558859 480595 558862
rect 480846 558860 480852 558862
rect 480916 558860 480922 558924
rect 483013 558922 483079 558925
rect 483422 558922 483428 558924
rect 483013 558920 483428 558922
rect 483013 558864 483018 558920
rect 483074 558864 483428 558920
rect 483013 558862 483428 558864
rect 483013 558859 483079 558862
rect 483422 558860 483428 558862
rect 483492 558860 483498 558924
rect 484485 558922 484551 558925
rect 485630 558922 485636 558924
rect 484485 558920 485636 558922
rect 484485 558864 484490 558920
rect 484546 558864 485636 558920
rect 484485 558862 485636 558864
rect 484485 558859 484551 558862
rect 485630 558860 485636 558862
rect 485700 558860 485706 558924
rect 485773 558922 485839 558925
rect 485998 558922 486004 558924
rect 485773 558920 486004 558922
rect 485773 558864 485778 558920
rect 485834 558864 486004 558920
rect 485773 558862 486004 558864
rect 485773 558859 485839 558862
rect 485998 558860 486004 558862
rect 486068 558860 486074 558924
rect 61694 558724 61700 558788
rect 61764 558786 61770 558788
rect 63534 558786 63540 558788
rect 61764 558726 63540 558786
rect 61764 558724 61770 558726
rect 63534 558724 63540 558726
rect 63604 558786 63610 558788
rect 64321 558786 64387 558789
rect 70209 558788 70275 558789
rect 63604 558784 64387 558786
rect 63604 558728 64326 558784
rect 64382 558728 64387 558784
rect 63604 558726 64387 558728
rect 63604 558724 63610 558726
rect 64321 558723 64387 558726
rect 70158 558724 70164 558788
rect 70228 558786 70275 558788
rect 80053 558786 80119 558789
rect 81014 558786 81020 558788
rect 70228 558784 70320 558786
rect 70270 558728 70320 558784
rect 70228 558726 70320 558728
rect 80053 558784 81020 558786
rect 80053 558728 80058 558784
rect 80114 558728 81020 558784
rect 80053 558726 81020 558728
rect 70228 558724 70275 558726
rect 70209 558723 70275 558724
rect 80053 558723 80119 558726
rect 81014 558724 81020 558726
rect 81084 558724 81090 558788
rect 81617 558786 81683 558789
rect 81750 558786 81756 558788
rect 81617 558784 81756 558786
rect 81617 558728 81622 558784
rect 81678 558728 81756 558784
rect 81617 558726 81756 558728
rect 81617 558723 81683 558726
rect 81750 558724 81756 558726
rect 81820 558724 81826 558788
rect 84142 558724 84148 558788
rect 84212 558786 84218 558788
rect 84285 558786 84351 558789
rect 84212 558784 84351 558786
rect 84212 558728 84290 558784
rect 84346 558728 84351 558784
rect 84212 558726 84351 558728
rect 84212 558724 84218 558726
rect 84285 558723 84351 558726
rect 86350 558724 86356 558788
rect 86420 558786 86426 558788
rect 86861 558786 86927 558789
rect 87873 558788 87939 558789
rect 87822 558786 87828 558788
rect 86420 558784 86927 558786
rect 86420 558728 86866 558784
rect 86922 558728 86927 558784
rect 86420 558726 86927 558728
rect 87782 558726 87828 558786
rect 87892 558784 87939 558788
rect 87934 558728 87939 558784
rect 86420 558724 86426 558726
rect 86861 558723 86927 558726
rect 87822 558724 87828 558726
rect 87892 558724 87939 558728
rect 87873 558723 87939 558724
rect 100293 558788 100359 558789
rect 100293 558784 100340 558788
rect 100404 558786 100410 558788
rect 100293 558728 100298 558784
rect 100293 558724 100340 558728
rect 100404 558726 100450 558786
rect 100404 558724 100410 558726
rect 101438 558724 101444 558788
rect 101508 558786 101514 558788
rect 102041 558786 102107 558789
rect 106273 558788 106339 558789
rect 106222 558786 106228 558788
rect 101508 558784 102107 558786
rect 101508 558728 102046 558784
rect 102102 558728 102107 558784
rect 101508 558726 102107 558728
rect 106182 558726 106228 558786
rect 106292 558784 106339 558788
rect 106334 558728 106339 558784
rect 101508 558724 101514 558726
rect 100293 558723 100359 558724
rect 102041 558723 102107 558726
rect 106222 558724 106228 558726
rect 106292 558724 106339 558728
rect 106273 558723 106339 558724
rect 108573 558788 108639 558789
rect 108573 558784 108620 558788
rect 108684 558786 108690 558788
rect 195973 558786 196039 558789
rect 196198 558786 196204 558788
rect 108573 558728 108578 558784
rect 108573 558724 108620 558728
rect 108684 558726 108730 558786
rect 195973 558784 196204 558786
rect 195973 558728 195978 558784
rect 196034 558728 196204 558784
rect 195973 558726 196204 558728
rect 108684 558724 108690 558726
rect 108573 558723 108639 558724
rect 195973 558723 196039 558726
rect 196198 558724 196204 558726
rect 196268 558724 196274 558788
rect 201493 558786 201559 558789
rect 201718 558786 201724 558788
rect 201493 558784 201724 558786
rect 201493 558728 201498 558784
rect 201554 558728 201724 558784
rect 201493 558726 201724 558728
rect 201493 558723 201559 558726
rect 201718 558724 201724 558726
rect 201788 558724 201794 558788
rect 202137 558786 202203 558789
rect 204897 558788 204963 558789
rect 202454 558786 202460 558788
rect 202137 558784 202460 558786
rect 202137 558728 202142 558784
rect 202198 558728 202460 558784
rect 202137 558726 202460 558728
rect 202137 558723 202203 558726
rect 202454 558724 202460 558726
rect 202524 558724 202530 558788
rect 204846 558786 204852 558788
rect 204806 558726 204852 558786
rect 204916 558784 204963 558788
rect 204958 558728 204963 558784
rect 204846 558724 204852 558726
rect 204916 558724 204963 558728
rect 204897 558723 204963 558724
rect 215293 558788 215359 558789
rect 215293 558784 215340 558788
rect 215404 558786 215410 558788
rect 215293 558728 215298 558784
rect 215293 558724 215340 558728
rect 215404 558726 215450 558786
rect 215404 558724 215410 558726
rect 216622 558724 216628 558788
rect 216692 558786 216698 558788
rect 216765 558786 216831 558789
rect 216692 558784 216831 558786
rect 216692 558728 216770 558784
rect 216826 558728 216831 558784
rect 216692 558726 216831 558728
rect 216692 558724 216698 558726
rect 215293 558723 215359 558724
rect 216765 558723 216831 558726
rect 217358 558724 217364 558788
rect 217428 558786 217434 558788
rect 217961 558786 218027 558789
rect 217428 558784 218027 558786
rect 217428 558728 217966 558784
rect 218022 558728 218027 558784
rect 217428 558726 218027 558728
rect 217428 558724 217434 558726
rect 217961 558723 218027 558726
rect 223573 558788 223639 558789
rect 223573 558784 223620 558788
rect 223684 558786 223690 558788
rect 224401 558786 224467 558789
rect 224534 558786 224540 558788
rect 223573 558728 223578 558784
rect 223573 558724 223620 558728
rect 223684 558726 223730 558786
rect 224401 558784 224540 558786
rect 224401 558728 224406 558784
rect 224462 558728 224540 558784
rect 224401 558726 224540 558728
rect 223684 558724 223690 558726
rect 223573 558723 223639 558724
rect 224401 558723 224467 558726
rect 224534 558724 224540 558726
rect 224604 558724 224610 558788
rect 225638 558724 225644 558788
rect 225708 558786 225714 558788
rect 226149 558786 226215 558789
rect 225708 558784 226215 558786
rect 225708 558728 226154 558784
rect 226210 558728 226215 558784
rect 225708 558726 226215 558728
rect 225708 558724 225714 558726
rect 226149 558723 226215 558726
rect 227713 558786 227779 558789
rect 227846 558786 227852 558788
rect 227713 558784 227852 558786
rect 227713 558728 227718 558784
rect 227774 558728 227852 558784
rect 227713 558726 227852 558728
rect 227713 558723 227779 558726
rect 227846 558724 227852 558726
rect 227916 558724 227922 558788
rect 232630 558724 232636 558788
rect 232700 558786 232706 558788
rect 233049 558786 233115 558789
rect 232700 558784 233115 558786
rect 232700 558728 233054 558784
rect 233110 558728 233115 558784
rect 232700 558726 233115 558728
rect 232700 558724 232706 558726
rect 233049 558723 233115 558726
rect 233233 558786 233299 558789
rect 233550 558786 233556 558788
rect 233233 558784 233556 558786
rect 233233 558728 233238 558784
rect 233294 558728 233556 558784
rect 233233 558726 233556 558728
rect 233233 558723 233299 558726
rect 233550 558724 233556 558726
rect 233620 558724 233626 558788
rect 235993 558786 236059 558789
rect 236126 558786 236132 558788
rect 235993 558784 236132 558786
rect 235993 558728 235998 558784
rect 236054 558728 236132 558784
rect 235993 558726 236132 558728
rect 235993 558723 236059 558726
rect 236126 558724 236132 558726
rect 236196 558724 236202 558788
rect 322289 558786 322355 558789
rect 322422 558786 322428 558788
rect 322289 558784 322428 558786
rect 322289 558728 322294 558784
rect 322350 558728 322428 558784
rect 322289 558726 322428 558728
rect 322289 558723 322355 558726
rect 322422 558724 322428 558726
rect 322492 558724 322498 558788
rect 327022 558724 327028 558788
rect 327092 558786 327098 558788
rect 327717 558786 327783 558789
rect 327092 558784 327783 558786
rect 327092 558728 327722 558784
rect 327778 558728 327783 558784
rect 327092 558726 327783 558728
rect 327092 558724 327098 558726
rect 327717 558723 327783 558726
rect 328494 558724 328500 558788
rect 328564 558786 328570 558788
rect 329097 558786 329163 558789
rect 328564 558784 329163 558786
rect 328564 558728 329102 558784
rect 329158 558728 329163 558784
rect 328564 558726 329163 558728
rect 328564 558724 328570 558726
rect 329097 558723 329163 558726
rect 332685 558788 332751 558789
rect 334065 558788 334131 558789
rect 332685 558784 332732 558788
rect 332796 558786 332802 558788
rect 334014 558786 334020 558788
rect 332685 558728 332690 558784
rect 332685 558724 332732 558728
rect 332796 558726 332842 558786
rect 333974 558726 334020 558786
rect 334084 558784 334131 558788
rect 334126 558728 334131 558784
rect 332796 558724 332802 558726
rect 334014 558724 334020 558726
rect 334084 558724 334131 558728
rect 332685 558723 332751 558724
rect 334065 558723 334131 558724
rect 335445 558788 335511 558789
rect 336641 558788 336707 558789
rect 335445 558784 335492 558788
rect 335556 558786 335562 558788
rect 336590 558786 336596 558788
rect 335445 558728 335450 558784
rect 335445 558724 335492 558728
rect 335556 558726 335602 558786
rect 336550 558726 336596 558786
rect 336660 558784 336707 558788
rect 336702 558728 336707 558784
rect 335556 558724 335562 558726
rect 336590 558724 336596 558726
rect 336660 558724 336707 558728
rect 335445 558723 335511 558724
rect 336641 558723 336707 558724
rect 338941 558788 339007 558789
rect 339861 558788 339927 558789
rect 340965 558788 341031 558789
rect 342529 558788 342595 558789
rect 338941 558784 338988 558788
rect 339052 558786 339058 558788
rect 338941 558728 338946 558784
rect 338941 558724 338988 558728
rect 339052 558726 339098 558786
rect 339861 558784 339908 558788
rect 339972 558786 339978 558788
rect 339861 558728 339866 558784
rect 339052 558724 339058 558726
rect 339861 558724 339908 558728
rect 339972 558726 340018 558786
rect 340965 558784 341012 558788
rect 341076 558786 341082 558788
rect 342478 558786 342484 558788
rect 340965 558728 340970 558784
rect 339972 558724 339978 558726
rect 340965 558724 341012 558728
rect 341076 558726 341122 558786
rect 342438 558726 342484 558786
rect 342548 558784 342595 558788
rect 342590 558728 342595 558784
rect 341076 558724 341082 558726
rect 342478 558724 342484 558726
rect 342548 558724 342595 558728
rect 343582 558724 343588 558788
rect 343652 558786 343658 558788
rect 343725 558786 343791 558789
rect 343652 558784 343791 558786
rect 343652 558728 343730 558784
rect 343786 558728 343791 558784
rect 343652 558726 343791 558728
rect 343652 558724 343658 558726
rect 338941 558723 339007 558724
rect 339861 558723 339927 558724
rect 340965 558723 341031 558724
rect 342529 558723 342595 558724
rect 343725 558723 343791 558726
rect 345974 558724 345980 558788
rect 346044 558786 346050 558788
rect 346301 558786 346367 558789
rect 346945 558788 347011 558789
rect 346894 558786 346900 558788
rect 346044 558784 346367 558786
rect 346044 558728 346306 558784
rect 346362 558728 346367 558784
rect 346044 558726 346367 558728
rect 346854 558726 346900 558786
rect 346964 558784 347011 558788
rect 347006 558728 347011 558784
rect 346044 558724 346050 558726
rect 346301 558723 346367 558726
rect 346894 558724 346900 558726
rect 346964 558724 347011 558728
rect 348182 558724 348188 558788
rect 348252 558786 348258 558788
rect 348325 558786 348391 558789
rect 349521 558788 349587 558789
rect 349470 558786 349476 558788
rect 348252 558784 348391 558786
rect 348252 558728 348330 558784
rect 348386 558728 348391 558784
rect 348252 558726 348391 558728
rect 349430 558726 349476 558786
rect 349540 558784 349587 558788
rect 349582 558728 349587 558784
rect 348252 558724 348258 558726
rect 346945 558723 347011 558724
rect 348325 558723 348391 558726
rect 349470 558724 349476 558726
rect 349540 558724 349587 558728
rect 349521 558723 349587 558724
rect 353293 558786 353359 558789
rect 353518 558786 353524 558788
rect 353293 558784 353524 558786
rect 353293 558728 353298 558784
rect 353354 558728 353524 558784
rect 353293 558726 353524 558728
rect 353293 558723 353359 558726
rect 353518 558724 353524 558726
rect 353588 558724 353594 558788
rect 357433 558786 357499 558789
rect 357566 558786 357572 558788
rect 357433 558784 357572 558786
rect 357433 558728 357438 558784
rect 357494 558728 357572 558784
rect 357433 558726 357572 558728
rect 357433 558723 357499 558726
rect 357566 558724 357572 558726
rect 357636 558724 357642 558788
rect 452694 558724 452700 558788
rect 452764 558786 452770 558788
rect 453297 558786 453363 558789
rect 452764 558784 453363 558786
rect 452764 558728 453302 558784
rect 453358 558728 453363 558784
rect 452764 558726 453363 558728
rect 452764 558724 452770 558726
rect 453297 558723 453363 558726
rect 459502 558724 459508 558788
rect 459572 558786 459578 558788
rect 460197 558786 460263 558789
rect 460657 558786 460723 558789
rect 459572 558784 460723 558786
rect 459572 558728 460202 558784
rect 460258 558728 460662 558784
rect 460718 558728 460723 558784
rect 459572 558726 460723 558728
rect 459572 558724 459578 558726
rect 460197 558723 460263 558726
rect 460657 558723 460723 558726
rect 461025 558786 461091 558789
rect 462957 558788 463023 558789
rect 464337 558788 464403 558789
rect 462078 558786 462084 558788
rect 461025 558784 462084 558786
rect 461025 558728 461030 558784
rect 461086 558728 462084 558784
rect 461025 558726 462084 558728
rect 461025 558723 461091 558726
rect 462078 558724 462084 558726
rect 462148 558724 462154 558788
rect 462957 558784 463004 558788
rect 463068 558786 463074 558788
rect 464286 558786 464292 558788
rect 462957 558728 462962 558784
rect 462957 558724 463004 558728
rect 463068 558726 463114 558786
rect 464246 558726 464292 558786
rect 464356 558784 464403 558788
rect 464398 558728 464403 558784
rect 463068 558724 463074 558726
rect 464286 558724 464292 558726
rect 464356 558724 464403 558728
rect 462957 558723 463023 558724
rect 464337 558723 464403 558724
rect 465165 558788 465231 558789
rect 465165 558784 465212 558788
rect 465276 558786 465282 558788
rect 467925 558786 467991 558789
rect 470041 558788 470107 558789
rect 469070 558786 469076 558788
rect 465165 558728 465170 558784
rect 465165 558724 465212 558728
rect 465276 558726 465322 558786
rect 467925 558784 469076 558786
rect 467925 558728 467930 558784
rect 467986 558728 469076 558784
rect 467925 558726 469076 558728
rect 465276 558724 465282 558726
rect 465165 558723 465231 558724
rect 467925 558723 467991 558726
rect 469070 558724 469076 558726
rect 469140 558724 469146 558788
rect 469990 558786 469996 558788
rect 469950 558726 469996 558786
rect 470060 558784 470107 558788
rect 470102 558728 470107 558784
rect 469990 558724 469996 558726
rect 470060 558724 470107 558728
rect 470041 558723 470107 558724
rect 471237 558788 471303 558789
rect 472249 558788 472315 558789
rect 473537 558788 473603 558789
rect 474825 558788 474891 558789
rect 475561 558788 475627 558789
rect 471237 558784 471284 558788
rect 471348 558786 471354 558788
rect 472198 558786 472204 558788
rect 471237 558728 471242 558784
rect 471237 558724 471284 558728
rect 471348 558726 471394 558786
rect 472158 558726 472204 558786
rect 472268 558784 472315 558788
rect 473486 558786 473492 558788
rect 472310 558728 472315 558784
rect 471348 558724 471354 558726
rect 472198 558724 472204 558726
rect 472268 558724 472315 558728
rect 473446 558726 473492 558786
rect 473556 558784 473603 558788
rect 474774 558786 474780 558788
rect 473598 558728 473603 558784
rect 473486 558724 473492 558726
rect 473556 558724 473603 558728
rect 474734 558726 474780 558786
rect 474844 558784 474891 558788
rect 474886 558728 474891 558784
rect 474774 558724 474780 558726
rect 474844 558724 474891 558728
rect 475510 558724 475516 558788
rect 475580 558786 475627 558788
rect 480437 558788 480503 558789
rect 480437 558786 480484 558788
rect 475580 558784 475672 558786
rect 475622 558728 475672 558784
rect 475580 558726 475672 558728
rect 480392 558784 480484 558786
rect 480392 558728 480442 558784
rect 480392 558726 480484 558728
rect 475580 558724 475627 558726
rect 471237 558723 471303 558724
rect 472249 558723 472315 558724
rect 473537 558723 473603 558724
rect 474825 558723 474891 558724
rect 475561 558723 475627 558724
rect 480437 558724 480484 558726
rect 480548 558724 480554 558788
rect 484393 558786 484459 558789
rect 484710 558786 484716 558788
rect 484393 558784 484716 558786
rect 484393 558728 484398 558784
rect 484454 558728 484716 558784
rect 484393 558726 484716 558728
rect 480437 558723 480503 558724
rect 484393 558723 484459 558726
rect 484710 558724 484716 558726
rect 484780 558724 484786 558788
rect 101857 558652 101923 558653
rect 101806 558650 101812 558652
rect 101766 558590 101812 558650
rect 101876 558648 101923 558652
rect 101918 558592 101923 558648
rect 101806 558588 101812 558590
rect 101876 558588 101923 558592
rect 101857 558587 101923 558588
rect 197353 558650 197419 558653
rect 197486 558650 197492 558652
rect 197353 558648 197492 558650
rect 197353 558592 197358 558648
rect 197414 558592 197492 558648
rect 197353 558590 197492 558592
rect 197353 558587 197419 558590
rect 197486 558588 197492 558590
rect 197556 558588 197562 558652
rect 203517 558650 203583 558653
rect 203742 558650 203748 558652
rect 203517 558648 203748 558650
rect 203517 558592 203522 558648
rect 203578 558592 203748 558648
rect 203517 558590 203748 558592
rect 203517 558587 203583 558590
rect 203742 558588 203748 558590
rect 203812 558588 203818 558652
rect 209037 558650 209103 558653
rect 209630 558650 209636 558652
rect 209037 558648 209636 558650
rect 209037 558592 209042 558648
rect 209098 558592 209636 558648
rect 209037 558590 209636 558592
rect 209037 558587 209103 558590
rect 209630 558588 209636 558590
rect 209700 558588 209706 558652
rect 230473 558650 230539 558653
rect 231853 558652 231919 558653
rect 234613 558652 234679 558653
rect 230606 558650 230612 558652
rect 230473 558648 230612 558650
rect 230473 558592 230478 558648
rect 230534 558592 230612 558648
rect 230473 558590 230612 558592
rect 230473 558587 230539 558590
rect 230606 558588 230612 558590
rect 230676 558588 230682 558652
rect 231853 558650 231900 558652
rect 231808 558648 231900 558650
rect 231808 558592 231858 558648
rect 231808 558590 231900 558592
rect 231853 558588 231900 558590
rect 231964 558588 231970 558652
rect 234613 558650 234660 558652
rect 234568 558648 234660 558650
rect 234568 558592 234618 558648
rect 234568 558590 234660 558592
rect 234613 558588 234660 558590
rect 234724 558588 234730 558652
rect 323526 558588 323532 558652
rect 323596 558650 323602 558652
rect 323669 558650 323735 558653
rect 323596 558648 323735 558650
rect 323596 558592 323674 558648
rect 323730 558592 323735 558648
rect 323596 558590 323735 558592
rect 323596 558588 323602 558590
rect 231853 558587 231919 558588
rect 234613 558587 234679 558588
rect 323669 558587 323735 558590
rect 324814 558588 324820 558652
rect 324884 558650 324890 558652
rect 324957 558650 325023 558653
rect 324884 558648 325023 558650
rect 324884 558592 324962 558648
rect 325018 558592 325023 558648
rect 324884 558590 325023 558592
rect 324884 558588 324890 558590
rect 324957 558587 325023 558590
rect 326102 558588 326108 558652
rect 326172 558650 326178 558652
rect 326337 558650 326403 558653
rect 326172 558648 326403 558650
rect 326172 558592 326342 558648
rect 326398 558592 326403 558648
rect 326172 558590 326403 558592
rect 326172 558588 326178 558590
rect 326337 558587 326403 558590
rect 329281 558650 329347 558653
rect 330477 558652 330543 558653
rect 356053 558652 356119 558653
rect 456057 558652 456123 558653
rect 329598 558650 329604 558652
rect 329281 558648 329604 558650
rect 329281 558592 329286 558648
rect 329342 558592 329604 558648
rect 329281 558590 329604 558592
rect 329281 558587 329347 558590
rect 329598 558588 329604 558590
rect 329668 558588 329674 558652
rect 330477 558648 330524 558652
rect 330588 558650 330594 558652
rect 356053 558650 356100 558652
rect 330477 558592 330482 558648
rect 330477 558588 330524 558592
rect 330588 558590 330634 558650
rect 356008 558648 356100 558650
rect 356008 558592 356058 558648
rect 356008 558590 356100 558592
rect 330588 558588 330594 558590
rect 356053 558588 356100 558590
rect 356164 558588 356170 558652
rect 456006 558650 456012 558652
rect 455966 558590 456012 558650
rect 456076 558648 456123 558652
rect 456118 558592 456123 558648
rect 456006 558588 456012 558590
rect 456076 558588 456123 558592
rect 457294 558588 457300 558652
rect 457364 558650 457370 558652
rect 457437 558650 457503 558653
rect 460841 558652 460907 558653
rect 466545 558652 466611 558653
rect 460790 558650 460796 558652
rect 457364 558648 457503 558650
rect 457364 558592 457442 558648
rect 457498 558592 457503 558648
rect 457364 558590 457503 558592
rect 460750 558590 460796 558650
rect 460860 558648 460907 558652
rect 466494 558650 466500 558652
rect 460902 558592 460907 558648
rect 457364 558588 457370 558590
rect 330477 558587 330543 558588
rect 356053 558587 356119 558588
rect 456057 558587 456123 558588
rect 457437 558587 457503 558590
rect 460790 558588 460796 558590
rect 460860 558588 460907 558592
rect 466454 558590 466500 558650
rect 466564 558648 466611 558652
rect 466606 558592 466611 558648
rect 466494 558588 466500 558590
rect 466564 558588 466611 558592
rect 467782 558588 467788 558652
rect 467852 558650 467858 558652
rect 468017 558650 468083 558653
rect 483013 558652 483079 558653
rect 488533 558652 488599 558653
rect 483013 558650 483060 558652
rect 467852 558648 468083 558650
rect 467852 558592 468022 558648
rect 468078 558592 468083 558648
rect 467852 558590 468083 558592
rect 482968 558648 483060 558650
rect 482968 558592 483018 558648
rect 482968 558590 483060 558592
rect 467852 558588 467858 558590
rect 460841 558587 460907 558588
rect 466545 558587 466611 558588
rect 468017 558587 468083 558590
rect 483013 558588 483060 558590
rect 483124 558588 483130 558652
rect 488533 558650 488580 558652
rect 488488 558648 488580 558650
rect 488488 558592 488538 558648
rect 488488 558590 488580 558592
rect 488533 558588 488580 558590
rect 488644 558588 488650 558652
rect 483013 558587 483079 558588
rect 488533 558587 488599 558588
rect 198733 558516 198799 558517
rect 200205 558516 200271 558517
rect 237373 558516 237439 558517
rect 238753 558516 238819 558517
rect 198733 558514 198780 558516
rect 198688 558512 198780 558514
rect 198688 558456 198738 558512
rect 198688 558454 198780 558456
rect 198733 558452 198780 558454
rect 198844 558452 198850 558516
rect 200205 558514 200252 558516
rect 200160 558512 200252 558514
rect 200160 558456 200210 558512
rect 200160 558454 200252 558456
rect 200205 558452 200252 558454
rect 200316 558452 200322 558516
rect 237373 558514 237420 558516
rect 237328 558512 237420 558514
rect 237328 558456 237378 558512
rect 237328 558454 237420 558456
rect 237373 558452 237420 558454
rect 237484 558452 237490 558516
rect 238702 558452 238708 558516
rect 238772 558514 238819 558516
rect 317413 558516 317479 558517
rect 317413 558514 317460 558516
rect 238772 558512 238864 558514
rect 238814 558456 238864 558512
rect 238772 558454 238864 558456
rect 317368 558512 317460 558514
rect 317368 558456 317418 558512
rect 317368 558454 317460 558456
rect 238772 558452 238819 558454
rect 198733 558451 198799 558452
rect 200205 558451 200271 558452
rect 237373 558451 237439 558452
rect 238753 558451 238819 558452
rect 317413 558452 317460 558454
rect 317524 558452 317530 558516
rect 336825 558514 336891 558517
rect 350533 558516 350599 558517
rect 337878 558514 337884 558516
rect 336825 558512 337884 558514
rect 336825 558456 336830 558512
rect 336886 558456 337884 558512
rect 336825 558454 337884 558456
rect 317413 558451 317479 558452
rect 336825 558451 336891 558454
rect 337878 558452 337884 558454
rect 337948 558452 337954 558516
rect 350533 558512 350580 558516
rect 350644 558514 350650 558516
rect 455413 558514 455479 558517
rect 481633 558516 481699 558517
rect 456558 558514 456564 558516
rect 350533 558456 350538 558512
rect 350533 558452 350580 558456
rect 350644 558454 350690 558514
rect 455413 558512 456564 558514
rect 455413 558456 455418 558512
rect 455474 558456 456564 558512
rect 455413 558454 456564 558456
rect 350644 558452 350650 558454
rect 350533 558451 350599 558452
rect 455413 558451 455479 558454
rect 456558 558452 456564 558454
rect 456628 558452 456634 558516
rect 481582 558452 481588 558516
rect 481652 558514 481699 558516
rect 487153 558514 487219 558517
rect 487286 558514 487292 558516
rect 481652 558512 481744 558514
rect 481694 558456 481744 558512
rect 481652 558454 481744 558456
rect 487153 558512 487292 558514
rect 487153 558456 487158 558512
rect 487214 558456 487292 558512
rect 487153 558454 487292 558456
rect 481652 558452 481699 558454
rect 481633 558451 481699 558452
rect 487153 558451 487219 558454
rect 487286 558452 487292 558454
rect 487356 558452 487362 558516
rect 77293 558378 77359 558381
rect 77702 558378 77708 558380
rect 77293 558376 77708 558378
rect 77293 558320 77298 558376
rect 77354 558320 77708 558376
rect 77293 558318 77708 558320
rect 77293 558315 77359 558318
rect 77702 558316 77708 558318
rect 77772 558316 77778 558380
rect 82813 558378 82879 558381
rect 329833 558380 329899 558381
rect 83406 558378 83412 558380
rect 82813 558376 83412 558378
rect 82813 558320 82818 558376
rect 82874 558320 83412 558376
rect 82813 558318 83412 558320
rect 82813 558315 82879 558318
rect 83406 558316 83412 558318
rect 83476 558316 83482 558380
rect 329782 558316 329788 558380
rect 329852 558378 329899 558380
rect 354673 558378 354739 558381
rect 354806 558378 354812 558380
rect 329852 558376 329944 558378
rect 329894 558320 329944 558376
rect 329852 558318 329944 558320
rect 354673 558376 354812 558378
rect 354673 558320 354678 558376
rect 354734 558320 354812 558376
rect 354673 558318 354812 558320
rect 329852 558316 329899 558318
rect 329833 558315 329899 558316
rect 354673 558315 354739 558318
rect 354806 558316 354812 558318
rect 354876 558316 354882 558380
rect 454033 558378 454099 558381
rect 455270 558378 455276 558380
rect 454033 558376 455276 558378
rect 454033 558320 454038 558376
rect 454094 558320 455276 558376
rect 454033 558318 455276 558320
rect 454033 558315 454099 558318
rect 455270 558316 455276 558318
rect 455340 558316 455346 558380
rect 456793 558378 456859 558381
rect 457478 558378 457484 558380
rect 456793 558376 457484 558378
rect 456793 558320 456798 558376
rect 456854 558320 457484 558376
rect 456793 558318 457484 558320
rect 456793 558315 456859 558318
rect 457478 558316 457484 558318
rect 457548 558316 457554 558380
rect 458173 558378 458239 558381
rect 458766 558378 458772 558380
rect 458173 558376 458772 558378
rect 458173 558320 458178 558376
rect 458234 558320 458772 558376
rect 458173 558318 458772 558320
rect 458173 558315 458239 558318
rect 458766 558316 458772 558318
rect 458836 558316 458842 558380
rect 488533 558378 488599 558381
rect 489126 558378 489132 558380
rect 488533 558376 489132 558378
rect 488533 558320 488538 558376
rect 488594 558320 489132 558376
rect 488533 558318 489132 558320
rect 488533 558315 488599 558318
rect 489126 558316 489132 558318
rect 489196 558316 489202 558380
rect 73153 558242 73219 558245
rect 74206 558242 74212 558244
rect 73153 558240 74212 558242
rect 73153 558184 73158 558240
rect 73214 558184 74212 558240
rect 73153 558182 74212 558184
rect 73153 558179 73219 558182
rect 74206 558180 74212 558182
rect 74276 558180 74282 558244
rect 328453 558242 328519 558245
rect 328862 558242 328868 558244
rect 328453 558240 328868 558242
rect 328453 558184 328458 558240
rect 328514 558184 328868 558240
rect 328453 558182 328868 558184
rect 328453 558179 328519 558182
rect 328862 558180 328868 558182
rect 328932 558180 328938 558244
rect 331213 558242 331279 558245
rect 332358 558242 332364 558244
rect 331213 558240 332364 558242
rect 331213 558184 331218 558240
rect 331274 558184 332364 558240
rect 331213 558182 332364 558184
rect 331213 558179 331279 558182
rect 332358 558180 332364 558182
rect 332428 558180 332434 558244
rect 452653 558242 452719 558245
rect 453798 558242 453804 558244
rect 452653 558240 453804 558242
rect 452653 558184 452658 558240
rect 452714 558184 453804 558240
rect 452653 558182 453804 558184
rect 452653 558179 452719 558182
rect 453798 558180 453804 558182
rect 453868 558180 453874 558244
rect 459553 558242 459619 558245
rect 459870 558242 459876 558244
rect 459553 558240 459876 558242
rect 459553 558184 459558 558240
rect 459614 558184 459876 558240
rect 459553 558182 459876 558184
rect 459553 558179 459619 558182
rect 459870 558180 459876 558182
rect 459940 558180 459946 558244
rect 483013 558242 483079 558245
rect 484158 558242 484164 558244
rect 483013 558240 484164 558242
rect 483013 558184 483018 558240
rect 483074 558184 484164 558240
rect 483013 558182 484164 558184
rect 483013 558179 483079 558182
rect 484158 558180 484164 558182
rect 484228 558180 484234 558244
rect 485773 558242 485839 558245
rect 486918 558242 486924 558244
rect 485773 558240 486924 558242
rect 485773 558184 485778 558240
rect 485834 558184 486924 558240
rect 485773 558182 486924 558184
rect 485773 558179 485839 558182
rect 486918 558180 486924 558182
rect 486988 558180 486994 558244
rect 487153 558242 487219 558245
rect 487838 558242 487844 558244
rect 487153 558240 487844 558242
rect 487153 558184 487158 558240
rect 487214 558184 487844 558240
rect 487153 558182 487844 558184
rect 487153 558179 487219 558182
rect 487838 558180 487844 558182
rect 487908 558180 487914 558244
rect 68502 558044 68508 558108
rect 68572 558106 68578 558108
rect 68921 558106 68987 558109
rect 68572 558104 68987 558106
rect 68572 558048 68926 558104
rect 68982 558048 68987 558104
rect 68572 558046 68987 558048
rect 68572 558044 68578 558046
rect 68921 558043 68987 558046
rect 206134 558044 206140 558108
rect 206204 558106 206210 558108
rect 206277 558106 206343 558109
rect 206204 558104 206343 558106
rect 206204 558048 206282 558104
rect 206338 558048 206343 558104
rect 206204 558046 206343 558048
rect 206204 558044 206210 558046
rect 206277 558043 206343 558046
rect 238334 558044 238340 558108
rect 238404 558106 238410 558108
rect 238661 558106 238727 558109
rect 238404 558104 238727 558106
rect 238404 558048 238666 558104
rect 238722 558048 238727 558104
rect 238404 558046 238727 558048
rect 238404 558044 238410 558046
rect 238661 558043 238727 558046
rect 476113 558106 476179 558109
rect 477350 558106 477356 558108
rect 476113 558104 477356 558106
rect 476113 558048 476118 558104
rect 476174 558048 477356 558104
rect 476113 558046 477356 558048
rect 476113 558043 476179 558046
rect 477350 558044 477356 558046
rect 477420 558044 477426 558108
rect 477493 558106 477559 558109
rect 478454 558106 478460 558108
rect 477493 558104 478460 558106
rect 477493 558048 477498 558104
rect 477554 558048 478460 558104
rect 477493 558046 478460 558048
rect 477493 558043 477559 558046
rect 478454 558044 478460 558046
rect 478524 558044 478530 558108
rect 78673 557972 78739 557973
rect 78622 557908 78628 557972
rect 78692 557970 78739 557972
rect 322933 557970 322999 557973
rect 324078 557970 324084 557972
rect 78692 557968 78784 557970
rect 78734 557912 78784 557968
rect 78692 557910 78784 557912
rect 322933 557968 324084 557970
rect 322933 557912 322938 557968
rect 322994 557912 324084 557968
rect 322933 557910 324084 557912
rect 78692 557908 78739 557910
rect 78673 557907 78739 557908
rect 322933 557907 322999 557910
rect 324078 557908 324084 557910
rect 324148 557908 324154 557972
rect 478873 557970 478939 557973
rect 479742 557970 479748 557972
rect 478873 557968 479748 557970
rect 478873 557912 478878 557968
rect 478934 557912 479748 557968
rect 478873 557910 479748 557912
rect 478873 557907 478939 557910
rect 479742 557908 479748 557910
rect 479812 557908 479818 557972
rect 74533 557834 74599 557837
rect 75126 557834 75132 557836
rect 74533 557832 75132 557834
rect 74533 557776 74538 557832
rect 74594 557776 75132 557832
rect 74533 557774 75132 557776
rect 74533 557771 74599 557774
rect 75126 557772 75132 557774
rect 75196 557772 75202 557836
rect 75913 557834 75979 557837
rect 320173 557836 320239 557837
rect 76414 557834 76420 557836
rect 75913 557832 76420 557834
rect 75913 557776 75918 557832
rect 75974 557776 76420 557832
rect 75913 557774 76420 557776
rect 75913 557771 75979 557774
rect 76414 557772 76420 557774
rect 76484 557772 76490 557836
rect 320173 557834 320220 557836
rect 320128 557832 320220 557834
rect 320128 557776 320178 557832
rect 320128 557774 320220 557776
rect 320173 557772 320220 557774
rect 320284 557772 320290 557836
rect 481633 557834 481699 557837
rect 482134 557834 482140 557836
rect 481633 557832 482140 557834
rect 481633 557776 481638 557832
rect 481694 557776 482140 557832
rect 481633 557774 482140 557776
rect 320173 557771 320239 557772
rect 481633 557771 481699 557774
rect 482134 557772 482140 557774
rect 482204 557772 482210 557836
rect 71773 557698 71839 557701
rect 72918 557698 72924 557700
rect 71773 557696 72924 557698
rect 71773 557640 71778 557696
rect 71834 557640 72924 557696
rect 71773 557638 72924 557640
rect 71773 557635 71839 557638
rect 72918 557636 72924 557638
rect 72988 557636 72994 557700
rect 78673 557698 78739 557701
rect 79910 557698 79916 557700
rect 78673 557696 79916 557698
rect 78673 557640 78678 557696
rect 78734 557640 79916 557696
rect 78673 557638 79916 557640
rect 78673 557635 78739 557638
rect 79910 557636 79916 557638
rect 79980 557636 79986 557700
rect 93158 557636 93164 557700
rect 93228 557698 93234 557700
rect 93669 557698 93735 557701
rect 93228 557696 93735 557698
rect 93228 557640 93674 557696
rect 93730 557640 93735 557696
rect 93228 557638 93735 557640
rect 93228 557636 93234 557638
rect 93669 557635 93735 557638
rect 207054 557636 207060 557700
rect 207124 557698 207130 557700
rect 207657 557698 207723 557701
rect 207124 557696 207723 557698
rect 207124 557640 207662 557696
rect 207718 557640 207723 557696
rect 207124 557638 207723 557640
rect 207124 557636 207130 557638
rect 207657 557635 207723 557638
rect 208342 557636 208348 557700
rect 208412 557698 208418 557700
rect 209221 557698 209287 557701
rect 208412 557696 209287 557698
rect 208412 557640 209226 557696
rect 209282 557640 209287 557696
rect 208412 557638 209287 557640
rect 208412 557636 208418 557638
rect 209221 557635 209287 557638
rect 210366 557636 210372 557700
rect 210436 557698 210442 557700
rect 210969 557698 211035 557701
rect 210436 557696 211035 557698
rect 210436 557640 210974 557696
rect 211030 557640 211035 557696
rect 210436 557638 211035 557640
rect 210436 557636 210442 557638
rect 210969 557635 211035 557638
rect 343725 557698 343791 557701
rect 344870 557698 344876 557700
rect 343725 557696 344876 557698
rect 343725 557640 343730 557696
rect 343786 557640 344876 557696
rect 343725 557638 344876 557640
rect 343725 557635 343791 557638
rect 344870 557636 344876 557638
rect 344940 557636 344946 557700
rect 352005 557698 352071 557701
rect 451365 557700 451431 557701
rect 353150 557698 353156 557700
rect 352005 557696 353156 557698
rect 352005 557640 352010 557696
rect 352066 557640 353156 557696
rect 352005 557638 353156 557640
rect 352005 557635 352071 557638
rect 353150 557636 353156 557638
rect 353220 557636 353226 557700
rect 451365 557698 451412 557700
rect 451320 557696 451412 557698
rect 451320 557640 451370 557696
rect 451320 557638 451412 557640
rect 451365 557636 451412 557638
rect 451476 557636 451482 557700
rect 474641 557698 474707 557701
rect 475510 557698 475516 557700
rect 474641 557696 475516 557698
rect 474641 557640 474646 557696
rect 474702 557640 475516 557696
rect 474641 557638 475516 557640
rect 451365 557635 451431 557636
rect 474641 557635 474707 557638
rect 475510 557636 475516 557638
rect 475580 557636 475586 557700
rect 483013 557698 483079 557701
rect 483606 557698 483612 557700
rect 483013 557696 483612 557698
rect 483013 557640 483018 557696
rect 483074 557640 483612 557696
rect 483013 557638 483612 557640
rect 483013 557635 483079 557638
rect 483606 557636 483612 557638
rect 483676 557636 483682 557700
rect 71446 557500 71452 557564
rect 71516 557562 71522 557564
rect 71589 557562 71655 557565
rect 91001 557564 91067 557565
rect 71516 557560 71655 557562
rect 71516 557504 71594 557560
rect 71650 557504 71655 557560
rect 71516 557502 71655 557504
rect 71516 557500 71522 557502
rect 71589 557499 71655 557502
rect 90950 557500 90956 557564
rect 91020 557562 91067 557564
rect 91020 557560 91112 557562
rect 91062 557504 91112 557560
rect 91020 557502 91112 557504
rect 91020 557500 91067 557502
rect 92054 557500 92060 557564
rect 92124 557562 92130 557564
rect 92381 557562 92447 557565
rect 93761 557564 93827 557565
rect 92124 557560 92447 557562
rect 92124 557504 92386 557560
rect 92442 557504 92447 557560
rect 92124 557502 92447 557504
rect 92124 557500 92130 557502
rect 91001 557499 91067 557500
rect 92381 557499 92447 557502
rect 93710 557500 93716 557564
rect 93780 557562 93827 557564
rect 93780 557560 93872 557562
rect 93822 557504 93872 557560
rect 93780 557502 93872 557504
rect 93780 557500 93827 557502
rect 94998 557500 95004 557564
rect 95068 557562 95074 557564
rect 95141 557562 95207 557565
rect 96521 557564 96587 557565
rect 95068 557560 95207 557562
rect 95068 557504 95146 557560
rect 95202 557504 95207 557560
rect 95068 557502 95207 557504
rect 95068 557500 95074 557502
rect 93761 557499 93827 557500
rect 95141 557499 95207 557502
rect 96470 557500 96476 557564
rect 96540 557562 96587 557564
rect 96540 557560 96632 557562
rect 96582 557504 96632 557560
rect 96540 557502 96632 557504
rect 96540 557500 96587 557502
rect 97758 557500 97764 557564
rect 97828 557562 97834 557564
rect 97901 557562 97967 557565
rect 97828 557560 97967 557562
rect 97828 557504 97906 557560
rect 97962 557504 97967 557560
rect 97828 557502 97967 557504
rect 97828 557500 97834 557502
rect 96521 557499 96587 557500
rect 97901 557499 97967 557502
rect 99046 557500 99052 557564
rect 99116 557562 99122 557564
rect 99281 557562 99347 557565
rect 206921 557564 206987 557565
rect 99116 557560 99347 557562
rect 99116 557504 99286 557560
rect 99342 557504 99347 557560
rect 99116 557502 99347 557504
rect 99116 557500 99122 557502
rect 99281 557499 99347 557502
rect 206870 557500 206876 557564
rect 206940 557562 206987 557564
rect 206940 557560 207032 557562
rect 206982 557504 207032 557560
rect 206940 557502 207032 557504
rect 206940 557500 206987 557502
rect 207974 557500 207980 557564
rect 208044 557562 208050 557564
rect 208301 557562 208367 557565
rect 208044 557560 208367 557562
rect 208044 557504 208306 557560
rect 208362 557504 208367 557560
rect 208044 557502 208367 557504
rect 208044 557500 208050 557502
rect 206921 557499 206987 557500
rect 208301 557499 208367 557502
rect 209262 557500 209268 557564
rect 209332 557562 209338 557564
rect 209681 557562 209747 557565
rect 212441 557564 212507 557565
rect 209332 557560 209747 557562
rect 209332 557504 209686 557560
rect 209742 557504 209747 557560
rect 209332 557502 209747 557504
rect 209332 557500 209338 557502
rect 209681 557499 209747 557502
rect 212390 557500 212396 557564
rect 212460 557562 212507 557564
rect 212460 557560 212552 557562
rect 212502 557504 212552 557560
rect 212460 557502 212552 557504
rect 212460 557500 212507 557502
rect 213494 557500 213500 557564
rect 213564 557562 213570 557564
rect 213821 557562 213887 557565
rect 213564 557560 213887 557562
rect 213564 557504 213826 557560
rect 213882 557504 213887 557560
rect 213564 557502 213887 557504
rect 213564 557500 213570 557502
rect 212441 557499 212507 557500
rect 213821 557499 213887 557502
rect 214782 557500 214788 557564
rect 214852 557562 214858 557564
rect 215201 557562 215267 557565
rect 214852 557560 215267 557562
rect 214852 557504 215206 557560
rect 215262 557504 215267 557560
rect 214852 557502 215267 557504
rect 214852 557500 214858 557502
rect 215201 557499 215267 557502
rect 350533 557562 350599 557565
rect 350942 557562 350948 557564
rect 350533 557560 350948 557562
rect 350533 557504 350538 557560
rect 350594 557504 350948 557560
rect 350533 557502 350948 557504
rect 350533 557499 350599 557502
rect 350942 557500 350948 557502
rect 351012 557500 351018 557564
rect 353293 557562 353359 557565
rect 354438 557562 354444 557564
rect 353293 557560 354444 557562
rect 353293 557504 353298 557560
rect 353354 557504 354444 557560
rect 353293 557502 354444 557504
rect 353293 557499 353359 557502
rect 354438 557500 354444 557502
rect 354508 557500 354514 557564
rect 354765 557562 354831 557565
rect 355542 557562 355548 557564
rect 354765 557560 355548 557562
rect 354765 557504 354770 557560
rect 354826 557504 355548 557560
rect 354765 557502 355548 557504
rect 354765 557499 354831 557502
rect 355542 557500 355548 557502
rect 355612 557500 355618 557564
rect 356053 557562 356119 557565
rect 356646 557562 356652 557564
rect 356053 557560 356652 557562
rect 356053 557504 356058 557560
rect 356114 557504 356652 557560
rect 356053 557502 356652 557504
rect 356053 557499 356119 557502
rect 356646 557500 356652 557502
rect 356716 557500 356722 557564
rect 357433 557562 357499 557565
rect 357934 557562 357940 557564
rect 357433 557560 357940 557562
rect 357433 557504 357438 557560
rect 357494 557504 357940 557560
rect 357433 557502 357940 557504
rect 357433 557499 357499 557502
rect 357934 557500 357940 557502
rect 358004 557500 358010 557564
rect 579613 557290 579679 557293
rect 583520 557290 584960 557380
rect 579613 557288 584960 557290
rect 579613 557232 579618 557288
rect 579674 557232 584960 557288
rect 579613 557230 584960 557232
rect 579613 557227 579679 557230
rect 583520 557140 584960 557230
rect 352189 555524 352255 555525
rect 352189 555522 352236 555524
rect 352144 555520 352236 555522
rect 352144 555464 352194 555520
rect 352144 555462 352236 555464
rect 352189 555460 352236 555462
rect 352300 555460 352306 555524
rect 358813 555522 358879 555525
rect 359222 555522 359228 555524
rect 358813 555520 359228 555522
rect 358813 555464 358818 555520
rect 358874 555464 359228 555520
rect 358813 555462 359228 555464
rect 352189 555459 352255 555460
rect 358813 555459 358879 555462
rect 359222 555460 359228 555462
rect 359292 555460 359298 555524
rect -960 553074 480 553164
rect 3877 553074 3943 553077
rect -960 553072 3943 553074
rect -960 553016 3882 553072
rect 3938 553016 3943 553072
rect -960 553014 3943 553016
rect -960 552924 480 553014
rect 3877 553011 3943 553014
rect 211245 550626 211311 550629
rect 211429 550626 211495 550629
rect 211245 550624 211495 550626
rect 211245 550568 211250 550624
rect 211306 550568 211434 550624
rect 211490 550568 211495 550624
rect 211245 550566 211495 550568
rect 211245 550563 211311 550566
rect 211429 550563 211495 550566
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 56593 543010 56659 543013
rect 158529 543010 158595 543013
rect 56593 543008 158595 543010
rect 56593 542952 56598 543008
rect 56654 542952 158534 543008
rect 158590 542952 158595 543008
rect 56593 542950 158595 542952
rect 56593 542947 56659 542950
rect 158529 542947 158595 542950
rect 57462 539140 57468 539204
rect 57532 539202 57538 539204
rect 580257 539202 580323 539205
rect 57532 539200 580323 539202
rect 57532 539144 580262 539200
rect 580318 539144 580323 539200
rect 57532 539142 580323 539144
rect 57532 539140 57538 539142
rect 580257 539139 580323 539142
rect 57646 539004 57652 539068
rect 57716 539066 57722 539068
rect 580441 539066 580507 539069
rect 57716 539064 580507 539066
rect 57716 539008 580446 539064
rect 580502 539008 580507 539064
rect 57716 539006 580507 539008
rect 57716 539004 57722 539006
rect 580441 539003 580507 539006
rect 57237 538930 57303 538933
rect 281717 538930 281783 538933
rect 57237 538928 60076 538930
rect 57237 538872 57242 538928
rect 57298 538872 60076 538928
rect 57237 538870 60076 538872
rect 279956 538928 281783 538930
rect 279956 538872 281722 538928
rect 281778 538872 281783 538928
rect 279956 538870 281783 538872
rect 57237 538867 57303 538870
rect 281717 538867 281783 538870
rect -960 538658 480 538748
rect 2957 538658 3023 538661
rect -960 538656 3023 538658
rect -960 538600 2962 538656
rect 3018 538600 3023 538656
rect -960 538598 3023 538600
rect -960 538508 480 538598
rect 2957 538595 3023 538598
rect 57237 536890 57303 536893
rect 57237 536888 60076 536890
rect 57237 536832 57242 536888
rect 57298 536832 60076 536888
rect 57237 536830 60076 536832
rect 57237 536827 57303 536830
rect 282821 536754 282887 536757
rect 279956 536752 282887 536754
rect 279956 536696 282826 536752
rect 282882 536696 282887 536752
rect 279956 536694 282887 536696
rect 282821 536691 282887 536694
rect 57237 534714 57303 534717
rect 57237 534712 60076 534714
rect 57237 534656 57242 534712
rect 57298 534656 60076 534712
rect 57237 534654 60076 534656
rect 57237 534651 57303 534654
rect 282821 534578 282887 534581
rect 279956 534576 282887 534578
rect 279956 534520 282826 534576
rect 282882 534520 282887 534576
rect 279956 534518 282887 534520
rect 282821 534515 282887 534518
rect 579797 533898 579863 533901
rect 583520 533898 584960 533988
rect 579797 533896 584960 533898
rect 579797 533840 579802 533896
rect 579858 533840 584960 533896
rect 579797 533838 584960 533840
rect 579797 533835 579863 533838
rect 583520 533748 584960 533838
rect 57237 532674 57303 532677
rect 57237 532672 60076 532674
rect 57237 532616 57242 532672
rect 57298 532616 60076 532672
rect 57237 532614 60076 532616
rect 57237 532611 57303 532614
rect 282821 532402 282887 532405
rect 279956 532400 282887 532402
rect 279956 532344 282826 532400
rect 282882 532344 282887 532400
rect 279956 532342 282887 532344
rect 282821 532339 282887 532342
rect 57237 530498 57303 530501
rect 57237 530496 60076 530498
rect 57237 530440 57242 530496
rect 57298 530440 60076 530496
rect 57237 530438 60076 530440
rect 57237 530435 57303 530438
rect 282821 530226 282887 530229
rect 279956 530224 282887 530226
rect 279956 530168 282826 530224
rect 282882 530168 282887 530224
rect 279956 530166 282887 530168
rect 282821 530163 282887 530166
rect 57237 528458 57303 528461
rect 57237 528456 60076 528458
rect 57237 528400 57242 528456
rect 57298 528400 60076 528456
rect 57237 528398 60076 528400
rect 57237 528395 57303 528398
rect 282821 527914 282887 527917
rect 279956 527912 282887 527914
rect 279956 527856 282826 527912
rect 282882 527856 282887 527912
rect 279956 527854 282887 527856
rect 282821 527851 282887 527854
rect 57237 526282 57303 526285
rect 57237 526280 60076 526282
rect 57237 526224 57242 526280
rect 57298 526224 60076 526280
rect 57237 526222 60076 526224
rect 57237 526219 57303 526222
rect 282821 525738 282887 525741
rect 279956 525736 282887 525738
rect 279956 525680 282826 525736
rect 282882 525680 282887 525736
rect 279956 525678 282887 525680
rect 282821 525675 282887 525678
rect -960 524092 480 524332
rect 57237 524242 57303 524245
rect 57237 524240 60076 524242
rect 57237 524184 57242 524240
rect 57298 524184 60076 524240
rect 57237 524182 60076 524184
rect 57237 524179 57303 524182
rect 282821 523562 282887 523565
rect 279956 523560 282887 523562
rect 279956 523504 282826 523560
rect 282882 523504 282887 523560
rect 279956 523502 282887 523504
rect 282821 523499 282887 523502
rect 57237 522066 57303 522069
rect 57237 522064 60076 522066
rect 57237 522008 57242 522064
rect 57298 522008 60076 522064
rect 57237 522006 60076 522008
rect 57237 522003 57303 522006
rect 583520 521916 584960 522156
rect 282821 521386 282887 521389
rect 279956 521384 282887 521386
rect 279956 521328 282826 521384
rect 282882 521328 282887 521384
rect 279956 521326 282887 521328
rect 282821 521323 282887 521326
rect 57237 520026 57303 520029
rect 57237 520024 60076 520026
rect 57237 519968 57242 520024
rect 57298 519968 60076 520024
rect 57237 519966 60076 519968
rect 57237 519963 57303 519966
rect 282821 519210 282887 519213
rect 279956 519208 282887 519210
rect 279956 519152 282826 519208
rect 282882 519152 282887 519208
rect 279956 519150 282887 519152
rect 282821 519147 282887 519150
rect 57237 517850 57303 517853
rect 57237 517848 60076 517850
rect 57237 517792 57242 517848
rect 57298 517792 60076 517848
rect 57237 517790 60076 517792
rect 57237 517787 57303 517790
rect 281901 516898 281967 516901
rect 279956 516896 281967 516898
rect 279956 516840 281906 516896
rect 281962 516840 281967 516896
rect 279956 516838 281967 516840
rect 281901 516835 281967 516838
rect 57237 515810 57303 515813
rect 57237 515808 60076 515810
rect 57237 515752 57242 515808
rect 57298 515752 60076 515808
rect 57237 515750 60076 515752
rect 57237 515747 57303 515750
rect 282821 514722 282887 514725
rect 279956 514720 282887 514722
rect 279956 514664 282826 514720
rect 282882 514664 282887 514720
rect 279956 514662 282887 514664
rect 282821 514659 282887 514662
rect 57237 513634 57303 513637
rect 57237 513632 60076 513634
rect 57237 513576 57242 513632
rect 57298 513576 60076 513632
rect 57237 513574 60076 513576
rect 57237 513571 57303 513574
rect 282085 512546 282151 512549
rect 279956 512544 282151 512546
rect 279956 512488 282090 512544
rect 282146 512488 282151 512544
rect 279956 512486 282151 512488
rect 282085 512483 282151 512486
rect 57237 511594 57303 511597
rect 57237 511592 60076 511594
rect 57237 511536 57242 511592
rect 57298 511536 60076 511592
rect 57237 511534 60076 511536
rect 57237 511531 57303 511534
rect 282821 510370 282887 510373
rect 279956 510368 282887 510370
rect 279956 510312 282826 510368
rect 282882 510312 282887 510368
rect 279956 510310 282887 510312
rect 282821 510307 282887 510310
rect 580257 510370 580323 510373
rect 583520 510370 584960 510460
rect 580257 510368 584960 510370
rect 580257 510312 580262 510368
rect 580318 510312 584960 510368
rect 580257 510310 584960 510312
rect 580257 510307 580323 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 2773 509962 2839 509965
rect -960 509960 2839 509962
rect -960 509904 2778 509960
rect 2834 509904 2839 509960
rect -960 509902 2839 509904
rect -960 509812 480 509902
rect 2773 509899 2839 509902
rect 57237 509418 57303 509421
rect 57237 509416 60076 509418
rect 57237 509360 57242 509416
rect 57298 509360 60076 509416
rect 57237 509358 60076 509360
rect 57237 509355 57303 509358
rect 282269 508194 282335 508197
rect 279956 508192 282335 508194
rect 279956 508136 282274 508192
rect 282330 508136 282335 508192
rect 279956 508134 282335 508136
rect 282269 508131 282335 508134
rect 57237 507378 57303 507381
rect 57237 507376 60076 507378
rect 57237 507320 57242 507376
rect 57298 507320 60076 507376
rect 57237 507318 60076 507320
rect 57237 507315 57303 507318
rect 281901 505882 281967 505885
rect 279956 505880 281967 505882
rect 279956 505824 281906 505880
rect 281962 505824 281967 505880
rect 279956 505822 281967 505824
rect 281901 505819 281967 505822
rect 57237 505202 57303 505205
rect 57237 505200 60076 505202
rect 57237 505144 57242 505200
rect 57298 505144 60076 505200
rect 57237 505142 60076 505144
rect 57237 505139 57303 505142
rect 282821 503706 282887 503709
rect 279956 503704 282887 503706
rect 279956 503648 282826 503704
rect 282882 503648 282887 503704
rect 279956 503646 282887 503648
rect 282821 503643 282887 503646
rect 57237 503162 57303 503165
rect 57237 503160 60076 503162
rect 57237 503104 57242 503160
rect 57298 503104 60076 503160
rect 57237 503102 60076 503104
rect 57237 503099 57303 503102
rect 282085 501530 282151 501533
rect 279956 501528 282151 501530
rect 279956 501472 282090 501528
rect 282146 501472 282151 501528
rect 279956 501470 282151 501472
rect 282085 501467 282151 501470
rect 57237 500986 57303 500989
rect 57237 500984 60076 500986
rect 57237 500928 57242 500984
rect 57298 500928 60076 500984
rect 57237 500926 60076 500928
rect 57237 500923 57303 500926
rect 282821 499354 282887 499357
rect 279956 499352 282887 499354
rect 279956 499296 282826 499352
rect 282882 499296 282887 499352
rect 279956 499294 282887 499296
rect 282821 499291 282887 499294
rect 57237 498946 57303 498949
rect 57237 498944 60076 498946
rect 57237 498888 57242 498944
rect 57298 498888 60076 498944
rect 57237 498886 60076 498888
rect 57237 498883 57303 498886
rect 580257 498674 580323 498677
rect 583520 498674 584960 498764
rect 580257 498672 584960 498674
rect 580257 498616 580262 498672
rect 580318 498616 584960 498672
rect 580257 498614 584960 498616
rect 580257 498611 580323 498614
rect 583520 498524 584960 498614
rect 282269 497178 282335 497181
rect 279956 497176 282335 497178
rect 279956 497120 282274 497176
rect 282330 497120 282335 497176
rect 279956 497118 282335 497120
rect 282269 497115 282335 497118
rect 56961 496770 57027 496773
rect 56961 496768 60076 496770
rect 56961 496712 56966 496768
rect 57022 496712 60076 496768
rect 56961 496710 60076 496712
rect 56961 496707 57027 496710
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 281901 494866 281967 494869
rect 279956 494864 281967 494866
rect 279956 494808 281906 494864
rect 281962 494808 281967 494864
rect 279956 494806 281967 494808
rect 281901 494803 281967 494806
rect 57237 494730 57303 494733
rect 57237 494728 60076 494730
rect 57237 494672 57242 494728
rect 57298 494672 60076 494728
rect 57237 494670 60076 494672
rect 57237 494667 57303 494670
rect 282453 492690 282519 492693
rect 279956 492688 282519 492690
rect 279956 492632 282458 492688
rect 282514 492632 282519 492688
rect 279956 492630 282519 492632
rect 282453 492627 282519 492630
rect 57237 492554 57303 492557
rect 57237 492552 60076 492554
rect 57237 492496 57242 492552
rect 57298 492496 60076 492552
rect 57237 492494 60076 492496
rect 57237 492491 57303 492494
rect 56961 490514 57027 490517
rect 282085 490514 282151 490517
rect 56961 490512 60076 490514
rect 56961 490456 56966 490512
rect 57022 490456 60076 490512
rect 56961 490454 60076 490456
rect 279956 490512 282151 490514
rect 279956 490456 282090 490512
rect 282146 490456 282151 490512
rect 279956 490454 282151 490456
rect 56961 490451 57027 490454
rect 282085 490451 282151 490454
rect 56593 488338 56659 488341
rect 282821 488338 282887 488341
rect 56593 488336 60076 488338
rect 56593 488280 56598 488336
rect 56654 488280 60076 488336
rect 56593 488278 60076 488280
rect 279956 488336 282887 488338
rect 279956 488280 282826 488336
rect 282882 488280 282887 488336
rect 279956 488278 282887 488280
rect 56593 488275 56659 488278
rect 282821 488275 282887 488278
rect 578877 486842 578943 486845
rect 583520 486842 584960 486932
rect 578877 486840 584960 486842
rect 578877 486784 578882 486840
rect 578938 486784 584960 486840
rect 578877 486782 584960 486784
rect 578877 486779 578943 486782
rect 583520 486692 584960 486782
rect 56593 486298 56659 486301
rect 56593 486296 60076 486298
rect 56593 486240 56598 486296
rect 56654 486240 60076 486296
rect 56593 486238 60076 486240
rect 56593 486235 56659 486238
rect 282821 486162 282887 486165
rect 279956 486160 282887 486162
rect 279956 486104 282826 486160
rect 282882 486104 282887 486160
rect 279956 486102 282887 486104
rect 282821 486099 282887 486102
rect 56593 484122 56659 484125
rect 56593 484120 60076 484122
rect 56593 484064 56598 484120
rect 56654 484064 60076 484120
rect 56593 484062 60076 484064
rect 56593 484059 56659 484062
rect 282821 483850 282887 483853
rect 279956 483848 282887 483850
rect 279956 483792 282826 483848
rect 282882 483792 282887 483848
rect 279956 483790 282887 483792
rect 282821 483787 282887 483790
rect 56593 482082 56659 482085
rect 56593 482080 60076 482082
rect 56593 482024 56598 482080
rect 56654 482024 60076 482080
rect 56593 482022 60076 482024
rect 56593 482019 56659 482022
rect 282453 481674 282519 481677
rect 279956 481672 282519 481674
rect 279956 481616 282458 481672
rect 282514 481616 282519 481672
rect 279956 481614 282519 481616
rect 282453 481611 282519 481614
rect -960 481130 480 481220
rect 3233 481130 3299 481133
rect -960 481128 3299 481130
rect -960 481072 3238 481128
rect 3294 481072 3299 481128
rect -960 481070 3299 481072
rect -960 480980 480 481070
rect 3233 481067 3299 481070
rect 56593 480042 56659 480045
rect 56593 480040 60076 480042
rect 56593 479984 56598 480040
rect 56654 479984 60076 480040
rect 56593 479982 60076 479984
rect 56593 479979 56659 479982
rect 282085 479498 282151 479501
rect 279956 479496 282151 479498
rect 279956 479440 282090 479496
rect 282146 479440 282151 479496
rect 279956 479438 282151 479440
rect 282085 479435 282151 479438
rect 56593 477866 56659 477869
rect 56593 477864 60076 477866
rect 56593 477808 56598 477864
rect 56654 477808 60076 477864
rect 56593 477806 60076 477808
rect 56593 477803 56659 477806
rect 282821 477322 282887 477325
rect 279956 477320 282887 477322
rect 279956 477264 282826 477320
rect 282882 477264 282887 477320
rect 279956 477262 282887 477264
rect 282821 477259 282887 477262
rect 56593 475826 56659 475829
rect 56593 475824 60076 475826
rect 56593 475768 56598 475824
rect 56654 475768 60076 475824
rect 56593 475766 60076 475768
rect 56593 475763 56659 475766
rect 282545 475146 282611 475149
rect 279956 475144 282611 475146
rect 279956 475088 282550 475144
rect 282606 475088 282611 475144
rect 279956 475086 282611 475088
rect 282545 475083 282611 475086
rect 583520 474996 584960 475236
rect 56593 473650 56659 473653
rect 56593 473648 60076 473650
rect 56593 473592 56598 473648
rect 56654 473592 60076 473648
rect 56593 473590 60076 473592
rect 56593 473587 56659 473590
rect 282085 472970 282151 472973
rect 279956 472968 282151 472970
rect 279956 472912 282090 472968
rect 282146 472912 282151 472968
rect 279956 472910 282151 472912
rect 282085 472907 282151 472910
rect 56593 471610 56659 471613
rect 56593 471608 60076 471610
rect 56593 471552 56598 471608
rect 56654 471552 60076 471608
rect 56593 471550 60076 471552
rect 56593 471547 56659 471550
rect 282453 470658 282519 470661
rect 279956 470656 282519 470658
rect 279956 470600 282458 470656
rect 282514 470600 282519 470656
rect 279956 470598 282519 470600
rect 282453 470595 282519 470598
rect 56501 469978 56567 469981
rect 56501 469976 60106 469978
rect 56501 469920 56506 469976
rect 56562 469920 60106 469976
rect 56501 469918 60106 469920
rect 56501 469915 56567 469918
rect 60046 469404 60106 469918
rect 282085 468482 282151 468485
rect 279956 468480 282151 468482
rect 279956 468424 282090 468480
rect 282146 468424 282151 468480
rect 279956 468422 282151 468424
rect 282085 468419 282151 468422
rect 56501 467802 56567 467805
rect 56501 467800 60106 467802
rect 56501 467744 56506 467800
rect 56562 467744 60106 467800
rect 56501 467742 60106 467744
rect 56501 467739 56567 467742
rect 60046 467364 60106 467742
rect -960 466700 480 466940
rect 282821 466306 282887 466309
rect 279956 466304 282887 466306
rect 279956 466248 282826 466304
rect 282882 466248 282887 466304
rect 279956 466246 282887 466248
rect 282821 466243 282887 466246
rect 56501 465762 56567 465765
rect 56501 465760 60106 465762
rect 56501 465704 56506 465760
rect 56562 465704 60106 465760
rect 56501 465702 60106 465704
rect 56501 465699 56567 465702
rect 60046 465188 60106 465702
rect 282269 464130 282335 464133
rect 279956 464128 282335 464130
rect 279956 464072 282274 464128
rect 282330 464072 282335 464128
rect 279956 464070 282335 464072
rect 282269 464067 282335 464070
rect 56501 463586 56567 463589
rect 56501 463584 60106 463586
rect 56501 463528 56506 463584
rect 56562 463528 60106 463584
rect 56501 463526 60106 463528
rect 56501 463523 56567 463526
rect 60046 463148 60106 463526
rect 579981 463450 580047 463453
rect 583520 463450 584960 463540
rect 579981 463448 584960 463450
rect 579981 463392 579986 463448
rect 580042 463392 584960 463448
rect 579981 463390 584960 463392
rect 579981 463387 580047 463390
rect 583520 463300 584960 463390
rect 282821 461954 282887 461957
rect 279956 461952 282887 461954
rect 279956 461896 282826 461952
rect 282882 461896 282887 461952
rect 279956 461894 282887 461896
rect 282821 461891 282887 461894
rect 56501 461546 56567 461549
rect 56501 461544 60106 461546
rect 56501 461488 56506 461544
rect 56562 461488 60106 461544
rect 56501 461486 60106 461488
rect 56501 461483 56567 461486
rect 60046 460972 60106 461486
rect 282453 459642 282519 459645
rect 279956 459640 282519 459642
rect 279956 459584 282458 459640
rect 282514 459584 282519 459640
rect 279956 459582 282519 459584
rect 282453 459579 282519 459582
rect 56593 458962 56659 458965
rect 56593 458960 60076 458962
rect 56593 458904 56598 458960
rect 56654 458904 60076 458960
rect 56593 458902 60076 458904
rect 56593 458899 56659 458902
rect 282085 457466 282151 457469
rect 279956 457464 282151 457466
rect 279956 457408 282090 457464
rect 282146 457408 282151 457464
rect 279956 457406 282151 457408
rect 282085 457403 282151 457406
rect 56593 456786 56659 456789
rect 56593 456784 60076 456786
rect 56593 456728 56598 456784
rect 56654 456728 60076 456784
rect 56593 456726 60076 456728
rect 56593 456723 56659 456726
rect 282821 455290 282887 455293
rect 279956 455288 282887 455290
rect 279956 455232 282826 455288
rect 282882 455232 282887 455288
rect 279956 455230 282887 455232
rect 282821 455227 282887 455230
rect 56593 454746 56659 454749
rect 56593 454744 60076 454746
rect 56593 454688 56598 454744
rect 56654 454688 60076 454744
rect 56593 454686 60076 454688
rect 56593 454683 56659 454686
rect 282821 453114 282887 453117
rect 279956 453112 282887 453114
rect 279956 453056 282826 453112
rect 282882 453056 282887 453112
rect 279956 453054 282887 453056
rect 282821 453051 282887 453054
rect 56593 452570 56659 452573
rect 56593 452568 60076 452570
rect -960 452434 480 452524
rect 56593 452512 56598 452568
rect 56654 452512 60076 452568
rect 56593 452510 60076 452512
rect 56593 452507 56659 452510
rect 3325 452434 3391 452437
rect -960 452432 3391 452434
rect -960 452376 3330 452432
rect 3386 452376 3391 452432
rect -960 452374 3391 452376
rect -960 452284 480 452374
rect 3325 452371 3391 452374
rect 580257 451754 580323 451757
rect 583520 451754 584960 451844
rect 580257 451752 584960 451754
rect 580257 451696 580262 451752
rect 580318 451696 584960 451752
rect 580257 451694 584960 451696
rect 580257 451691 580323 451694
rect 583520 451604 584960 451694
rect 282821 450938 282887 450941
rect 279956 450936 282887 450938
rect 279956 450880 282826 450936
rect 282882 450880 282887 450936
rect 279956 450878 282887 450880
rect 282821 450875 282887 450878
rect 56593 450530 56659 450533
rect 56593 450528 60076 450530
rect 56593 450472 56598 450528
rect 56654 450472 60076 450528
rect 56593 450470 60076 450472
rect 56593 450467 56659 450470
rect 282453 448626 282519 448629
rect 279956 448624 282519 448626
rect 279956 448568 282458 448624
rect 282514 448568 282519 448624
rect 279956 448566 282519 448568
rect 282453 448563 282519 448566
rect 57513 448354 57579 448357
rect 57513 448352 60076 448354
rect 57513 448296 57518 448352
rect 57574 448296 60076 448352
rect 57513 448294 60076 448296
rect 57513 448291 57579 448294
rect 282821 446450 282887 446453
rect 279956 446448 282887 446450
rect 279956 446392 282826 446448
rect 282882 446392 282887 446448
rect 279956 446390 282887 446392
rect 282821 446387 282887 446390
rect 57513 446314 57579 446317
rect 57513 446312 60076 446314
rect 57513 446256 57518 446312
rect 57574 446256 60076 446312
rect 57513 446254 60076 446256
rect 57513 446251 57579 446254
rect 282821 444274 282887 444277
rect 279956 444272 282887 444274
rect 279956 444216 282826 444272
rect 282882 444216 282887 444272
rect 279956 444214 282887 444216
rect 282821 444211 282887 444214
rect 56593 444138 56659 444141
rect 56593 444136 60076 444138
rect 56593 444080 56598 444136
rect 56654 444080 60076 444136
rect 56593 444078 60076 444080
rect 56593 444075 56659 444078
rect 58433 442098 58499 442101
rect 282821 442098 282887 442101
rect 58433 442096 60076 442098
rect 58433 442040 58438 442096
rect 58494 442040 60076 442096
rect 58433 442038 60076 442040
rect 279956 442096 282887 442098
rect 279956 442040 282826 442096
rect 282882 442040 282887 442096
rect 279956 442038 282887 442040
rect 58433 442035 58499 442038
rect 282821 442035 282887 442038
rect 57421 439922 57487 439925
rect 282821 439922 282887 439925
rect 57421 439920 60076 439922
rect 57421 439864 57426 439920
rect 57482 439864 60076 439920
rect 57421 439862 60076 439864
rect 279956 439920 282887 439922
rect 279956 439864 282826 439920
rect 282882 439864 282887 439920
rect 279956 439862 282887 439864
rect 57421 439859 57487 439862
rect 282821 439859 282887 439862
rect 579613 439922 579679 439925
rect 583520 439922 584960 440012
rect 579613 439920 584960 439922
rect 579613 439864 579618 439920
rect 579674 439864 584960 439920
rect 579613 439862 584960 439864
rect 579613 439859 579679 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 4061 438018 4127 438021
rect -960 438016 4127 438018
rect -960 437960 4066 438016
rect 4122 437960 4127 438016
rect -960 437958 4127 437960
rect -960 437868 480 437958
rect 4061 437955 4127 437958
rect 57605 437882 57671 437885
rect 57605 437880 60076 437882
rect 57605 437824 57610 437880
rect 57666 437824 60076 437880
rect 57605 437822 60076 437824
rect 57605 437819 57671 437822
rect 282453 437610 282519 437613
rect 279956 437608 282519 437610
rect 279956 437552 282458 437608
rect 282514 437552 282519 437608
rect 279956 437550 282519 437552
rect 282453 437547 282519 437550
rect 58525 435706 58591 435709
rect 58525 435704 60076 435706
rect 58525 435648 58530 435704
rect 58586 435648 60076 435704
rect 58525 435646 60076 435648
rect 58525 435643 58591 435646
rect 282821 435434 282887 435437
rect 279956 435432 282887 435434
rect 279956 435376 282826 435432
rect 282882 435376 282887 435432
rect 279956 435374 282887 435376
rect 282821 435371 282887 435374
rect 56685 433666 56751 433669
rect 56685 433664 60076 433666
rect 56685 433608 56690 433664
rect 56746 433608 60076 433664
rect 56685 433606 60076 433608
rect 56685 433603 56751 433606
rect 282821 433258 282887 433261
rect 279956 433256 282887 433258
rect 279956 433200 282826 433256
rect 282882 433200 282887 433256
rect 279956 433198 282887 433200
rect 282821 433195 282887 433198
rect 58709 431490 58775 431493
rect 58709 431488 60076 431490
rect 58709 431432 58714 431488
rect 58770 431432 60076 431488
rect 58709 431430 60076 431432
rect 58709 431427 58775 431430
rect 282821 431082 282887 431085
rect 279956 431080 282887 431082
rect 279956 431024 282826 431080
rect 282882 431024 282887 431080
rect 279956 431022 282887 431024
rect 282821 431019 282887 431022
rect 58801 429450 58867 429453
rect 58801 429448 60076 429450
rect 58801 429392 58806 429448
rect 58862 429392 60076 429448
rect 58801 429390 60076 429392
rect 58801 429387 58867 429390
rect 282821 428906 282887 428909
rect 279956 428904 282887 428906
rect 279956 428848 282826 428904
rect 282882 428848 282887 428904
rect 279956 428846 282887 428848
rect 282821 428843 282887 428846
rect 583520 428076 584960 428316
rect 56777 427274 56843 427277
rect 56777 427272 60076 427274
rect 56777 427216 56782 427272
rect 56838 427216 60076 427272
rect 56777 427214 60076 427216
rect 56777 427211 56843 427214
rect 282821 426594 282887 426597
rect 279956 426592 282887 426594
rect 279956 426536 282826 426592
rect 282882 426536 282887 426592
rect 279956 426534 282887 426536
rect 282821 426531 282887 426534
rect 58893 425234 58959 425237
rect 58893 425232 60076 425234
rect 58893 425176 58898 425232
rect 58954 425176 60076 425232
rect 58893 425174 60076 425176
rect 58893 425171 58959 425174
rect 282453 424418 282519 424421
rect 279956 424416 282519 424418
rect 279956 424360 282458 424416
rect 282514 424360 282519 424416
rect 279956 424358 282519 424360
rect 282453 424355 282519 424358
rect -960 423738 480 423828
rect 3969 423738 4035 423741
rect -960 423736 4035 423738
rect -960 423680 3974 423736
rect 4030 423680 4035 423736
rect -960 423678 4035 423680
rect -960 423588 480 423678
rect 3969 423675 4035 423678
rect 58985 423058 59051 423061
rect 58985 423056 60076 423058
rect 58985 423000 58990 423056
rect 59046 423000 60076 423056
rect 58985 422998 60076 423000
rect 58985 422995 59051 422998
rect 282085 422242 282151 422245
rect 279956 422240 282151 422242
rect 279956 422184 282090 422240
rect 282146 422184 282151 422240
rect 279956 422182 282151 422184
rect 282085 422179 282151 422182
rect 56869 421018 56935 421021
rect 56869 421016 60076 421018
rect 56869 420960 56874 421016
rect 56930 420960 60076 421016
rect 56869 420958 60076 420960
rect 56869 420955 56935 420958
rect 281717 420066 281783 420069
rect 279956 420064 281783 420066
rect 279956 420008 281722 420064
rect 281778 420008 281783 420064
rect 279956 420006 281783 420008
rect 281717 420003 281783 420006
rect 57697 418978 57763 418981
rect 57697 418976 60076 418978
rect 57697 418920 57702 418976
rect 57758 418920 60076 418976
rect 57697 418918 60076 418920
rect 57697 418915 57763 418918
rect 282821 417890 282887 417893
rect 279956 417888 282887 417890
rect 279956 417832 282826 417888
rect 282882 417832 282887 417888
rect 279956 417830 282887 417832
rect 282821 417827 282887 417830
rect 59077 416802 59143 416805
rect 59077 416800 60076 416802
rect 59077 416744 59082 416800
rect 59138 416744 60076 416800
rect 59077 416742 60076 416744
rect 59077 416739 59143 416742
rect 580257 416530 580323 416533
rect 583520 416530 584960 416620
rect 580257 416528 584960 416530
rect 580257 416472 580262 416528
rect 580318 416472 584960 416528
rect 580257 416470 584960 416472
rect 580257 416467 580323 416470
rect 583520 416380 584960 416470
rect 282821 415714 282887 415717
rect 279956 415712 282887 415714
rect 279956 415656 282826 415712
rect 282882 415656 282887 415712
rect 279956 415654 282887 415656
rect 282821 415651 282887 415654
rect 59537 414762 59603 414765
rect 59537 414760 60076 414762
rect 59537 414704 59542 414760
rect 59598 414704 60076 414760
rect 59537 414702 60076 414704
rect 59537 414699 59603 414702
rect 281901 413402 281967 413405
rect 279956 413400 281967 413402
rect 279956 413344 281906 413400
rect 281962 413344 281967 413400
rect 279956 413342 281967 413344
rect 281901 413339 281967 413342
rect 57789 412586 57855 412589
rect 57789 412584 60076 412586
rect 57789 412528 57794 412584
rect 57850 412528 60076 412584
rect 57789 412526 60076 412528
rect 57789 412523 57855 412526
rect 282821 411226 282887 411229
rect 279956 411224 282887 411226
rect 279956 411168 282826 411224
rect 282882 411168 282887 411224
rect 279956 411166 282887 411168
rect 282821 411163 282887 411166
rect 59169 410546 59235 410549
rect 59169 410544 60076 410546
rect 59169 410488 59174 410544
rect 59230 410488 60076 410544
rect 59169 410486 60076 410488
rect 59169 410483 59235 410486
rect -960 409172 480 409412
rect 282085 409050 282151 409053
rect 279956 409048 282151 409050
rect 279956 408992 282090 409048
rect 282146 408992 282151 409048
rect 279956 408990 282151 408992
rect 282085 408987 282151 408990
rect 59721 408370 59787 408373
rect 59721 408368 60076 408370
rect 59721 408312 59726 408368
rect 59782 408312 60076 408368
rect 59721 408310 60076 408312
rect 59721 408307 59787 408310
rect 282821 406874 282887 406877
rect 279956 406872 282887 406874
rect 279956 406816 282826 406872
rect 282882 406816 282887 406872
rect 279956 406814 282887 406816
rect 282821 406811 282887 406814
rect 57881 406330 57947 406333
rect 57881 406328 60076 406330
rect 57881 406272 57886 406328
rect 57942 406272 60076 406328
rect 57881 406270 60076 406272
rect 57881 406267 57947 406270
rect 580901 404834 580967 404837
rect 583520 404834 584960 404924
rect 580901 404832 584960 404834
rect 580901 404776 580906 404832
rect 580962 404776 584960 404832
rect 580901 404774 584960 404776
rect 580901 404771 580967 404774
rect 282821 404698 282887 404701
rect 279956 404696 282887 404698
rect 279956 404640 282826 404696
rect 282882 404640 282887 404696
rect 583520 404684 584960 404774
rect 279956 404638 282887 404640
rect 282821 404635 282887 404638
rect 58341 404154 58407 404157
rect 58341 404152 60076 404154
rect 58341 404096 58346 404152
rect 58402 404096 60076 404152
rect 58341 404094 60076 404096
rect 58341 404091 58407 404094
rect 281901 402386 281967 402389
rect 279956 402384 281967 402386
rect 279956 402328 281906 402384
rect 281962 402328 281967 402384
rect 279956 402326 281967 402328
rect 281901 402323 281967 402326
rect 59445 402114 59511 402117
rect 59445 402112 60076 402114
rect 59445 402056 59450 402112
rect 59506 402056 60076 402112
rect 59445 402054 60076 402056
rect 59445 402051 59511 402054
rect 282821 400210 282887 400213
rect 279956 400208 282887 400210
rect 279956 400152 282826 400208
rect 282882 400152 282887 400208
rect 279956 400150 282887 400152
rect 282821 400147 282887 400150
rect 59353 399938 59419 399941
rect 59353 399936 60076 399938
rect 59353 399880 59358 399936
rect 59414 399880 60076 399936
rect 59353 399878 60076 399880
rect 59353 399875 59419 399878
rect 282085 398034 282151 398037
rect 279956 398032 282151 398034
rect 279956 397976 282090 398032
rect 282146 397976 282151 398032
rect 279956 397974 282151 397976
rect 282085 397971 282151 397974
rect 59261 397898 59327 397901
rect 59261 397896 60076 397898
rect 59261 397840 59266 397896
rect 59322 397840 60076 397896
rect 59261 397838 60076 397840
rect 59261 397835 59327 397838
rect 282085 395858 282151 395861
rect 279956 395856 282151 395858
rect 279956 395800 282090 395856
rect 282146 395800 282151 395856
rect 279956 395798 282151 395800
rect 282085 395795 282151 395798
rect 59629 395722 59695 395725
rect 59629 395720 60076 395722
rect 59629 395664 59634 395720
rect 59690 395664 60076 395720
rect 59629 395662 60076 395664
rect 59629 395659 59695 395662
rect -960 395042 480 395132
rect 3785 395042 3851 395045
rect -960 395040 3851 395042
rect -960 394984 3790 395040
rect 3846 394984 3851 395040
rect -960 394982 3851 394984
rect -960 394892 480 394982
rect 3785 394979 3851 394982
rect 57830 393620 57836 393684
rect 57900 393682 57906 393684
rect 282269 393682 282335 393685
rect 57900 393622 60076 393682
rect 279956 393680 282335 393682
rect 279956 393624 282274 393680
rect 282330 393624 282335 393680
rect 279956 393622 282335 393624
rect 57900 393620 57906 393622
rect 282269 393619 282335 393622
rect 579613 393002 579679 393005
rect 583520 393002 584960 393092
rect 579613 393000 584960 393002
rect 579613 392944 579618 393000
rect 579674 392944 584960 393000
rect 579613 392942 584960 392944
rect 579613 392939 579679 392942
rect 583520 392852 584960 392942
rect 59118 391444 59124 391508
rect 59188 391506 59194 391508
rect 59188 391446 60076 391506
rect 59188 391444 59194 391446
rect 281901 391370 281967 391373
rect 279956 391368 281967 391370
rect 279956 391312 281906 391368
rect 281962 391312 281967 391368
rect 279956 391310 281967 391312
rect 281901 391307 281967 391310
rect 58198 389404 58204 389468
rect 58268 389466 58274 389468
rect 58268 389406 60076 389466
rect 58268 389404 58274 389406
rect 282453 389194 282519 389197
rect 279956 389192 282519 389194
rect 279956 389136 282458 389192
rect 282514 389136 282519 389192
rect 279956 389134 282519 389136
rect 282453 389131 282519 389134
rect 57462 387228 57468 387292
rect 57532 387290 57538 387292
rect 57532 387230 60076 387290
rect 57532 387228 57538 387230
rect 282085 387018 282151 387021
rect 279956 387016 282151 387018
rect 279956 386960 282090 387016
rect 282146 386960 282151 387016
rect 279956 386958 282151 386960
rect 282085 386955 282151 386958
rect 58617 385250 58683 385253
rect 58617 385248 60076 385250
rect 58617 385192 58622 385248
rect 58678 385192 60076 385248
rect 58617 385190 60076 385192
rect 58617 385187 58683 385190
rect 282821 384842 282887 384845
rect 279956 384840 282887 384842
rect 279956 384784 282826 384840
rect 282882 384784 282887 384840
rect 279956 384782 282887 384784
rect 282821 384779 282887 384782
rect 57973 383074 58039 383077
rect 57973 383072 60076 383074
rect 57973 383016 57978 383072
rect 58034 383016 60076 383072
rect 57973 383014 60076 383016
rect 57973 383011 58039 383014
rect 282821 382666 282887 382669
rect 279956 382664 282887 382666
rect 279956 382608 282826 382664
rect 282882 382608 282887 382664
rect 279956 382606 282887 382608
rect 282821 382603 282887 382606
rect 583520 381156 584960 381396
rect 57053 381034 57119 381037
rect 57053 381032 60076 381034
rect 57053 380976 57058 381032
rect 57114 380976 60076 381032
rect 57053 380974 60076 380976
rect 57053 380971 57119 380974
rect -960 380626 480 380716
rect 3693 380626 3759 380629
rect -960 380624 3759 380626
rect -960 380568 3698 380624
rect 3754 380568 3759 380624
rect -960 380566 3759 380568
rect -960 380476 480 380566
rect 3693 380563 3759 380566
rect 282821 380354 282887 380357
rect 279956 380352 282887 380354
rect 279956 380296 282826 380352
rect 282882 380296 282887 380352
rect 279956 380294 282887 380296
rect 282821 380291 282887 380294
rect 57646 378796 57652 378860
rect 57716 378858 57722 378860
rect 57716 378798 60076 378858
rect 57716 378796 57722 378798
rect 282453 378178 282519 378181
rect 279956 378176 282519 378178
rect 279956 378120 282458 378176
rect 282514 378120 282519 378176
rect 279956 378118 282519 378120
rect 282453 378115 282519 378118
rect 58065 376818 58131 376821
rect 58065 376816 60076 376818
rect 58065 376760 58070 376816
rect 58126 376760 60076 376816
rect 58065 376758 60076 376760
rect 58065 376755 58131 376758
rect 282085 376002 282151 376005
rect 279956 376000 282151 376002
rect 279956 375944 282090 376000
rect 282146 375944 282151 376000
rect 279956 375942 282151 375944
rect 282085 375939 282151 375942
rect 57329 374642 57395 374645
rect 57329 374640 60076 374642
rect 57329 374584 57334 374640
rect 57390 374584 60076 374640
rect 57329 374582 60076 374584
rect 57329 374579 57395 374582
rect 282821 373826 282887 373829
rect 279956 373824 282887 373826
rect 279956 373768 282826 373824
rect 282882 373768 282887 373824
rect 279956 373766 282887 373768
rect 282821 373763 282887 373766
rect 58249 372602 58315 372605
rect 58249 372600 60076 372602
rect 58249 372544 58254 372600
rect 58310 372544 60076 372600
rect 58249 372542 60076 372544
rect 58249 372539 58315 372542
rect 282545 371650 282611 371653
rect 279956 371648 282611 371650
rect 279956 371592 282550 371648
rect 282606 371592 282611 371648
rect 279956 371590 282611 371592
rect 282545 371587 282611 371590
rect 58157 370426 58223 370429
rect 58157 370424 60076 370426
rect 58157 370368 58162 370424
rect 58218 370368 60076 370424
rect 58157 370366 60076 370368
rect 58157 370363 58223 370366
rect 579521 369610 579587 369613
rect 583520 369610 584960 369700
rect 579521 369608 584960 369610
rect 579521 369552 579526 369608
rect 579582 369552 584960 369608
rect 579521 369550 584960 369552
rect 579521 369547 579587 369550
rect 583520 369460 584960 369550
rect 282821 369338 282887 369341
rect 279956 369336 282887 369338
rect 279956 369280 282826 369336
rect 282882 369280 282887 369336
rect 279956 369278 282887 369280
rect 282821 369275 282887 369278
rect 57605 368386 57671 368389
rect 57605 368384 60076 368386
rect 57605 368328 57610 368384
rect 57666 368328 60076 368384
rect 57605 368326 60076 368328
rect 57605 368323 57671 368326
rect 282453 367162 282519 367165
rect 279956 367160 282519 367162
rect 279956 367104 282458 367160
rect 282514 367104 282519 367160
rect 279956 367102 282519 367104
rect 282453 367099 282519 367102
rect -960 366210 480 366300
rect 2957 366210 3023 366213
rect -960 366208 3023 366210
rect -960 366152 2962 366208
rect 3018 366152 3023 366208
rect -960 366150 3023 366152
rect -960 366060 480 366150
rect 2957 366147 3023 366150
rect 57145 366210 57211 366213
rect 57145 366208 60076 366210
rect 57145 366152 57150 366208
rect 57206 366152 60076 366208
rect 57145 366150 60076 366152
rect 57145 366147 57211 366150
rect 282085 364986 282151 364989
rect 279956 364984 282151 364986
rect 279956 364928 282090 364984
rect 282146 364928 282151 364984
rect 279956 364926 282151 364928
rect 282085 364923 282151 364926
rect 57697 364170 57763 364173
rect 57697 364168 60076 364170
rect 57697 364112 57702 364168
rect 57758 364112 60076 364168
rect 57697 364110 60076 364112
rect 57697 364107 57763 364110
rect 282821 362810 282887 362813
rect 279956 362808 282887 362810
rect 279956 362752 282826 362808
rect 282882 362752 282887 362808
rect 279956 362750 282887 362752
rect 282821 362747 282887 362750
rect 57053 361994 57119 361997
rect 57053 361992 60076 361994
rect 57053 361936 57058 361992
rect 57114 361936 60076 361992
rect 57053 361934 60076 361936
rect 57053 361931 57119 361934
rect 282545 360634 282611 360637
rect 279956 360632 282611 360634
rect 279956 360576 282550 360632
rect 282606 360576 282611 360632
rect 279956 360574 282611 360576
rect 282545 360571 282611 360574
rect 57697 359954 57763 359957
rect 57697 359952 60076 359954
rect 57697 359896 57702 359952
rect 57758 359896 60076 359952
rect 57697 359894 60076 359896
rect 57697 359891 57763 359894
rect 282821 358458 282887 358461
rect 279956 358456 282887 358458
rect 279956 358400 282826 358456
rect 282882 358400 282887 358456
rect 279956 358398 282887 358400
rect 282821 358395 282887 358398
rect 57421 357914 57487 357917
rect 579521 357914 579587 357917
rect 583520 357914 584960 358004
rect 57421 357912 60076 357914
rect 57421 357856 57426 357912
rect 57482 357856 60076 357912
rect 57421 357854 60076 357856
rect 579521 357912 584960 357914
rect 579521 357856 579526 357912
rect 579582 357856 584960 357912
rect 579521 357854 584960 357856
rect 57421 357851 57487 357854
rect 579521 357851 579587 357854
rect 583520 357764 584960 357854
rect 282453 356146 282519 356149
rect 279956 356144 282519 356146
rect 279956 356088 282458 356144
rect 282514 356088 282519 356144
rect 279956 356086 282519 356088
rect 282453 356083 282519 356086
rect 57145 355738 57211 355741
rect 57145 355736 60076 355738
rect 57145 355680 57150 355736
rect 57206 355680 60076 355736
rect 57145 355678 60076 355680
rect 57145 355675 57211 355678
rect 282085 353970 282151 353973
rect 279956 353968 282151 353970
rect 279956 353912 282090 353968
rect 282146 353912 282151 353968
rect 279956 353910 282151 353912
rect 282085 353907 282151 353910
rect 56593 353698 56659 353701
rect 56593 353696 60076 353698
rect 56593 353640 56598 353696
rect 56654 353640 60076 353696
rect 56593 353638 60076 353640
rect 56593 353635 56659 353638
rect -960 351780 480 352020
rect 282821 351794 282887 351797
rect 279956 351792 282887 351794
rect 279956 351736 282826 351792
rect 282882 351736 282887 351792
rect 279956 351734 282887 351736
rect 282821 351731 282887 351734
rect 57513 351522 57579 351525
rect 57513 351520 60076 351522
rect 57513 351464 57518 351520
rect 57574 351464 60076 351520
rect 57513 351462 60076 351464
rect 57513 351459 57579 351462
rect 282545 349618 282611 349621
rect 279956 349616 282611 349618
rect 279956 349560 282550 349616
rect 282606 349560 282611 349616
rect 279956 349558 282611 349560
rect 282545 349555 282611 349558
rect 57329 349482 57395 349485
rect 57329 349480 60076 349482
rect 57329 349424 57334 349480
rect 57390 349424 60076 349480
rect 57329 349422 60076 349424
rect 57329 349419 57395 349422
rect 282821 347442 282887 347445
rect 279956 347440 282887 347442
rect 279956 347384 282826 347440
rect 282882 347384 282887 347440
rect 279956 347382 282887 347384
rect 282821 347379 282887 347382
rect 57789 347306 57855 347309
rect 57789 347304 60076 347306
rect 57789 347248 57794 347304
rect 57850 347248 60076 347304
rect 57789 347246 60076 347248
rect 57789 347243 57855 347246
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 57605 345266 57671 345269
rect 57605 345264 60076 345266
rect 57605 345208 57610 345264
rect 57666 345208 60076 345264
rect 57605 345206 60076 345208
rect 57605 345203 57671 345206
rect 282453 345130 282519 345133
rect 279956 345128 282519 345130
rect 279956 345072 282458 345128
rect 282514 345072 282519 345128
rect 279956 345070 282519 345072
rect 282453 345067 282519 345070
rect 56685 343090 56751 343093
rect 56685 343088 60076 343090
rect 56685 343032 56690 343088
rect 56746 343032 60076 343088
rect 56685 343030 60076 343032
rect 56685 343027 56751 343030
rect 282821 342954 282887 342957
rect 279956 342952 282887 342954
rect 279956 342896 282826 342952
rect 282882 342896 282887 342952
rect 279956 342894 282887 342896
rect 282821 342891 282887 342894
rect 57881 341050 57947 341053
rect 57881 341048 60076 341050
rect 57881 340992 57886 341048
rect 57942 340992 60076 341048
rect 57881 340990 60076 340992
rect 57881 340987 57947 340990
rect 282821 340778 282887 340781
rect 279956 340776 282887 340778
rect 279956 340720 282826 340776
rect 282882 340720 282887 340776
rect 279956 340718 282887 340720
rect 282821 340715 282887 340718
rect 56777 338874 56843 338877
rect 56777 338872 60076 338874
rect 56777 338816 56782 338872
rect 56838 338816 60076 338872
rect 56777 338814 60076 338816
rect 56777 338811 56843 338814
rect 282821 338602 282887 338605
rect 279956 338600 282887 338602
rect 279956 338544 282826 338600
rect 282882 338544 282887 338600
rect 279956 338542 282887 338544
rect 282821 338539 282887 338542
rect -960 337514 480 337604
rect 3325 337514 3391 337517
rect -960 337512 3391 337514
rect -960 337456 3330 337512
rect 3386 337456 3391 337512
rect -960 337454 3391 337456
rect -960 337364 480 337454
rect 3325 337451 3391 337454
rect 56961 336834 57027 336837
rect 56961 336832 60076 336834
rect 56961 336776 56966 336832
rect 57022 336776 60076 336832
rect 56961 336774 60076 336776
rect 56961 336771 57027 336774
rect 282821 336426 282887 336429
rect 279956 336424 282887 336426
rect 279956 336368 282826 336424
rect 282882 336368 282887 336424
rect 279956 336366 282887 336368
rect 282821 336363 282887 336366
rect 56869 334658 56935 334661
rect 56869 334656 60076 334658
rect 56869 334600 56874 334656
rect 56930 334600 60076 334656
rect 56869 334598 60076 334600
rect 56869 334595 56935 334598
rect 583520 334236 584960 334476
rect 282361 334114 282427 334117
rect 279956 334112 282427 334114
rect 279956 334056 282366 334112
rect 282422 334056 282427 334112
rect 279956 334054 282427 334056
rect 282361 334051 282427 334054
rect 57053 332618 57119 332621
rect 57053 332616 60076 332618
rect 57053 332560 57058 332616
rect 57114 332560 60076 332616
rect 57053 332558 60076 332560
rect 57053 332555 57119 332558
rect 282821 331938 282887 331941
rect 279956 331936 282887 331938
rect 279956 331880 282826 331936
rect 282882 331880 282887 331936
rect 279956 331878 282887 331880
rect 282821 331875 282887 331878
rect 57329 330442 57395 330445
rect 57329 330440 60076 330442
rect 57329 330384 57334 330440
rect 57390 330384 60076 330440
rect 57329 330382 60076 330384
rect 57329 330379 57395 330382
rect 282821 329762 282887 329765
rect 279956 329760 282887 329762
rect 279956 329704 282826 329760
rect 282882 329704 282887 329760
rect 279956 329702 282887 329704
rect 282821 329699 282887 329702
rect 57145 328402 57211 328405
rect 57145 328400 60076 328402
rect 57145 328344 57150 328400
rect 57206 328344 60076 328400
rect 57145 328342 60076 328344
rect 57145 328339 57211 328342
rect 282821 327586 282887 327589
rect 279956 327584 282887 327586
rect 279956 327528 282826 327584
rect 282882 327528 282887 327584
rect 279956 327526 282887 327528
rect 282821 327523 282887 327526
rect 57421 326226 57487 326229
rect 57421 326224 60076 326226
rect 57421 326168 57426 326224
rect 57482 326168 60076 326224
rect 57421 326166 60076 326168
rect 57421 326163 57487 326166
rect 282821 325410 282887 325413
rect 279956 325408 282887 325410
rect 279956 325352 282826 325408
rect 282882 325352 282887 325408
rect 279956 325350 282887 325352
rect 282821 325347 282887 325350
rect 57697 324186 57763 324189
rect 57697 324184 60076 324186
rect 57697 324128 57702 324184
rect 57758 324128 60076 324184
rect 57697 324126 60076 324128
rect 57697 324123 57763 324126
rect -960 323098 480 323188
rect 3049 323098 3115 323101
rect 282361 323098 282427 323101
rect -960 323096 3115 323098
rect -960 323040 3054 323096
rect 3110 323040 3115 323096
rect -960 323038 3115 323040
rect 279956 323096 282427 323098
rect 279956 323040 282366 323096
rect 282422 323040 282427 323096
rect 279956 323038 282427 323040
rect -960 322948 480 323038
rect 3049 323035 3115 323038
rect 282361 323035 282427 323038
rect 580257 322690 580323 322693
rect 583520 322690 584960 322780
rect 580257 322688 584960 322690
rect 580257 322632 580262 322688
rect 580318 322632 584960 322688
rect 580257 322630 584960 322632
rect 580257 322627 580323 322630
rect 583520 322540 584960 322630
rect 57789 322010 57855 322013
rect 57789 322008 60076 322010
rect 57789 321952 57794 322008
rect 57850 321952 60076 322008
rect 57789 321950 60076 321952
rect 57789 321947 57855 321950
rect 282821 320922 282887 320925
rect 279956 320920 282887 320922
rect 279956 320864 282826 320920
rect 282882 320864 282887 320920
rect 279956 320862 282887 320864
rect 282821 320859 282887 320862
rect 59353 319970 59419 319973
rect 59353 319968 60076 319970
rect 59353 319912 59358 319968
rect 59414 319912 60076 319968
rect 59353 319910 60076 319912
rect 59353 319907 59419 319910
rect 282821 318746 282887 318749
rect 279956 318744 282887 318746
rect 279956 318688 282826 318744
rect 282882 318688 282887 318744
rect 279956 318686 282887 318688
rect 282821 318683 282887 318686
rect 57789 317794 57855 317797
rect 57789 317792 60076 317794
rect 57789 317736 57794 317792
rect 57850 317736 60076 317792
rect 57789 317734 60076 317736
rect 57789 317731 57855 317734
rect 282821 316570 282887 316573
rect 279956 316568 282887 316570
rect 279956 316512 282826 316568
rect 282882 316512 282887 316568
rect 279956 316510 282887 316512
rect 282821 316507 282887 316510
rect 57329 316028 57395 316029
rect 57278 316026 57284 316028
rect 57238 315966 57284 316026
rect 57348 316024 57395 316028
rect 57390 315968 57395 316024
rect 57278 315964 57284 315966
rect 57348 315964 57395 315968
rect 57329 315963 57395 315964
rect 57697 315754 57763 315757
rect 57697 315752 60076 315754
rect 57697 315696 57702 315752
rect 57758 315696 60076 315752
rect 57697 315694 60076 315696
rect 57697 315691 57763 315694
rect 282821 314394 282887 314397
rect 279956 314392 282887 314394
rect 279956 314336 282826 314392
rect 282882 314336 282887 314392
rect 279956 314334 282887 314336
rect 282821 314331 282887 314334
rect 59077 313578 59143 313581
rect 59077 313576 60076 313578
rect 59077 313520 59082 313576
rect 59138 313520 60076 313576
rect 59077 313518 60076 313520
rect 59077 313515 59143 313518
rect 282361 312082 282427 312085
rect 279956 312080 282427 312082
rect 279956 312024 282366 312080
rect 282422 312024 282427 312080
rect 279956 312022 282427 312024
rect 282361 312019 282427 312022
rect 57462 311476 57468 311540
rect 57532 311538 57538 311540
rect 57532 311478 60076 311538
rect 57532 311476 57538 311478
rect 580349 310858 580415 310861
rect 583520 310858 584960 310948
rect 580349 310856 584960 310858
rect 580349 310800 580354 310856
rect 580410 310800 584960 310856
rect 580349 310798 584960 310800
rect 580349 310795 580415 310798
rect 583520 310708 584960 310798
rect 281901 309906 281967 309909
rect 279956 309904 281967 309906
rect 279956 309848 281906 309904
rect 281962 309848 281967 309904
rect 279956 309846 281967 309848
rect 281901 309843 281967 309846
rect 56593 309362 56659 309365
rect 56593 309360 60076 309362
rect 56593 309304 56598 309360
rect 56654 309304 60076 309360
rect 56593 309302 60076 309304
rect 56593 309299 56659 309302
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 282821 307730 282887 307733
rect 279956 307728 282887 307730
rect 279956 307672 282826 307728
rect 282882 307672 282887 307728
rect 279956 307670 282887 307672
rect 282821 307667 282887 307670
rect 59169 307322 59235 307325
rect 59169 307320 60076 307322
rect 59169 307264 59174 307320
rect 59230 307264 60076 307320
rect 59169 307262 60076 307264
rect 59169 307259 59235 307262
rect 57329 306508 57395 306509
rect 57278 306444 57284 306508
rect 57348 306506 57395 306508
rect 57348 306504 57440 306506
rect 57390 306448 57440 306504
rect 57348 306446 57440 306448
rect 57348 306444 57395 306446
rect 57329 306443 57395 306444
rect 282085 305554 282151 305557
rect 279956 305552 282151 305554
rect 279956 305496 282090 305552
rect 282146 305496 282151 305552
rect 279956 305494 282151 305496
rect 282085 305491 282151 305494
rect 57830 305084 57836 305148
rect 57900 305146 57906 305148
rect 57900 305086 60076 305146
rect 57900 305084 57906 305086
rect 281533 303378 281599 303381
rect 279956 303376 281599 303378
rect 279956 303320 281538 303376
rect 281594 303320 281599 303376
rect 279956 303318 281599 303320
rect 281533 303315 281599 303318
rect 57646 303044 57652 303108
rect 57716 303106 57722 303108
rect 57716 303046 60076 303106
rect 57716 303044 57722 303046
rect 281625 301202 281691 301205
rect 279956 301200 281691 301202
rect 279956 301144 281630 301200
rect 281686 301144 281691 301200
rect 279956 301142 281691 301144
rect 281625 301139 281691 301142
rect 59261 301066 59327 301069
rect 59261 301064 60076 301066
rect 59261 301008 59266 301064
rect 59322 301008 60076 301064
rect 59261 301006 60076 301008
rect 59261 301003 59327 301006
rect 60825 300658 60891 300661
rect 61142 300658 61148 300660
rect 60825 300656 61148 300658
rect 60825 300600 60830 300656
rect 60886 300600 61148 300656
rect 60825 300598 61148 300600
rect 60825 300595 60891 300598
rect 61142 300596 61148 300598
rect 61212 300658 61218 300660
rect 61694 300658 61700 300660
rect 61212 300598 61700 300658
rect 61212 300596 61218 300598
rect 61694 300596 61700 300598
rect 61764 300596 61770 300660
rect 61101 299572 61167 299573
rect 61101 299568 61148 299572
rect 61212 299570 61218 299572
rect 61101 299512 61106 299568
rect 61101 299508 61148 299512
rect 61212 299510 61258 299570
rect 61212 299508 61218 299510
rect 61101 299507 61167 299508
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 115841 297666 115907 297669
rect 247769 297666 247835 297669
rect 115841 297664 247835 297666
rect 115841 297608 115846 297664
rect 115902 297608 247774 297664
rect 247830 297608 247835 297664
rect 115841 297606 247835 297608
rect 115841 297603 115907 297606
rect 247769 297603 247835 297606
rect 121361 297530 121427 297533
rect 257521 297530 257587 297533
rect 121361 297528 257587 297530
rect 121361 297472 121366 297528
rect 121422 297472 257526 297528
rect 257582 297472 257587 297528
rect 121361 297470 257587 297472
rect 121361 297467 121427 297470
rect 257521 297467 257587 297470
rect 122741 297394 122807 297397
rect 259453 297394 259519 297397
rect 122741 297392 259519 297394
rect 122741 297336 122746 297392
rect 122802 297336 259458 297392
rect 259514 297336 259519 297392
rect 122741 297334 259519 297336
rect 122741 297331 122807 297334
rect 259453 297331 259519 297334
rect 56777 296714 56843 296717
rect 57605 296714 57671 296717
rect 56777 296712 57671 296714
rect 56777 296656 56782 296712
rect 56838 296656 57610 296712
rect 57666 296656 57671 296712
rect 56777 296654 57671 296656
rect 56777 296651 56843 296654
rect 57605 296651 57671 296654
rect -960 294402 480 294492
rect 2957 294402 3023 294405
rect -960 294400 3023 294402
rect -960 294344 2962 294400
rect 3018 294344 3023 294400
rect -960 294342 3023 294344
rect -960 294252 480 294342
rect 2957 294339 3023 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3325 280122 3391 280125
rect -960 280120 3391 280122
rect -960 280064 3330 280120
rect 3386 280064 3391 280120
rect -960 280062 3391 280064
rect -960 279972 480 280062
rect 3325 280059 3391 280062
rect 56777 277402 56843 277405
rect 57329 277402 57395 277405
rect 56777 277400 57395 277402
rect 56777 277344 56782 277400
rect 56838 277344 57334 277400
rect 57390 277344 57395 277400
rect 56777 277342 57395 277344
rect 56777 277339 56843 277342
rect 57329 277339 57395 277342
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 3141 265706 3207 265709
rect -960 265704 3207 265706
rect -960 265648 3146 265704
rect 3202 265648 3207 265704
rect -960 265646 3207 265648
rect -960 265556 480 265646
rect 3141 265643 3207 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3601 251290 3667 251293
rect -960 251288 3667 251290
rect -960 251232 3606 251288
rect 3662 251232 3667 251288
rect -960 251230 3667 251232
rect -960 251140 480 251230
rect 3601 251227 3667 251230
rect 583520 240396 584960 240636
rect 67357 240138 67423 240141
rect 67541 240138 67607 240141
rect 67357 240136 67607 240138
rect 67357 240080 67362 240136
rect 67418 240080 67546 240136
rect 67602 240080 67607 240136
rect 67357 240078 67607 240080
rect 67357 240075 67423 240078
rect 67541 240075 67607 240078
rect -960 237010 480 237100
rect 3233 237010 3299 237013
rect -960 237008 3299 237010
rect -960 236952 3238 237008
rect 3294 236952 3299 237008
rect -960 236950 3299 236952
rect -960 236860 480 236950
rect 3233 236947 3299 236950
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 3325 222594 3391 222597
rect -960 222592 3391 222594
rect -960 222536 3330 222592
rect 3386 222536 3391 222592
rect -960 222534 3391 222536
rect -960 222444 480 222534
rect 3325 222531 3391 222534
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 3509 208178 3575 208181
rect -960 208176 3575 208178
rect -960 208120 3514 208176
rect 3570 208120 3575 208176
rect -960 208118 3575 208120
rect -960 208028 480 208118
rect 3509 208115 3575 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect -960 193898 480 193988
rect 3509 193898 3575 193901
rect -960 193896 3575 193898
rect -960 193840 3514 193896
rect 3570 193840 3575 193896
rect -960 193838 3575 193840
rect -960 193748 480 193838
rect 3509 193835 3575 193838
rect 583520 193476 584960 193716
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 67398 177244 67404 177308
rect 67468 177306 67474 177308
rect 67541 177306 67607 177309
rect 67468 177304 67607 177306
rect 67468 177248 67546 177304
rect 67602 177248 67607 177304
rect 67468 177246 67607 177248
rect 67468 177244 67474 177246
rect 67541 177243 67607 177246
rect 60917 173906 60983 173909
rect 61101 173906 61167 173909
rect 60917 173904 61167 173906
rect 60917 173848 60922 173904
rect 60978 173848 61106 173904
rect 61162 173848 61167 173904
rect 60917 173846 61167 173848
rect 60917 173843 60983 173846
rect 61101 173843 61167 173846
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3417 165066 3483 165069
rect -960 165064 3483 165066
rect -960 165008 3422 165064
rect 3478 165008 3483 165064
rect -960 165006 3483 165008
rect -960 164916 480 165006
rect 3417 165003 3483 165006
rect 67398 164188 67404 164252
rect 67468 164250 67474 164252
rect 67541 164250 67607 164253
rect 67468 164248 67607 164250
rect 67468 164192 67546 164248
rect 67602 164192 67607 164248
rect 67468 164190 67607 164192
rect 67468 164188 67474 164190
rect 67541 164187 67607 164190
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect 60917 143578 60983 143581
rect 61193 143578 61259 143581
rect 60917 143576 61259 143578
rect 60917 143520 60922 143576
rect 60978 143520 61198 143576
rect 61254 143520 61259 143576
rect 60917 143518 61259 143520
rect 60917 143515 60983 143518
rect 61193 143515 61259 143518
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 67398 125972 67404 126036
rect 67468 126034 67474 126036
rect 67541 126034 67607 126037
rect 67468 126032 67607 126034
rect 67468 125976 67546 126032
rect 67602 125976 67607 126032
rect 67468 125974 67607 125976
rect 67468 125972 67474 125974
rect 67541 125971 67607 125974
rect 67398 125564 67404 125628
rect 67468 125626 67474 125628
rect 67541 125626 67607 125629
rect 67468 125624 67607 125626
rect 67468 125568 67546 125624
rect 67602 125568 67607 125624
rect 67468 125566 67607 125568
rect 67468 125564 67474 125566
rect 67541 125563 67607 125566
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 60733 106314 60799 106317
rect 61009 106314 61075 106317
rect 60733 106312 61075 106314
rect 60733 106256 60738 106312
rect 60794 106256 61014 106312
rect 61070 106256 61075 106312
rect 60733 106254 61075 106256
rect 60733 106251 60799 106254
rect 61009 106251 61075 106254
rect 583520 99636 584960 99876
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 125542 76468 125548 76532
rect 125612 76530 125618 76532
rect 135161 76530 135227 76533
rect 125612 76528 135227 76530
rect 125612 76472 135166 76528
rect 135222 76472 135227 76528
rect 125612 76470 135227 76472
rect 125612 76468 125618 76470
rect 135161 76467 135227 76470
rect 115790 76394 115796 76396
rect 108806 76334 115796 76394
rect 57462 76196 57468 76260
rect 57532 76258 57538 76260
rect 77201 76258 77267 76261
rect 57532 76198 60658 76258
rect 57532 76196 57538 76198
rect 60598 75986 60658 76198
rect 77201 76256 79978 76258
rect 77201 76200 77206 76256
rect 77262 76200 79978 76256
rect 77201 76198 79978 76200
rect 77201 76195 77267 76198
rect 67582 76122 67588 76124
rect 60782 76062 67588 76122
rect 60782 75986 60842 76062
rect 67582 76060 67588 76062
rect 67652 76060 67658 76124
rect 60598 75926 60842 75986
rect 79918 75986 79978 76198
rect 89529 76122 89595 76125
rect 80102 76120 89595 76122
rect 80102 76064 89534 76120
rect 89590 76064 89595 76120
rect 80102 76062 89595 76064
rect 80102 75986 80162 76062
rect 89529 76059 89595 76062
rect 89805 76122 89871 76125
rect 108806 76122 108866 76334
rect 115790 76332 115796 76334
rect 115860 76332 115866 76396
rect 140037 76394 140103 76397
rect 135302 76392 140103 76394
rect 135302 76336 140042 76392
rect 140098 76336 140103 76392
rect 135302 76334 140103 76336
rect 118877 76258 118943 76261
rect 125542 76258 125548 76260
rect 118877 76256 125548 76258
rect 118877 76200 118882 76256
rect 118938 76200 125548 76256
rect 118877 76198 125548 76200
rect 118877 76195 118943 76198
rect 125542 76196 125548 76198
rect 125612 76196 125618 76260
rect 89805 76120 96538 76122
rect 89805 76064 89810 76120
rect 89866 76064 96538 76120
rect 89805 76062 96538 76064
rect 89805 76059 89871 76062
rect 79918 75926 80162 75986
rect 96478 75986 96538 76062
rect 99422 76062 108866 76122
rect 135161 76122 135227 76125
rect 135302 76122 135362 76334
rect 140037 76331 140103 76334
rect 154481 76258 154547 76261
rect 583520 76258 584960 76348
rect 154481 76256 161490 76258
rect 154481 76200 154486 76256
rect 154542 76200 161490 76256
rect 154481 76198 161490 76200
rect 154481 76195 154547 76198
rect 147581 76122 147647 76125
rect 135161 76120 135362 76122
rect 135161 76064 135166 76120
rect 135222 76064 135362 76120
rect 135161 76062 135362 76064
rect 144870 76120 147647 76122
rect 144870 76064 147586 76120
rect 147642 76064 147647 76120
rect 144870 76062 147647 76064
rect 161430 76122 161490 76198
rect 171182 76198 180810 76258
rect 161430 76062 171058 76122
rect 99422 75986 99482 76062
rect 135161 76059 135227 76062
rect 96478 75926 99482 75986
rect 115790 75924 115796 75988
rect 115860 75986 115866 75988
rect 115933 75986 115999 75989
rect 115860 75984 115999 75986
rect 115860 75928 115938 75984
rect 115994 75928 115999 75984
rect 115860 75926 115999 75928
rect 115860 75924 115866 75926
rect 115933 75923 115999 75926
rect 140037 75986 140103 75989
rect 144870 75986 144930 76062
rect 147581 76059 147647 76062
rect 140037 75984 144930 75986
rect 140037 75928 140042 75984
rect 140098 75928 144930 75984
rect 140037 75926 144930 75928
rect 170998 75986 171058 76062
rect 171182 75986 171242 76198
rect 180750 76122 180810 76198
rect 190502 76198 200130 76258
rect 180750 76062 190378 76122
rect 170998 75926 171242 75986
rect 190318 75986 190378 76062
rect 190502 75986 190562 76198
rect 200070 76122 200130 76198
rect 209822 76198 219450 76258
rect 200070 76062 209698 76122
rect 190318 75926 190562 75986
rect 209638 75986 209698 76062
rect 209822 75986 209882 76198
rect 219390 76122 219450 76198
rect 229142 76198 238770 76258
rect 219390 76062 229018 76122
rect 209638 75926 209882 75986
rect 228958 75986 229018 76062
rect 229142 75986 229202 76198
rect 238710 76122 238770 76198
rect 248462 76198 258090 76258
rect 238710 76062 248338 76122
rect 228958 75926 229202 75986
rect 248278 75986 248338 76062
rect 248462 75986 248522 76198
rect 258030 76122 258090 76198
rect 267782 76198 277410 76258
rect 258030 76062 267658 76122
rect 248278 75926 248522 75986
rect 267598 75986 267658 76062
rect 267782 75986 267842 76198
rect 277350 76122 277410 76198
rect 287102 76198 296730 76258
rect 277350 76062 286978 76122
rect 267598 75926 267842 75986
rect 286918 75986 286978 76062
rect 287102 75986 287162 76198
rect 296670 76122 296730 76198
rect 306422 76198 316050 76258
rect 296670 76062 306298 76122
rect 286918 75926 287162 75986
rect 306238 75986 306298 76062
rect 306422 75986 306482 76198
rect 315990 76122 316050 76198
rect 325742 76198 335370 76258
rect 315990 76062 325618 76122
rect 306238 75926 306482 75986
rect 325558 75986 325618 76062
rect 325742 75986 325802 76198
rect 335310 76122 335370 76198
rect 345062 76198 354690 76258
rect 335310 76062 344938 76122
rect 325558 75926 325802 75986
rect 344878 75986 344938 76062
rect 345062 75986 345122 76198
rect 354630 76122 354690 76198
rect 364382 76198 374010 76258
rect 354630 76062 364258 76122
rect 344878 75926 345122 75986
rect 364198 75986 364258 76062
rect 364382 75986 364442 76198
rect 373950 76122 374010 76198
rect 383702 76198 393330 76258
rect 373950 76062 383578 76122
rect 364198 75926 364442 75986
rect 383518 75986 383578 76062
rect 383702 75986 383762 76198
rect 393270 76122 393330 76198
rect 403022 76198 412650 76258
rect 393270 76062 402898 76122
rect 383518 75926 383762 75986
rect 402838 75986 402898 76062
rect 403022 75986 403082 76198
rect 412590 76122 412650 76198
rect 422342 76198 431970 76258
rect 412590 76062 422218 76122
rect 402838 75926 403082 75986
rect 422158 75986 422218 76062
rect 422342 75986 422402 76198
rect 431910 76122 431970 76198
rect 441662 76198 451290 76258
rect 431910 76062 441538 76122
rect 422158 75926 422402 75986
rect 441478 75986 441538 76062
rect 441662 75986 441722 76198
rect 451230 76122 451290 76198
rect 460982 76198 470610 76258
rect 451230 76062 460858 76122
rect 441478 75926 441722 75986
rect 460798 75986 460858 76062
rect 460982 75986 461042 76198
rect 470550 76122 470610 76198
rect 480302 76198 489930 76258
rect 470550 76062 480178 76122
rect 460798 75926 461042 75986
rect 480118 75986 480178 76062
rect 480302 75986 480362 76198
rect 489870 76122 489930 76198
rect 499622 76198 509250 76258
rect 489870 76062 499498 76122
rect 480118 75926 480362 75986
rect 499438 75986 499498 76062
rect 499622 75986 499682 76198
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 499438 75926 499682 75986
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 140037 75923 140103 75926
rect 67582 75788 67588 75852
rect 67652 75850 67658 75852
rect 77201 75850 77267 75853
rect 67652 75848 77267 75850
rect 67652 75792 77206 75848
rect 77262 75792 77267 75848
rect 67652 75790 77267 75792
rect 67652 75788 67658 75790
rect 77201 75787 77267 75790
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 125542 40564 125548 40628
rect 125612 40626 125618 40628
rect 135161 40626 135227 40629
rect 125612 40624 135227 40626
rect 125612 40568 135166 40624
rect 135222 40568 135227 40624
rect 125612 40566 135227 40568
rect 125612 40564 125618 40566
rect 135161 40563 135227 40566
rect 115790 40490 115796 40492
rect 108806 40430 115796 40490
rect 57646 40292 57652 40356
rect 57716 40354 57722 40356
rect 77201 40354 77267 40357
rect 57716 40294 60658 40354
rect 57716 40292 57722 40294
rect 60598 40082 60658 40294
rect 77201 40352 79978 40354
rect 77201 40296 77206 40352
rect 77262 40296 79978 40352
rect 77201 40294 79978 40296
rect 77201 40291 77267 40294
rect 67582 40218 67588 40220
rect 60782 40158 67588 40218
rect 60782 40082 60842 40158
rect 67582 40156 67588 40158
rect 67652 40156 67658 40220
rect 60598 40022 60842 40082
rect 79918 40082 79978 40294
rect 89529 40218 89595 40221
rect 80102 40216 89595 40218
rect 80102 40160 89534 40216
rect 89590 40160 89595 40216
rect 80102 40158 89595 40160
rect 80102 40082 80162 40158
rect 89529 40155 89595 40158
rect 91737 40218 91803 40221
rect 108806 40218 108866 40430
rect 115790 40428 115796 40430
rect 115860 40428 115866 40492
rect 140037 40490 140103 40493
rect 135302 40488 140103 40490
rect 135302 40432 140042 40488
rect 140098 40432 140103 40488
rect 135302 40430 140103 40432
rect 118877 40354 118943 40357
rect 125542 40354 125548 40356
rect 118877 40352 125548 40354
rect 118877 40296 118882 40352
rect 118938 40296 125548 40352
rect 118877 40294 125548 40296
rect 118877 40291 118943 40294
rect 125542 40292 125548 40294
rect 125612 40292 125618 40356
rect 91737 40216 96538 40218
rect 91737 40160 91742 40216
rect 91798 40160 96538 40216
rect 91737 40158 96538 40160
rect 91737 40155 91803 40158
rect 79918 40022 80162 40082
rect 96478 40082 96538 40158
rect 99422 40158 108866 40218
rect 135161 40218 135227 40221
rect 135302 40218 135362 40430
rect 140037 40427 140103 40430
rect 154481 40354 154547 40357
rect 154481 40352 161490 40354
rect 154481 40296 154486 40352
rect 154542 40296 161490 40352
rect 154481 40294 161490 40296
rect 154481 40291 154547 40294
rect 147581 40218 147647 40221
rect 135161 40216 135362 40218
rect 135161 40160 135166 40216
rect 135222 40160 135362 40216
rect 135161 40158 135362 40160
rect 144870 40216 147647 40218
rect 144870 40160 147586 40216
rect 147642 40160 147647 40216
rect 144870 40158 147647 40160
rect 161430 40218 161490 40294
rect 171182 40294 180810 40354
rect 161430 40158 171058 40218
rect 99422 40082 99482 40158
rect 135161 40155 135227 40158
rect 96478 40022 99482 40082
rect 115790 40020 115796 40084
rect 115860 40082 115866 40084
rect 115933 40082 115999 40085
rect 115860 40080 115999 40082
rect 115860 40024 115938 40080
rect 115994 40024 115999 40080
rect 115860 40022 115999 40024
rect 115860 40020 115866 40022
rect 115933 40019 115999 40022
rect 140037 40082 140103 40085
rect 144870 40082 144930 40158
rect 147581 40155 147647 40158
rect 140037 40080 144930 40082
rect 140037 40024 140042 40080
rect 140098 40024 144930 40080
rect 140037 40022 144930 40024
rect 170998 40082 171058 40158
rect 171182 40082 171242 40294
rect 180750 40218 180810 40294
rect 190502 40294 200130 40354
rect 180750 40158 190378 40218
rect 170998 40022 171242 40082
rect 190318 40082 190378 40158
rect 190502 40082 190562 40294
rect 200070 40218 200130 40294
rect 209822 40294 219450 40354
rect 200070 40158 209698 40218
rect 190318 40022 190562 40082
rect 209638 40082 209698 40158
rect 209822 40082 209882 40294
rect 219390 40218 219450 40294
rect 229142 40294 238770 40354
rect 219390 40158 229018 40218
rect 209638 40022 209882 40082
rect 228958 40082 229018 40158
rect 229142 40082 229202 40294
rect 238710 40218 238770 40294
rect 248462 40294 258090 40354
rect 238710 40158 248338 40218
rect 228958 40022 229202 40082
rect 248278 40082 248338 40158
rect 248462 40082 248522 40294
rect 258030 40218 258090 40294
rect 267782 40294 277410 40354
rect 258030 40158 267658 40218
rect 248278 40022 248522 40082
rect 267598 40082 267658 40158
rect 267782 40082 267842 40294
rect 277350 40218 277410 40294
rect 287102 40294 296730 40354
rect 277350 40158 286978 40218
rect 267598 40022 267842 40082
rect 286918 40082 286978 40158
rect 287102 40082 287162 40294
rect 296670 40218 296730 40294
rect 306422 40294 316050 40354
rect 296670 40158 306298 40218
rect 286918 40022 287162 40082
rect 306238 40082 306298 40158
rect 306422 40082 306482 40294
rect 315990 40218 316050 40294
rect 325742 40294 335370 40354
rect 315990 40158 325618 40218
rect 306238 40022 306482 40082
rect 325558 40082 325618 40158
rect 325742 40082 325802 40294
rect 335310 40218 335370 40294
rect 345062 40294 354690 40354
rect 335310 40158 344938 40218
rect 325558 40022 325802 40082
rect 344878 40082 344938 40158
rect 345062 40082 345122 40294
rect 354630 40218 354690 40294
rect 364382 40294 374010 40354
rect 354630 40158 364258 40218
rect 344878 40022 345122 40082
rect 364198 40082 364258 40158
rect 364382 40082 364442 40294
rect 373950 40218 374010 40294
rect 383702 40294 393330 40354
rect 373950 40158 383578 40218
rect 364198 40022 364442 40082
rect 383518 40082 383578 40158
rect 383702 40082 383762 40294
rect 393270 40218 393330 40294
rect 403022 40294 412650 40354
rect 393270 40158 402898 40218
rect 383518 40022 383762 40082
rect 402838 40082 402898 40158
rect 403022 40082 403082 40294
rect 412590 40218 412650 40294
rect 422342 40294 431970 40354
rect 412590 40158 422218 40218
rect 402838 40022 403082 40082
rect 422158 40082 422218 40158
rect 422342 40082 422402 40294
rect 431910 40218 431970 40294
rect 441662 40294 451290 40354
rect 431910 40158 441538 40218
rect 422158 40022 422402 40082
rect 441478 40082 441538 40158
rect 441662 40082 441722 40294
rect 451230 40218 451290 40294
rect 460982 40294 470610 40354
rect 451230 40158 460858 40218
rect 441478 40022 441722 40082
rect 460798 40082 460858 40158
rect 460982 40082 461042 40294
rect 470550 40218 470610 40294
rect 480302 40294 489930 40354
rect 470550 40158 480178 40218
rect 460798 40022 461042 40082
rect 480118 40082 480178 40158
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 140037 40019 140103 40022
rect 67582 39884 67588 39948
rect 67652 39946 67658 39948
rect 77201 39946 77267 39949
rect 67652 39944 77267 39946
rect 67652 39888 77206 39944
rect 77262 39888 77267 39944
rect 67652 39886 77267 39888
rect 67652 39884 67658 39886
rect 77201 39883 77267 39886
rect 67449 37226 67515 37229
rect 67725 37226 67791 37229
rect 67449 37224 67791 37226
rect 67449 37168 67454 37224
rect 67510 37168 67730 37224
rect 67786 37168 67791 37224
rect 67449 37166 67791 37168
rect 67449 37163 67515 37166
rect 67725 37163 67791 37166
rect -960 35866 480 35956
rect 2773 35866 2839 35869
rect -960 35864 2839 35866
rect -960 35808 2778 35864
rect 2834 35808 2839 35864
rect -960 35806 2839 35808
rect -960 35716 480 35806
rect 2773 35803 2839 35806
rect 86902 29548 86908 29612
rect 86972 29610 86978 29612
rect 91737 29610 91803 29613
rect 86972 29608 91803 29610
rect 86972 29552 91742 29608
rect 91798 29552 91803 29608
rect 86972 29550 91803 29552
rect 86972 29548 86978 29550
rect 91737 29547 91803 29550
rect 115790 29474 115796 29476
rect 108806 29414 115796 29474
rect 57830 29276 57836 29340
rect 57900 29338 57906 29340
rect 57900 29278 79794 29338
rect 57900 29276 57906 29278
rect 79734 29202 79794 29278
rect 86902 29202 86908 29204
rect 79734 29142 86908 29202
rect 86902 29140 86908 29142
rect 86972 29140 86978 29204
rect 91737 29202 91803 29205
rect 108806 29202 108866 29414
rect 115790 29412 115796 29414
rect 115860 29412 115866 29476
rect 133822 29412 133828 29476
rect 133892 29474 133898 29476
rect 143441 29474 143507 29477
rect 133892 29472 143507 29474
rect 133892 29416 143446 29472
rect 143502 29416 143507 29472
rect 133892 29414 143507 29416
rect 133892 29412 133898 29414
rect 143441 29411 143507 29414
rect 120809 29338 120875 29341
rect 128261 29338 128327 29341
rect 120809 29336 128327 29338
rect 120809 29280 120814 29336
rect 120870 29280 128266 29336
rect 128322 29280 128327 29336
rect 120809 29278 128327 29280
rect 120809 29275 120875 29278
rect 128261 29275 128327 29278
rect 154481 29338 154547 29341
rect 583520 29338 584960 29428
rect 154481 29336 161490 29338
rect 154481 29280 154486 29336
rect 154542 29280 161490 29336
rect 154481 29278 161490 29280
rect 154481 29275 154547 29278
rect 91737 29200 96538 29202
rect 91737 29144 91742 29200
rect 91798 29144 96538 29200
rect 91737 29142 96538 29144
rect 91737 29139 91803 29142
rect 96478 29066 96538 29142
rect 99422 29142 108866 29202
rect 128445 29202 128511 29205
rect 133822 29202 133828 29204
rect 128445 29200 133828 29202
rect 128445 29144 128450 29200
rect 128506 29144 133828 29200
rect 128445 29142 133828 29144
rect 99422 29066 99482 29142
rect 128445 29139 128511 29142
rect 133822 29140 133828 29142
rect 133892 29140 133898 29204
rect 147581 29202 147647 29205
rect 144870 29200 147647 29202
rect 144870 29144 147586 29200
rect 147642 29144 147647 29200
rect 144870 29142 147647 29144
rect 161430 29202 161490 29278
rect 171182 29278 180810 29338
rect 161430 29142 171058 29202
rect 96478 29006 99482 29066
rect 115790 29004 115796 29068
rect 115860 29066 115866 29068
rect 115933 29066 115999 29069
rect 115860 29064 115999 29066
rect 115860 29008 115938 29064
rect 115994 29008 115999 29064
rect 115860 29006 115999 29008
rect 115860 29004 115866 29006
rect 115933 29003 115999 29006
rect 143441 29066 143507 29069
rect 144870 29066 144930 29142
rect 147581 29139 147647 29142
rect 143441 29064 144930 29066
rect 143441 29008 143446 29064
rect 143502 29008 144930 29064
rect 143441 29006 144930 29008
rect 170998 29066 171058 29142
rect 171182 29066 171242 29278
rect 180750 29202 180810 29278
rect 190502 29278 200130 29338
rect 180750 29142 190378 29202
rect 170998 29006 171242 29066
rect 190318 29066 190378 29142
rect 190502 29066 190562 29278
rect 200070 29202 200130 29278
rect 209822 29278 219450 29338
rect 200070 29142 209698 29202
rect 190318 29006 190562 29066
rect 209638 29066 209698 29142
rect 209822 29066 209882 29278
rect 219390 29202 219450 29278
rect 229142 29278 238770 29338
rect 219390 29142 229018 29202
rect 209638 29006 209882 29066
rect 228958 29066 229018 29142
rect 229142 29066 229202 29278
rect 238710 29202 238770 29278
rect 248462 29278 258090 29338
rect 238710 29142 248338 29202
rect 228958 29006 229202 29066
rect 248278 29066 248338 29142
rect 248462 29066 248522 29278
rect 258030 29202 258090 29278
rect 267782 29278 277410 29338
rect 258030 29142 267658 29202
rect 248278 29006 248522 29066
rect 267598 29066 267658 29142
rect 267782 29066 267842 29278
rect 277350 29202 277410 29278
rect 287102 29278 296730 29338
rect 277350 29142 286978 29202
rect 267598 29006 267842 29066
rect 286918 29066 286978 29142
rect 287102 29066 287162 29278
rect 296670 29202 296730 29278
rect 306422 29278 316050 29338
rect 296670 29142 306298 29202
rect 286918 29006 287162 29066
rect 306238 29066 306298 29142
rect 306422 29066 306482 29278
rect 315990 29202 316050 29278
rect 325742 29278 335370 29338
rect 315990 29142 325618 29202
rect 306238 29006 306482 29066
rect 325558 29066 325618 29142
rect 325742 29066 325802 29278
rect 335310 29202 335370 29278
rect 345062 29278 354690 29338
rect 335310 29142 344938 29202
rect 325558 29006 325802 29066
rect 344878 29066 344938 29142
rect 345062 29066 345122 29278
rect 354630 29202 354690 29278
rect 364382 29278 374010 29338
rect 354630 29142 364258 29202
rect 344878 29006 345122 29066
rect 364198 29066 364258 29142
rect 364382 29066 364442 29278
rect 373950 29202 374010 29278
rect 383702 29278 393330 29338
rect 373950 29142 383578 29202
rect 364198 29006 364442 29066
rect 383518 29066 383578 29142
rect 383702 29066 383762 29278
rect 393270 29202 393330 29278
rect 403022 29278 412650 29338
rect 393270 29142 402898 29202
rect 383518 29006 383762 29066
rect 402838 29066 402898 29142
rect 403022 29066 403082 29278
rect 412590 29202 412650 29278
rect 422342 29278 431970 29338
rect 412590 29142 422218 29202
rect 402838 29006 403082 29066
rect 422158 29066 422218 29142
rect 422342 29066 422402 29278
rect 431910 29202 431970 29278
rect 441662 29278 451290 29338
rect 431910 29142 441538 29202
rect 422158 29006 422402 29066
rect 441478 29066 441538 29142
rect 441662 29066 441722 29278
rect 451230 29202 451290 29278
rect 460982 29278 470610 29338
rect 451230 29142 460858 29202
rect 441478 29006 441722 29066
rect 460798 29066 460858 29142
rect 460982 29066 461042 29278
rect 470550 29202 470610 29278
rect 480302 29278 489930 29338
rect 470550 29142 480178 29202
rect 460798 29006 461042 29066
rect 480118 29066 480178 29142
rect 480302 29066 480362 29278
rect 489870 29202 489930 29278
rect 499622 29278 509250 29338
rect 489870 29142 499498 29202
rect 480118 29006 480362 29066
rect 499438 29066 499498 29142
rect 499622 29066 499682 29278
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 499438 29006 499682 29066
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 143441 29003 143507 29006
rect -960 21450 480 21540
rect 2865 21450 2931 21453
rect -960 21448 2931 21450
rect -960 21392 2870 21448
rect 2926 21392 2931 21448
rect -960 21390 2931 21392
rect -960 21300 480 21390
rect 2865 21387 2931 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 90909 5266 90975 5269
rect 208393 5266 208459 5269
rect 90909 5264 208459 5266
rect 90909 5208 90914 5264
rect 90970 5208 208398 5264
rect 208454 5208 208459 5264
rect 90909 5206 208459 5208
rect 90909 5203 90975 5206
rect 208393 5203 208459 5206
rect 94497 5130 94563 5133
rect 213913 5130 213979 5133
rect 94497 5128 213979 5130
rect 94497 5072 94502 5128
rect 94558 5072 213918 5128
rect 213974 5072 213979 5128
rect 94497 5070 213979 5072
rect 94497 5067 94563 5070
rect 213913 5067 213979 5070
rect 101581 4994 101647 4997
rect 226333 4994 226399 4997
rect 101581 4992 226399 4994
rect 101581 4936 101586 4992
rect 101642 4936 226338 4992
rect 226394 4936 226399 4992
rect 101581 4934 226399 4936
rect 101581 4931 101647 4934
rect 226333 4931 226399 4934
rect 131389 4858 131455 4861
rect 274633 4858 274699 4861
rect 131389 4856 274699 4858
rect 131389 4800 131394 4856
rect 131450 4800 274638 4856
rect 274694 4800 274699 4856
rect 131389 4798 274699 4800
rect 131389 4795 131455 4798
rect 274633 4795 274699 4798
rect 78949 4042 79015 4045
rect 82997 4042 83063 4045
rect 78949 4040 83063 4042
rect 78949 3984 78954 4040
rect 79010 3984 83002 4040
rect 83058 3984 83063 4040
rect 78949 3982 83063 3984
rect 78949 3979 79015 3982
rect 82997 3979 83063 3982
rect 86033 4042 86099 4045
rect 89713 4042 89779 4045
rect 86033 4040 89779 4042
rect 86033 3984 86038 4040
rect 86094 3984 89718 4040
rect 89774 3984 89779 4040
rect 86033 3982 89779 3984
rect 86033 3979 86099 3982
rect 89713 3979 89779 3982
rect 93209 3906 93275 3909
rect 93853 3906 93919 3909
rect 93209 3904 93919 3906
rect 93209 3848 93214 3904
rect 93270 3848 93858 3904
rect 93914 3848 93919 3904
rect 93209 3846 93919 3848
rect 93209 3843 93275 3846
rect 93853 3843 93919 3846
rect 95509 3906 95575 3909
rect 96613 3906 96679 3909
rect 95509 3904 96679 3906
rect 95509 3848 95514 3904
rect 95570 3848 96618 3904
rect 96674 3848 96679 3904
rect 95509 3846 96679 3848
rect 95509 3843 95575 3846
rect 96613 3843 96679 3846
rect 102685 3906 102751 3909
rect 104893 3906 104959 3909
rect 102685 3904 104959 3906
rect 102685 3848 102690 3904
rect 102746 3848 104898 3904
rect 104954 3848 104959 3904
rect 102685 3846 104959 3848
rect 102685 3843 102751 3846
rect 104893 3843 104959 3846
rect 109861 3906 109927 3909
rect 117313 3906 117379 3909
rect 109861 3904 117379 3906
rect 109861 3848 109866 3904
rect 109922 3848 117318 3904
rect 117374 3848 117379 3904
rect 109861 3846 117379 3848
rect 109861 3843 109927 3846
rect 117313 3843 117379 3846
rect 84929 3770 84995 3773
rect 198733 3770 198799 3773
rect 84929 3768 198799 3770
rect 84929 3712 84934 3768
rect 84990 3712 198738 3768
rect 198794 3712 198799 3768
rect 84929 3710 198799 3712
rect 84929 3707 84995 3710
rect 198733 3707 198799 3710
rect 74625 3634 74691 3637
rect 84009 3634 84075 3637
rect 74625 3632 84075 3634
rect 74625 3576 74630 3632
rect 74686 3576 84014 3632
rect 84070 3576 84075 3632
rect 74625 3574 84075 3576
rect 74625 3571 74691 3574
rect 84009 3571 84075 3574
rect 92105 3634 92171 3637
rect 209773 3634 209839 3637
rect 92105 3632 209839 3634
rect 92105 3576 92110 3632
rect 92166 3576 209778 3632
rect 209834 3576 209839 3632
rect 92105 3574 209839 3576
rect 92105 3571 92171 3574
rect 209773 3571 209839 3574
rect 68645 3498 68711 3501
rect 84101 3498 84167 3501
rect 68645 3496 84167 3498
rect 68645 3440 68650 3496
rect 68706 3440 84106 3496
rect 84162 3440 84167 3496
rect 68645 3438 84167 3440
rect 68645 3435 68711 3438
rect 84101 3435 84167 3438
rect 99281 3498 99347 3501
rect 222193 3498 222259 3501
rect 99281 3496 222259 3498
rect 99281 3440 99286 3496
rect 99342 3440 222198 3496
rect 222254 3440 222259 3496
rect 99281 3438 222259 3440
rect 99281 3435 99347 3438
rect 222193 3435 222259 3438
rect 93853 3362 93919 3365
rect 99373 3362 99439 3365
rect 93853 3360 99439 3362
rect 93853 3304 93858 3360
rect 93914 3304 99378 3360
rect 99434 3304 99439 3360
rect 93853 3302 99439 3304
rect 93853 3299 93919 3302
rect 99373 3299 99439 3302
rect 103973 3362 104039 3365
rect 229093 3362 229159 3365
rect 103973 3360 229159 3362
rect 103973 3304 103978 3360
rect 104034 3304 229098 3360
rect 229154 3304 229159 3360
rect 103973 3302 229159 3304
rect 103973 3299 104039 3302
rect 229093 3299 229159 3302
rect 93945 3226 94011 3229
rect 99465 3226 99531 3229
rect 93945 3224 99531 3226
rect 93945 3168 93950 3224
rect 94006 3168 99470 3224
rect 99526 3168 99531 3224
rect 93945 3166 99531 3168
rect 93945 3163 94011 3166
rect 99465 3163 99531 3166
<< via3 >>
rect 550588 697308 550652 697372
rect 59124 697172 59188 697236
rect 550588 696900 550652 696964
rect 183508 686428 183572 686492
rect 376708 686428 376772 686492
rect 434668 686428 434732 686492
rect 164188 686292 164252 686356
rect 357388 686292 357452 686356
rect 550588 686292 550652 686356
rect 57836 686156 57900 686220
rect 183508 686156 183572 686220
rect 164188 685884 164252 685948
rect 299428 686156 299492 686220
rect 299428 685884 299492 685948
rect 376708 686156 376772 686220
rect 357388 685884 357452 685948
rect 434668 686020 434732 686084
rect 550588 685884 550652 685948
rect 183508 674052 183572 674116
rect 376708 674052 376772 674116
rect 357388 673916 357452 673980
rect 58204 673780 58268 673844
rect 183508 673780 183572 673844
rect 299428 673780 299492 673844
rect 299428 673508 299492 673572
rect 376708 673780 376772 673844
rect 357388 673508 357452 673572
rect 129228 652896 129292 652900
rect 129228 652840 129278 652896
rect 129278 652840 129292 652896
rect 129228 652836 129292 652840
rect 133644 652896 133708 652900
rect 133644 652840 133658 652896
rect 133658 652840 133708 652896
rect 133644 652836 133708 652840
rect 259132 652896 259196 652900
rect 259132 652840 259182 652896
rect 259182 652840 259196 652896
rect 259132 652836 259196 652840
rect 263732 652896 263796 652900
rect 263732 652840 263782 652896
rect 263782 652840 263796 652896
rect 263732 652836 263796 652840
rect 378548 652896 378612 652900
rect 378548 652840 378562 652896
rect 378562 652840 378612 652896
rect 378548 652836 378612 652840
rect 383516 652896 383580 652900
rect 383516 652840 383530 652896
rect 383530 652840 383580 652896
rect 383516 652836 383580 652840
rect 507900 652896 507964 652900
rect 507900 652840 507914 652896
rect 507914 652840 507964 652896
rect 507900 652836 507964 652840
rect 513420 652896 513484 652900
rect 513420 652840 513434 652896
rect 513434 652840 513484 652896
rect 513420 652836 513484 652840
rect 211108 560008 211172 560012
rect 211108 559952 211122 560008
rect 211122 559952 211172 560008
rect 211108 559948 211172 559952
rect 210556 559812 210620 559876
rect 351868 559268 351932 559332
rect 358860 559268 358924 559332
rect 67404 558860 67468 558924
rect 69796 558860 69860 558924
rect 72372 558920 72436 558924
rect 72372 558864 72422 558920
rect 72422 558864 72436 558920
rect 72372 558860 72436 558864
rect 73660 558920 73724 558924
rect 73660 558864 73710 558920
rect 73710 558864 73724 558920
rect 73660 558860 73724 558864
rect 74948 558860 75012 558924
rect 75868 558860 75932 558924
rect 77340 558920 77404 558924
rect 77340 558864 77390 558920
rect 77390 558864 77404 558920
rect 77340 558860 77404 558864
rect 78444 558920 78508 558924
rect 78444 558864 78494 558920
rect 78494 558864 78508 558920
rect 78444 558860 78508 558864
rect 79364 558860 79428 558924
rect 80652 558920 80716 558924
rect 80652 558864 80702 558920
rect 80702 558864 80716 558920
rect 80652 558860 80716 558864
rect 82124 558860 82188 558924
rect 82860 558920 82924 558924
rect 82860 558864 82910 558920
rect 82910 558864 82924 558920
rect 82860 558860 82924 558864
rect 84700 558860 84764 558924
rect 85436 558920 85500 558924
rect 85436 558864 85450 558920
rect 85450 558864 85500 558920
rect 85436 558860 85500 558864
rect 85620 558920 85684 558924
rect 85620 558864 85670 558920
rect 85670 558864 85684 558920
rect 85620 558860 85684 558864
rect 86724 558860 86788 558924
rect 88196 558860 88260 558924
rect 88932 558920 88996 558924
rect 88932 558864 88982 558920
rect 88982 558864 88996 558920
rect 88932 558860 88996 558864
rect 89116 558860 89180 558924
rect 90036 558920 90100 558924
rect 90036 558864 90086 558920
rect 90086 558864 90100 558920
rect 90036 558860 90100 558864
rect 91324 558920 91388 558924
rect 91324 558864 91374 558920
rect 91374 558864 91388 558920
rect 91324 558860 91388 558864
rect 92428 558920 92492 558924
rect 92428 558864 92478 558920
rect 92478 558864 92492 558920
rect 92428 558860 92492 558864
rect 93532 558920 93596 558924
rect 93532 558864 93582 558920
rect 93582 558864 93596 558920
rect 93532 558860 93596 558864
rect 94636 558920 94700 558924
rect 94636 558864 94650 558920
rect 94650 558864 94700 558920
rect 94636 558860 94700 558864
rect 95372 558920 95436 558924
rect 95372 558864 95386 558920
rect 95386 558864 95436 558920
rect 95372 558860 95436 558864
rect 96660 558920 96724 558924
rect 96660 558864 96674 558920
rect 96674 558864 96724 558920
rect 96660 558860 96724 558864
rect 98316 558920 98380 558924
rect 98316 558864 98330 558920
rect 98330 558864 98380 558920
rect 98316 558860 98380 558864
rect 99604 558920 99668 558924
rect 99604 558864 99618 558920
rect 99618 558864 99668 558920
rect 99604 558860 99668 558864
rect 100156 558860 100220 558924
rect 101996 558920 102060 558924
rect 101996 558864 102010 558920
rect 102010 558864 102060 558920
rect 101996 558860 102060 558864
rect 102732 558920 102796 558924
rect 102732 558864 102746 558920
rect 102746 558864 102796 558920
rect 102732 558860 102796 558864
rect 103284 558860 103348 558924
rect 104020 558920 104084 558924
rect 104020 558864 104034 558920
rect 104034 558864 104084 558920
rect 104020 558860 104084 558864
rect 104756 558920 104820 558924
rect 104756 558864 104806 558920
rect 104806 558864 104820 558920
rect 104756 558860 104820 558864
rect 105308 558920 105372 558924
rect 105308 558864 105358 558920
rect 105358 558864 105372 558920
rect 105308 558860 105372 558864
rect 106044 558860 106108 558924
rect 107148 558860 107212 558924
rect 107700 558860 107764 558924
rect 108436 558860 108500 558924
rect 109540 558860 109604 558924
rect 193812 558920 193876 558924
rect 193812 558864 193826 558920
rect 193826 558864 193876 558920
rect 193812 558860 193876 558864
rect 202644 558860 202708 558924
rect 203932 558860 203996 558924
rect 205404 558860 205468 558924
rect 211844 558920 211908 558924
rect 211844 558864 211894 558920
rect 211894 558864 211908 558920
rect 211844 558860 211908 558864
rect 213132 558920 213196 558924
rect 213132 558864 213182 558920
rect 213182 558864 213196 558920
rect 213132 558860 213196 558864
rect 214052 558860 214116 558924
rect 216260 558860 216324 558924
rect 217548 558920 217612 558924
rect 217548 558864 217598 558920
rect 217598 558864 217612 558920
rect 217548 558860 217612 558864
rect 217916 558920 217980 558924
rect 217916 558864 217930 558920
rect 217930 558864 217980 558920
rect 217916 558860 217980 558864
rect 218836 558920 218900 558924
rect 218836 558864 218886 558920
rect 218886 558864 218900 558920
rect 218836 558860 218900 558864
rect 219204 558860 219268 558924
rect 220124 558920 220188 558924
rect 220124 558864 220138 558920
rect 220138 558864 220188 558920
rect 220124 558860 220188 558864
rect 220676 558920 220740 558924
rect 220676 558864 220726 558920
rect 220726 558864 220740 558920
rect 220676 558860 220740 558864
rect 221044 558920 221108 558924
rect 221044 558864 221094 558920
rect 221094 558864 221108 558920
rect 221044 558860 221108 558864
rect 221964 558860 222028 558924
rect 222332 558920 222396 558924
rect 222332 558864 222346 558920
rect 222346 558864 222396 558920
rect 222332 558860 222396 558864
rect 223252 558860 223316 558924
rect 224356 558860 224420 558924
rect 225828 558920 225892 558924
rect 225828 558864 225842 558920
rect 225842 558864 225892 558920
rect 225828 558860 225892 558864
rect 226196 558920 226260 558924
rect 226196 558864 226246 558920
rect 226246 558864 226260 558920
rect 226196 558860 226260 558864
rect 227116 558920 227180 558924
rect 227116 558864 227166 558920
rect 227166 558864 227180 558920
rect 227116 558860 227180 558864
rect 227484 558860 227548 558924
rect 228772 558860 228836 558924
rect 229508 558920 229572 558924
rect 229508 558864 229522 558920
rect 229522 558864 229572 558920
rect 229508 558860 229572 558864
rect 230244 558860 230308 558924
rect 230796 558860 230860 558924
rect 232820 558860 232884 558924
rect 233004 558860 233068 558924
rect 234476 558920 234540 558924
rect 234476 558864 234526 558920
rect 234526 558864 234540 558920
rect 234476 558860 234540 558864
rect 235764 558860 235828 558924
rect 237236 558920 237300 558924
rect 237236 558864 237286 558920
rect 237286 558864 237300 558920
rect 237236 558860 237300 558864
rect 239628 558860 239692 558924
rect 313780 558920 313844 558924
rect 313780 558864 313794 558920
rect 313794 558864 313844 558920
rect 313780 558860 313844 558864
rect 316172 558860 316236 558924
rect 318932 558860 318996 558924
rect 320956 558860 321020 558924
rect 322796 558860 322860 558924
rect 325188 558860 325252 558924
rect 326292 558860 326356 558924
rect 327580 558860 327644 558924
rect 331076 558860 331140 558924
rect 331812 558920 331876 558924
rect 331812 558864 331826 558920
rect 331826 558864 331876 558920
rect 331812 558860 331876 558864
rect 333284 558860 333348 558924
rect 334572 558860 334636 558924
rect 335860 558860 335924 558924
rect 336780 558920 336844 558924
rect 336780 558864 336794 558920
rect 336794 558864 336844 558920
rect 336780 558860 336844 558864
rect 337700 558860 337764 558924
rect 339172 558860 339236 558924
rect 340460 558860 340524 558924
rect 341748 558860 341812 558924
rect 342668 558860 342732 558924
rect 343956 558860 344020 558924
rect 344324 558920 344388 558924
rect 344324 558864 344338 558920
rect 344338 558864 344388 558920
rect 344324 558860 344388 558864
rect 346164 558860 346228 558924
rect 347452 558860 347516 558924
rect 348740 558860 348804 558924
rect 349660 558860 349724 558924
rect 352420 558860 352484 558924
rect 443132 558920 443196 558924
rect 443132 558864 443146 558920
rect 443146 558864 443196 558920
rect 443132 558860 443196 558864
rect 446260 558860 446324 558924
rect 447364 558860 447428 558924
rect 448468 558860 448532 558924
rect 449940 558860 450004 558924
rect 452884 558860 452948 558924
rect 453620 558860 453684 558924
rect 454724 558920 454788 558924
rect 454724 558864 454738 558920
rect 454738 558864 454788 558920
rect 454724 558860 454788 558864
rect 458404 558860 458468 558924
rect 460980 558920 461044 558924
rect 460980 558864 460994 558920
rect 460994 558864 461044 558920
rect 460980 558860 461044 558864
rect 461716 558920 461780 558924
rect 461716 558864 461766 558920
rect 461766 558864 461780 558920
rect 461716 558860 461780 558864
rect 463372 558860 463436 558924
rect 464476 558860 464540 558924
rect 465764 558860 465828 558924
rect 466868 558860 466932 558924
rect 467972 558860 468036 558924
rect 468708 558860 468772 558924
rect 470364 558860 470428 558924
rect 471468 558860 471532 558924
rect 472756 558860 472820 558924
rect 474044 558860 474108 558924
rect 474964 558860 475028 558924
rect 476252 558920 476316 558924
rect 476252 558864 476266 558920
rect 476266 558864 476316 558920
rect 476252 558860 476316 558864
rect 477172 558920 477236 558924
rect 477172 558864 477186 558920
rect 477186 558864 477236 558920
rect 477172 558860 477236 558864
rect 478276 558920 478340 558924
rect 478276 558864 478326 558920
rect 478326 558864 478340 558920
rect 478276 558860 478340 558864
rect 479380 558920 479444 558924
rect 479380 558864 479430 558920
rect 479430 558864 479444 558920
rect 479380 558860 479444 558864
rect 480852 558860 480916 558924
rect 483428 558860 483492 558924
rect 485636 558860 485700 558924
rect 486004 558860 486068 558924
rect 61700 558724 61764 558788
rect 63540 558724 63604 558788
rect 70164 558784 70228 558788
rect 70164 558728 70214 558784
rect 70214 558728 70228 558784
rect 70164 558724 70228 558728
rect 81020 558724 81084 558788
rect 81756 558724 81820 558788
rect 84148 558724 84212 558788
rect 86356 558724 86420 558788
rect 87828 558784 87892 558788
rect 87828 558728 87878 558784
rect 87878 558728 87892 558784
rect 87828 558724 87892 558728
rect 100340 558784 100404 558788
rect 100340 558728 100354 558784
rect 100354 558728 100404 558784
rect 100340 558724 100404 558728
rect 101444 558724 101508 558788
rect 106228 558784 106292 558788
rect 106228 558728 106278 558784
rect 106278 558728 106292 558784
rect 106228 558724 106292 558728
rect 108620 558784 108684 558788
rect 108620 558728 108634 558784
rect 108634 558728 108684 558784
rect 108620 558724 108684 558728
rect 196204 558724 196268 558788
rect 201724 558724 201788 558788
rect 202460 558724 202524 558788
rect 204852 558784 204916 558788
rect 204852 558728 204902 558784
rect 204902 558728 204916 558784
rect 204852 558724 204916 558728
rect 215340 558784 215404 558788
rect 215340 558728 215354 558784
rect 215354 558728 215404 558784
rect 215340 558724 215404 558728
rect 216628 558724 216692 558788
rect 217364 558724 217428 558788
rect 223620 558784 223684 558788
rect 223620 558728 223634 558784
rect 223634 558728 223684 558784
rect 223620 558724 223684 558728
rect 224540 558724 224604 558788
rect 225644 558724 225708 558788
rect 227852 558724 227916 558788
rect 232636 558724 232700 558788
rect 233556 558724 233620 558788
rect 236132 558724 236196 558788
rect 322428 558724 322492 558788
rect 327028 558724 327092 558788
rect 328500 558724 328564 558788
rect 332732 558784 332796 558788
rect 332732 558728 332746 558784
rect 332746 558728 332796 558784
rect 332732 558724 332796 558728
rect 334020 558784 334084 558788
rect 334020 558728 334070 558784
rect 334070 558728 334084 558784
rect 334020 558724 334084 558728
rect 335492 558784 335556 558788
rect 335492 558728 335506 558784
rect 335506 558728 335556 558784
rect 335492 558724 335556 558728
rect 336596 558784 336660 558788
rect 336596 558728 336646 558784
rect 336646 558728 336660 558784
rect 336596 558724 336660 558728
rect 338988 558784 339052 558788
rect 338988 558728 339002 558784
rect 339002 558728 339052 558784
rect 338988 558724 339052 558728
rect 339908 558784 339972 558788
rect 339908 558728 339922 558784
rect 339922 558728 339972 558784
rect 339908 558724 339972 558728
rect 341012 558784 341076 558788
rect 341012 558728 341026 558784
rect 341026 558728 341076 558784
rect 341012 558724 341076 558728
rect 342484 558784 342548 558788
rect 342484 558728 342534 558784
rect 342534 558728 342548 558784
rect 342484 558724 342548 558728
rect 343588 558724 343652 558788
rect 345980 558724 346044 558788
rect 346900 558784 346964 558788
rect 346900 558728 346950 558784
rect 346950 558728 346964 558784
rect 346900 558724 346964 558728
rect 348188 558724 348252 558788
rect 349476 558784 349540 558788
rect 349476 558728 349526 558784
rect 349526 558728 349540 558784
rect 349476 558724 349540 558728
rect 353524 558724 353588 558788
rect 357572 558724 357636 558788
rect 452700 558724 452764 558788
rect 459508 558724 459572 558788
rect 462084 558724 462148 558788
rect 463004 558784 463068 558788
rect 463004 558728 463018 558784
rect 463018 558728 463068 558784
rect 463004 558724 463068 558728
rect 464292 558784 464356 558788
rect 464292 558728 464342 558784
rect 464342 558728 464356 558784
rect 464292 558724 464356 558728
rect 465212 558784 465276 558788
rect 465212 558728 465226 558784
rect 465226 558728 465276 558784
rect 465212 558724 465276 558728
rect 469076 558724 469140 558788
rect 469996 558784 470060 558788
rect 469996 558728 470046 558784
rect 470046 558728 470060 558784
rect 469996 558724 470060 558728
rect 471284 558784 471348 558788
rect 471284 558728 471298 558784
rect 471298 558728 471348 558784
rect 471284 558724 471348 558728
rect 472204 558784 472268 558788
rect 472204 558728 472254 558784
rect 472254 558728 472268 558784
rect 472204 558724 472268 558728
rect 473492 558784 473556 558788
rect 473492 558728 473542 558784
rect 473542 558728 473556 558784
rect 473492 558724 473556 558728
rect 474780 558784 474844 558788
rect 474780 558728 474830 558784
rect 474830 558728 474844 558784
rect 474780 558724 474844 558728
rect 475516 558784 475580 558788
rect 475516 558728 475566 558784
rect 475566 558728 475580 558784
rect 475516 558724 475580 558728
rect 480484 558784 480548 558788
rect 480484 558728 480498 558784
rect 480498 558728 480548 558784
rect 480484 558724 480548 558728
rect 484716 558724 484780 558788
rect 101812 558648 101876 558652
rect 101812 558592 101862 558648
rect 101862 558592 101876 558648
rect 101812 558588 101876 558592
rect 197492 558588 197556 558652
rect 203748 558588 203812 558652
rect 209636 558588 209700 558652
rect 230612 558588 230676 558652
rect 231900 558648 231964 558652
rect 231900 558592 231914 558648
rect 231914 558592 231964 558648
rect 231900 558588 231964 558592
rect 234660 558648 234724 558652
rect 234660 558592 234674 558648
rect 234674 558592 234724 558648
rect 234660 558588 234724 558592
rect 323532 558588 323596 558652
rect 324820 558588 324884 558652
rect 326108 558588 326172 558652
rect 329604 558588 329668 558652
rect 330524 558648 330588 558652
rect 330524 558592 330538 558648
rect 330538 558592 330588 558648
rect 330524 558588 330588 558592
rect 356100 558648 356164 558652
rect 356100 558592 356114 558648
rect 356114 558592 356164 558648
rect 356100 558588 356164 558592
rect 456012 558648 456076 558652
rect 456012 558592 456062 558648
rect 456062 558592 456076 558648
rect 456012 558588 456076 558592
rect 457300 558588 457364 558652
rect 460796 558648 460860 558652
rect 460796 558592 460846 558648
rect 460846 558592 460860 558648
rect 460796 558588 460860 558592
rect 466500 558648 466564 558652
rect 466500 558592 466550 558648
rect 466550 558592 466564 558648
rect 466500 558588 466564 558592
rect 467788 558588 467852 558652
rect 483060 558648 483124 558652
rect 483060 558592 483074 558648
rect 483074 558592 483124 558648
rect 483060 558588 483124 558592
rect 488580 558648 488644 558652
rect 488580 558592 488594 558648
rect 488594 558592 488644 558648
rect 488580 558588 488644 558592
rect 198780 558512 198844 558516
rect 198780 558456 198794 558512
rect 198794 558456 198844 558512
rect 198780 558452 198844 558456
rect 200252 558512 200316 558516
rect 200252 558456 200266 558512
rect 200266 558456 200316 558512
rect 200252 558452 200316 558456
rect 237420 558512 237484 558516
rect 237420 558456 237434 558512
rect 237434 558456 237484 558512
rect 237420 558452 237484 558456
rect 238708 558512 238772 558516
rect 238708 558456 238758 558512
rect 238758 558456 238772 558512
rect 238708 558452 238772 558456
rect 317460 558512 317524 558516
rect 317460 558456 317474 558512
rect 317474 558456 317524 558512
rect 317460 558452 317524 558456
rect 337884 558452 337948 558516
rect 350580 558512 350644 558516
rect 350580 558456 350594 558512
rect 350594 558456 350644 558512
rect 350580 558452 350644 558456
rect 456564 558452 456628 558516
rect 481588 558512 481652 558516
rect 481588 558456 481638 558512
rect 481638 558456 481652 558512
rect 481588 558452 481652 558456
rect 487292 558452 487356 558516
rect 77708 558316 77772 558380
rect 83412 558316 83476 558380
rect 329788 558376 329852 558380
rect 329788 558320 329838 558376
rect 329838 558320 329852 558376
rect 329788 558316 329852 558320
rect 354812 558316 354876 558380
rect 455276 558316 455340 558380
rect 457484 558316 457548 558380
rect 458772 558316 458836 558380
rect 489132 558316 489196 558380
rect 74212 558180 74276 558244
rect 328868 558180 328932 558244
rect 332364 558180 332428 558244
rect 453804 558180 453868 558244
rect 459876 558180 459940 558244
rect 484164 558180 484228 558244
rect 486924 558180 486988 558244
rect 487844 558180 487908 558244
rect 68508 558044 68572 558108
rect 206140 558044 206204 558108
rect 238340 558044 238404 558108
rect 477356 558044 477420 558108
rect 478460 558044 478524 558108
rect 78628 557968 78692 557972
rect 78628 557912 78678 557968
rect 78678 557912 78692 557968
rect 78628 557908 78692 557912
rect 324084 557908 324148 557972
rect 479748 557908 479812 557972
rect 75132 557772 75196 557836
rect 76420 557772 76484 557836
rect 320220 557832 320284 557836
rect 320220 557776 320234 557832
rect 320234 557776 320284 557832
rect 320220 557772 320284 557776
rect 482140 557772 482204 557836
rect 72924 557636 72988 557700
rect 79916 557636 79980 557700
rect 93164 557636 93228 557700
rect 207060 557636 207124 557700
rect 208348 557636 208412 557700
rect 210372 557636 210436 557700
rect 344876 557636 344940 557700
rect 353156 557636 353220 557700
rect 451412 557696 451476 557700
rect 451412 557640 451426 557696
rect 451426 557640 451476 557696
rect 451412 557636 451476 557640
rect 475516 557636 475580 557700
rect 483612 557636 483676 557700
rect 71452 557500 71516 557564
rect 90956 557560 91020 557564
rect 90956 557504 91006 557560
rect 91006 557504 91020 557560
rect 90956 557500 91020 557504
rect 92060 557500 92124 557564
rect 93716 557560 93780 557564
rect 93716 557504 93766 557560
rect 93766 557504 93780 557560
rect 93716 557500 93780 557504
rect 95004 557500 95068 557564
rect 96476 557560 96540 557564
rect 96476 557504 96526 557560
rect 96526 557504 96540 557560
rect 96476 557500 96540 557504
rect 97764 557500 97828 557564
rect 99052 557500 99116 557564
rect 206876 557560 206940 557564
rect 206876 557504 206926 557560
rect 206926 557504 206940 557560
rect 206876 557500 206940 557504
rect 207980 557500 208044 557564
rect 209268 557500 209332 557564
rect 212396 557560 212460 557564
rect 212396 557504 212446 557560
rect 212446 557504 212460 557560
rect 212396 557500 212460 557504
rect 213500 557500 213564 557564
rect 214788 557500 214852 557564
rect 350948 557500 351012 557564
rect 354444 557500 354508 557564
rect 355548 557500 355612 557564
rect 356652 557500 356716 557564
rect 357940 557500 358004 557564
rect 352236 555520 352300 555524
rect 352236 555464 352250 555520
rect 352250 555464 352300 555520
rect 352236 555460 352300 555464
rect 359228 555460 359292 555524
rect 57468 539140 57532 539204
rect 57652 539004 57716 539068
rect 57836 393620 57900 393684
rect 59124 391444 59188 391508
rect 58204 389404 58268 389468
rect 57468 387228 57532 387292
rect 57652 378796 57716 378860
rect 57284 316024 57348 316028
rect 57284 315968 57334 316024
rect 57334 315968 57348 316024
rect 57284 315964 57348 315968
rect 57468 311476 57532 311540
rect 57284 306504 57348 306508
rect 57284 306448 57334 306504
rect 57334 306448 57348 306504
rect 57284 306444 57348 306448
rect 57836 305084 57900 305148
rect 57652 303044 57716 303108
rect 61148 300596 61212 300660
rect 61700 300596 61764 300660
rect 61148 299568 61212 299572
rect 61148 299512 61162 299568
rect 61162 299512 61212 299568
rect 61148 299508 61212 299512
rect 67404 177244 67468 177308
rect 67404 164188 67468 164252
rect 67404 125972 67468 126036
rect 67404 125564 67468 125628
rect 125548 76468 125612 76532
rect 57468 76196 57532 76260
rect 67588 76060 67652 76124
rect 115796 76332 115860 76396
rect 125548 76196 125612 76260
rect 115796 75924 115860 75988
rect 67588 75788 67652 75852
rect 125548 40564 125612 40628
rect 57652 40292 57716 40356
rect 67588 40156 67652 40220
rect 115796 40428 115860 40492
rect 125548 40292 125612 40356
rect 115796 40020 115860 40084
rect 67588 39884 67652 39948
rect 86908 29548 86972 29612
rect 57836 29276 57900 29340
rect 86908 29140 86972 29204
rect 115796 29412 115860 29476
rect 133828 29412 133892 29476
rect 133828 29140 133892 29204
rect 115796 29004 115860 29068
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 57835 686220 57901 686221
rect 57835 686156 57836 686220
rect 57900 686156 57901 686220
rect 57835 686155 57901 686156
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 57467 539204 57533 539205
rect 57467 539140 57468 539204
rect 57532 539140 57533 539204
rect 57467 539139 57533 539140
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 57470 387293 57530 539139
rect 57651 539068 57717 539069
rect 57651 539004 57652 539068
rect 57716 539004 57717 539068
rect 57651 539003 57717 539004
rect 57467 387292 57533 387293
rect 57467 387228 57468 387292
rect 57532 387228 57533 387292
rect 57467 387227 57533 387228
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 57654 378861 57714 539003
rect 57838 393685 57898 686155
rect 58203 673844 58269 673845
rect 58203 673780 58204 673844
rect 58268 673780 58269 673844
rect 58203 673779 58269 673780
rect 57835 393684 57901 393685
rect 57835 393620 57836 393684
rect 57900 393620 57901 393684
rect 57835 393619 57901 393620
rect 58206 389469 58266 673779
rect 58404 672054 59004 707102
rect 59123 697236 59189 697237
rect 59123 697172 59124 697236
rect 59188 697172 59189 697236
rect 59123 697171 59189 697172
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 654247 59004 671498
rect 58404 543000 59004 557000
rect 59126 391509 59186 697171
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 654247 62604 675098
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 654247 66204 678698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 654247 73404 685898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654247 77004 689498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 654247 80604 657098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 654247 84204 660698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 654247 91404 667898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 654247 95004 671498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 654247 98604 675098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 654247 102204 678698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 654247 109404 685898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654247 113004 689498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 654247 116604 657098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 654247 120204 660698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 654247 127404 667898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 654247 131004 671498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 654247 134604 675098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 654247 138204 678698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 129227 652900 129293 652901
rect 129227 652836 129228 652900
rect 129292 652836 129293 652900
rect 129227 652835 129293 652836
rect 133643 652900 133709 652901
rect 133643 652836 133644 652900
rect 133708 652836 133709 652900
rect 133643 652835 133709 652836
rect 129230 651130 129290 652835
rect 133646 651810 133706 652835
rect 128608 651070 129290 651130
rect 133573 651750 133706 651810
rect 133573 651100 133633 651750
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 136938 643254 137262 643276
rect 136938 643018 136982 643254
rect 137218 643018 137262 643254
rect 136938 642934 137262 643018
rect 136938 642698 136982 642934
rect 137218 642698 137262 642934
rect 136938 642676 137262 642698
rect 136938 639654 137262 639676
rect 136938 639418 136982 639654
rect 137218 639418 137262 639654
rect 136938 639334 137262 639418
rect 136938 639098 136982 639334
rect 137218 639098 137262 639334
rect 136938 639076 137262 639098
rect 136938 636054 137262 636076
rect 136938 635818 136982 636054
rect 137218 635818 137262 636054
rect 136938 635734 137262 635818
rect 136938 635498 136982 635734
rect 137218 635498 137262 635734
rect 136938 635476 137262 635498
rect 136938 632454 137262 632476
rect 136938 632218 136982 632454
rect 137218 632218 137262 632454
rect 136938 632134 137262 632218
rect 136938 631898 136982 632134
rect 137218 631898 137262 632134
rect 136938 631876 137262 631898
rect 136494 625254 136814 625276
rect 136494 625018 136536 625254
rect 136772 625018 136814 625254
rect 136494 624934 136814 625018
rect 136494 624698 136536 624934
rect 136772 624698 136814 624934
rect 136494 624676 136814 624698
rect 136494 621654 136814 621676
rect 136494 621418 136536 621654
rect 136772 621418 136814 621654
rect 136494 621334 136814 621418
rect 136494 621098 136536 621334
rect 136772 621098 136814 621334
rect 136494 621076 136814 621098
rect 136494 618054 136814 618076
rect 136494 617818 136536 618054
rect 136772 617818 136814 618054
rect 136494 617734 136814 617818
rect 136494 617498 136536 617734
rect 136772 617498 136814 617734
rect 136494 617476 136814 617498
rect 136494 614454 136814 614476
rect 136494 614218 136536 614454
rect 136772 614218 136814 614454
rect 136494 614134 136814 614218
rect 136494 613898 136536 614134
rect 136772 613898 136814 614134
rect 136494 613876 136814 613898
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 136938 607254 137262 607276
rect 136938 607018 136982 607254
rect 137218 607018 137262 607254
rect 136938 606934 137262 607018
rect 136938 606698 136982 606934
rect 137218 606698 137262 606934
rect 136938 606676 137262 606698
rect 136938 603654 137262 603676
rect 136938 603418 136982 603654
rect 137218 603418 137262 603654
rect 136938 603334 137262 603418
rect 136938 603098 136982 603334
rect 137218 603098 137262 603334
rect 136938 603076 137262 603098
rect 136938 600054 137262 600076
rect 136938 599818 136982 600054
rect 137218 599818 137262 600054
rect 136938 599734 137262 599818
rect 136938 599498 136982 599734
rect 137218 599498 137262 599734
rect 136938 599476 137262 599498
rect 136938 596454 137262 596476
rect 136938 596218 136982 596454
rect 137218 596218 137262 596454
rect 136938 596134 137262 596218
rect 136938 595898 136982 596134
rect 137218 595898 137262 596134
rect 136938 595876 137262 595898
rect 136494 589254 136814 589276
rect 136494 589018 136536 589254
rect 136772 589018 136814 589254
rect 136494 588934 136814 589018
rect 136494 588698 136536 588934
rect 136772 588698 136814 588934
rect 136494 588676 136814 588698
rect 136494 585654 136814 585676
rect 136494 585418 136536 585654
rect 136772 585418 136814 585654
rect 136494 585334 136814 585418
rect 136494 585098 136536 585334
rect 136772 585098 136814 585334
rect 136494 585076 136814 585098
rect 136494 582054 136814 582076
rect 136494 581818 136536 582054
rect 136772 581818 136814 582054
rect 136494 581734 136814 581818
rect 136494 581498 136536 581734
rect 136772 581498 136814 581734
rect 136494 581476 136814 581498
rect 136494 578454 136814 578476
rect 136494 578218 136536 578454
rect 136772 578218 136814 578454
rect 136494 578134 136814 578218
rect 136494 577898 136536 578134
rect 136772 577898 136814 578134
rect 136494 577876 136814 577898
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 136938 571254 137262 571276
rect 136938 571018 136982 571254
rect 137218 571018 137262 571254
rect 136938 570934 137262 571018
rect 136938 570698 136982 570934
rect 137218 570698 137262 570934
rect 136938 570676 137262 570698
rect 136938 567654 137262 567676
rect 136938 567418 136982 567654
rect 137218 567418 137262 567654
rect 136938 567334 137262 567418
rect 136938 567098 136982 567334
rect 137218 567098 137262 567334
rect 136938 567076 137262 567098
rect 136938 564054 137262 564076
rect 136938 563818 136982 564054
rect 137218 563818 137262 564054
rect 136938 563734 137262 563818
rect 136938 563498 136982 563734
rect 137218 563498 137262 563734
rect 136938 563476 137262 563498
rect 72374 560430 72672 560490
rect 73964 560430 74274 560490
rect 63542 560290 63833 560350
rect 66832 560290 67466 560350
rect 68000 560290 68570 560350
rect 69168 560290 69858 560350
rect 63542 558789 63602 560290
rect 67406 558925 67466 560290
rect 67403 558924 67469 558925
rect 67403 558860 67404 558924
rect 67468 558860 67469 558924
rect 67403 558859 67469 558860
rect 61699 558788 61765 558789
rect 61699 558724 61700 558788
rect 61764 558724 61765 558788
rect 61699 558723 61765 558724
rect 63539 558788 63605 558789
rect 63539 558724 63540 558788
rect 63604 558724 63605 558788
rect 63539 558723 63605 558724
rect 59123 391508 59189 391509
rect 59123 391444 59124 391508
rect 59188 391444 59189 391508
rect 59123 391443 59189 391444
rect 58203 389468 58269 389469
rect 58203 389404 58204 389468
rect 58268 389404 58269 389468
rect 58203 389403 58269 389404
rect 57651 378860 57717 378861
rect 57651 378796 57652 378860
rect 57716 378796 57717 378860
rect 57651 378795 57717 378796
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 57283 316028 57349 316029
rect 57283 315964 57284 316028
rect 57348 315964 57349 316028
rect 57283 315963 57349 315964
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 57286 306509 57346 315963
rect 57467 311540 57533 311541
rect 57467 311476 57468 311540
rect 57532 311476 57533 311540
rect 57467 311475 57533 311476
rect 57283 306508 57349 306509
rect 57283 306444 57284 306508
rect 57348 306444 57349 306508
rect 57283 306443 57349 306444
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 57470 76261 57530 311475
rect 57835 305148 57901 305149
rect 57835 305084 57836 305148
rect 57900 305084 57901 305148
rect 57835 305083 57901 305084
rect 57651 303108 57717 303109
rect 57651 303044 57652 303108
rect 57716 303044 57717 303108
rect 57651 303043 57717 303044
rect 57467 76260 57533 76261
rect 57467 76196 57468 76260
rect 57532 76196 57533 76260
rect 57467 76195 57533 76196
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 57654 40357 57714 303043
rect 57651 40356 57717 40357
rect 57651 40292 57652 40356
rect 57716 40292 57717 40356
rect 57651 40291 57717 40292
rect 57838 29341 57898 305083
rect 61702 300661 61762 558723
rect 68510 558109 68570 560290
rect 69798 558925 69858 560290
rect 70166 560290 70336 560350
rect 69795 558924 69861 558925
rect 69795 558860 69796 558924
rect 69860 558860 69861 558924
rect 69795 558859 69861 558860
rect 70166 558789 70226 560290
rect 70163 558788 70229 558789
rect 70163 558724 70164 558788
rect 70228 558724 70229 558788
rect 70163 558723 70229 558724
rect 68507 558108 68573 558109
rect 68507 558044 68508 558108
rect 68572 558044 68573 558108
rect 68507 558043 68573 558044
rect 71454 557565 71514 560350
rect 72374 558925 72434 560430
rect 72796 560290 72986 560350
rect 72371 558924 72437 558925
rect 72371 558860 72372 558924
rect 72436 558860 72437 558924
rect 72371 558859 72437 558860
rect 72926 557701 72986 560290
rect 73662 560290 73840 560350
rect 73662 558925 73722 560290
rect 73659 558924 73725 558925
rect 73659 558860 73660 558924
rect 73724 558860 73725 558924
rect 73659 558859 73725 558860
rect 74214 558245 74274 560430
rect 75870 560430 76176 560490
rect 77468 560430 77770 560490
rect 74950 558925 75010 560350
rect 75132 560290 75194 560350
rect 74947 558924 75013 558925
rect 74947 558860 74948 558924
rect 75012 558860 75013 558924
rect 74947 558859 75013 558860
rect 74211 558244 74277 558245
rect 74211 558180 74212 558244
rect 74276 558180 74277 558244
rect 74211 558179 74277 558180
rect 75134 557837 75194 560290
rect 75870 558925 75930 560430
rect 76300 560290 76482 560350
rect 75867 558924 75933 558925
rect 75867 558860 75868 558924
rect 75932 558860 75933 558924
rect 75867 558859 75933 558860
rect 76422 557837 76482 560290
rect 77314 559330 77374 560320
rect 77314 559270 77402 559330
rect 77342 558925 77402 559270
rect 77339 558924 77405 558925
rect 77339 558860 77340 558924
rect 77404 558860 77405 558924
rect 77339 558859 77405 558860
rect 77710 558381 77770 560430
rect 79366 560430 79680 560490
rect 82862 560430 83184 560490
rect 84476 560430 84762 560490
rect 78446 560290 78512 560350
rect 78446 558925 78506 560290
rect 78443 558924 78509 558925
rect 78443 558860 78444 558924
rect 78508 558860 78509 558924
rect 78443 558859 78509 558860
rect 77707 558380 77773 558381
rect 77707 558316 77708 558380
rect 77772 558316 77773 558380
rect 77707 558315 77773 558316
rect 78630 557973 78690 560350
rect 79366 558925 79426 560430
rect 79804 560290 79978 560350
rect 79363 558924 79429 558925
rect 79363 558860 79364 558924
rect 79428 558860 79429 558924
rect 79363 558859 79429 558860
rect 78627 557972 78693 557973
rect 78627 557908 78628 557972
rect 78692 557908 78693 557972
rect 78627 557907 78693 557908
rect 75131 557836 75197 557837
rect 75131 557772 75132 557836
rect 75196 557772 75197 557836
rect 75131 557771 75197 557772
rect 76419 557836 76485 557837
rect 76419 557772 76420 557836
rect 76484 557772 76485 557836
rect 76419 557771 76485 557772
rect 79918 557701 79978 560290
rect 80654 560290 80848 560350
rect 80654 558925 80714 560290
rect 80942 560010 81002 560320
rect 81758 560290 82016 560350
rect 80942 559950 81082 560010
rect 80651 558924 80717 558925
rect 80651 558860 80652 558924
rect 80716 558860 80717 558924
rect 80651 558859 80717 558860
rect 81022 558789 81082 559950
rect 81758 558789 81818 560290
rect 82126 558925 82186 560350
rect 82862 558925 82922 560430
rect 83308 560290 83474 560350
rect 82123 558924 82189 558925
rect 82123 558860 82124 558924
rect 82188 558860 82189 558924
rect 82123 558859 82189 558860
rect 82859 558924 82925 558925
rect 82859 558860 82860 558924
rect 82924 558860 82925 558924
rect 82859 558859 82925 558860
rect 81019 558788 81085 558789
rect 81019 558724 81020 558788
rect 81084 558724 81085 558788
rect 81019 558723 81085 558724
rect 81755 558788 81821 558789
rect 81755 558724 81756 558788
rect 81820 558724 81821 558788
rect 81755 558723 81821 558724
rect 83414 558381 83474 560290
rect 84150 560290 84352 560350
rect 84150 558789 84210 560290
rect 84702 558925 84762 560430
rect 86358 560430 86688 560490
rect 87980 560430 88258 560490
rect 85438 560290 85520 560350
rect 85438 558925 85498 560290
rect 85622 558925 85682 560350
rect 84699 558924 84765 558925
rect 84699 558860 84700 558924
rect 84764 558860 84765 558924
rect 84699 558859 84765 558860
rect 85435 558924 85501 558925
rect 85435 558860 85436 558924
rect 85500 558860 85501 558924
rect 85435 558859 85501 558860
rect 85619 558924 85685 558925
rect 85619 558860 85620 558924
rect 85684 558860 85685 558924
rect 85619 558859 85685 558860
rect 86358 558789 86418 560430
rect 86782 559330 86842 560320
rect 87826 560010 87886 560320
rect 87826 559950 87890 560010
rect 86726 559270 86842 559330
rect 86726 558925 86786 559270
rect 86723 558924 86789 558925
rect 86723 558860 86724 558924
rect 86788 558860 86789 558924
rect 86723 558859 86789 558860
rect 87830 558789 87890 559950
rect 88198 558925 88258 560430
rect 102734 560430 103040 560490
rect 106230 560430 106544 560490
rect 88934 560290 89024 560350
rect 88934 558925 88994 560290
rect 89118 558925 89178 560320
rect 90038 560290 90192 560350
rect 90316 560290 91018 560350
rect 90038 558925 90098 560290
rect 88195 558924 88261 558925
rect 88195 558860 88196 558924
rect 88260 558860 88261 558924
rect 88195 558859 88261 558860
rect 88931 558924 88997 558925
rect 88931 558860 88932 558924
rect 88996 558860 88997 558924
rect 88931 558859 88997 558860
rect 89115 558924 89181 558925
rect 89115 558860 89116 558924
rect 89180 558860 89181 558924
rect 89115 558859 89181 558860
rect 90035 558924 90101 558925
rect 90035 558860 90036 558924
rect 90100 558860 90101 558924
rect 90035 558859 90101 558860
rect 84147 558788 84213 558789
rect 84147 558724 84148 558788
rect 84212 558724 84213 558788
rect 84147 558723 84213 558724
rect 86355 558788 86421 558789
rect 86355 558724 86356 558788
rect 86420 558724 86421 558788
rect 86355 558723 86421 558724
rect 87827 558788 87893 558789
rect 87827 558724 87828 558788
rect 87892 558724 87893 558788
rect 87827 558723 87893 558724
rect 83411 558380 83477 558381
rect 83411 558316 83412 558380
rect 83476 558316 83477 558380
rect 83411 558315 83477 558316
rect 72923 557700 72989 557701
rect 72923 557636 72924 557700
rect 72988 557636 72989 557700
rect 72923 557635 72989 557636
rect 79915 557700 79981 557701
rect 79915 557636 79916 557700
rect 79980 557636 79981 557700
rect 79915 557635 79981 557636
rect 90958 557565 91018 560290
rect 91326 558925 91386 560350
rect 91484 560290 92122 560350
rect 91323 558924 91389 558925
rect 91323 558860 91324 558924
rect 91388 558860 91389 558924
rect 91323 558859 91389 558860
rect 92062 557565 92122 560290
rect 92498 560010 92558 560320
rect 92652 560290 93226 560350
rect 92430 559950 92558 560010
rect 92430 558925 92490 559950
rect 92427 558924 92493 558925
rect 92427 558860 92428 558924
rect 92492 558860 92493 558924
rect 92427 558859 92493 558860
rect 93166 557701 93226 560290
rect 93534 560290 93696 560350
rect 93534 558925 93594 560290
rect 93790 559330 93850 560320
rect 93718 559270 93850 559330
rect 94638 560290 94864 560350
rect 94988 560290 95066 560350
rect 93531 558924 93597 558925
rect 93531 558860 93532 558924
rect 93596 558860 93597 558924
rect 93531 558859 93597 558860
rect 93163 557700 93229 557701
rect 93163 557636 93164 557700
rect 93228 557636 93229 557700
rect 93163 557635 93229 557636
rect 93718 557565 93778 559270
rect 94638 558925 94698 560290
rect 94635 558924 94701 558925
rect 94635 558860 94636 558924
rect 94700 558860 94701 558924
rect 94635 558859 94701 558860
rect 95006 557565 95066 560290
rect 95374 560290 96032 560350
rect 96156 560290 96538 560350
rect 95374 558925 95434 560290
rect 95371 558924 95437 558925
rect 95371 558860 95372 558924
rect 95436 558860 95437 558924
rect 95371 558859 95437 558860
rect 96478 557565 96538 560290
rect 96662 560290 97200 560350
rect 97324 560290 97826 560350
rect 96662 558925 96722 560290
rect 96659 558924 96725 558925
rect 96659 558860 96660 558924
rect 96724 558860 96725 558924
rect 96659 558859 96725 558860
rect 97766 557565 97826 560290
rect 98318 558925 98378 560350
rect 98492 560290 99114 560350
rect 98315 558924 98381 558925
rect 98315 558860 98316 558924
rect 98380 558860 98381 558924
rect 98315 558859 98381 558860
rect 99054 557565 99114 560290
rect 99506 559330 99566 560320
rect 99660 560290 100218 560350
rect 99506 559270 99666 559330
rect 99606 558925 99666 559270
rect 100158 558925 100218 560290
rect 100342 560290 100704 560350
rect 100828 560290 101506 560350
rect 99603 558924 99669 558925
rect 99603 558860 99604 558924
rect 99668 558860 99669 558924
rect 99603 558859 99669 558860
rect 100155 558924 100221 558925
rect 100155 558860 100156 558924
rect 100220 558860 100221 558924
rect 100155 558859 100221 558860
rect 100342 558789 100402 560290
rect 101446 558789 101506 560290
rect 100339 558788 100405 558789
rect 100339 558724 100340 558788
rect 100404 558724 100405 558788
rect 100339 558723 100405 558724
rect 101443 558788 101509 558789
rect 101443 558724 101444 558788
rect 101508 558724 101509 558788
rect 101443 558723 101509 558724
rect 101814 558653 101874 560350
rect 101996 560290 102058 560350
rect 101998 558925 102058 560290
rect 102734 558925 102794 560430
rect 103164 560290 103346 560350
rect 103286 558925 103346 560290
rect 104022 560290 104208 560350
rect 104332 560290 104818 560350
rect 104022 558925 104082 560290
rect 104758 558925 104818 560290
rect 105310 560290 105376 560350
rect 105500 560290 106106 560350
rect 105310 558925 105370 560290
rect 106046 558925 106106 560290
rect 101995 558924 102061 558925
rect 101995 558860 101996 558924
rect 102060 558860 102061 558924
rect 101995 558859 102061 558860
rect 102731 558924 102797 558925
rect 102731 558860 102732 558924
rect 102796 558860 102797 558924
rect 102731 558859 102797 558860
rect 103283 558924 103349 558925
rect 103283 558860 103284 558924
rect 103348 558860 103349 558924
rect 103283 558859 103349 558860
rect 104019 558924 104085 558925
rect 104019 558860 104020 558924
rect 104084 558860 104085 558924
rect 104019 558859 104085 558860
rect 104755 558924 104821 558925
rect 104755 558860 104756 558924
rect 104820 558860 104821 558924
rect 104755 558859 104821 558860
rect 105307 558924 105373 558925
rect 105307 558860 105308 558924
rect 105372 558860 105373 558924
rect 105307 558859 105373 558860
rect 106043 558924 106109 558925
rect 106043 558860 106044 558924
rect 106108 558860 106109 558924
rect 106043 558859 106109 558860
rect 106230 558789 106290 560430
rect 106668 560290 107210 560350
rect 107150 558925 107210 560290
rect 107682 559330 107742 560320
rect 107836 560290 108498 560350
rect 107682 559270 107762 559330
rect 107702 558925 107762 559270
rect 108438 558925 108498 560290
rect 108622 560290 108880 560350
rect 109004 560290 109602 560350
rect 107147 558924 107213 558925
rect 107147 558860 107148 558924
rect 107212 558860 107213 558924
rect 107147 558859 107213 558860
rect 107699 558924 107765 558925
rect 107699 558860 107700 558924
rect 107764 558860 107765 558924
rect 107699 558859 107765 558860
rect 108435 558924 108501 558925
rect 108435 558860 108436 558924
rect 108500 558860 108501 558924
rect 108435 558859 108501 558860
rect 108622 558789 108682 560290
rect 109542 558925 109602 560290
rect 109539 558924 109605 558925
rect 109539 558860 109540 558924
rect 109604 558860 109605 558924
rect 109539 558859 109605 558860
rect 106227 558788 106293 558789
rect 106227 558724 106228 558788
rect 106292 558724 106293 558788
rect 106227 558723 106293 558724
rect 108619 558788 108685 558789
rect 108619 558724 108620 558788
rect 108684 558724 108685 558788
rect 108619 558723 108685 558724
rect 101811 558652 101877 558653
rect 101811 558588 101812 558652
rect 101876 558588 101877 558652
rect 101811 558587 101877 558588
rect 71451 557564 71517 557565
rect 71451 557500 71452 557564
rect 71516 557500 71517 557564
rect 71451 557499 71517 557500
rect 90955 557564 91021 557565
rect 90955 557500 90956 557564
rect 91020 557500 91021 557564
rect 90955 557499 91021 557500
rect 92059 557564 92125 557565
rect 92059 557500 92060 557564
rect 92124 557500 92125 557564
rect 92059 557499 92125 557500
rect 93715 557564 93781 557565
rect 93715 557500 93716 557564
rect 93780 557500 93781 557564
rect 93715 557499 93781 557500
rect 95003 557564 95069 557565
rect 95003 557500 95004 557564
rect 95068 557500 95069 557564
rect 95003 557499 95069 557500
rect 96475 557564 96541 557565
rect 96475 557500 96476 557564
rect 96540 557500 96541 557564
rect 96475 557499 96541 557500
rect 97763 557564 97829 557565
rect 97763 557500 97764 557564
rect 97828 557500 97829 557564
rect 97763 557499 97829 557500
rect 99051 557564 99117 557565
rect 99051 557500 99052 557564
rect 99116 557500 99117 557564
rect 99051 557499 99117 557500
rect 62004 543000 62604 557000
rect 65604 543000 66204 557000
rect 72804 543000 73404 557000
rect 76404 546054 77004 557000
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 543000 77004 545498
rect 80004 549654 80604 557000
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 543000 80604 549098
rect 83604 553254 84204 557000
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 543000 84204 552698
rect 90804 543000 91404 557000
rect 94404 543000 95004 557000
rect 98004 543000 98604 557000
rect 101604 543000 102204 557000
rect 108804 543000 109404 557000
rect 112404 546054 113004 557000
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 543000 113004 545498
rect 116004 549654 116604 557000
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 543000 116604 549098
rect 119604 553254 120204 557000
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 543000 120204 552698
rect 126804 543000 127404 557000
rect 130404 543000 131004 557000
rect 134004 543000 134604 557000
rect 137604 543000 138204 557000
rect 144804 543000 145404 577898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 543000 149004 545498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 543000 152604 549098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 543000 156204 552698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 164187 686356 164253 686357
rect 164187 686292 164188 686356
rect 164252 686292 164253 686356
rect 164187 686291 164253 686292
rect 164190 685949 164250 686291
rect 164187 685948 164253 685949
rect 164187 685884 164188 685948
rect 164252 685884 164253 685948
rect 164187 685883 164253 685884
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 543000 163404 559898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 543000 167004 563498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 543000 170604 567098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 543000 174204 570698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 183507 686492 183573 686493
rect 183507 686428 183508 686492
rect 183572 686428 183573 686492
rect 183507 686427 183573 686428
rect 183510 686221 183570 686427
rect 180804 686134 181404 686218
rect 183507 686220 183573 686221
rect 183507 686156 183508 686220
rect 183572 686156 183573 686220
rect 183507 686155 183573 686156
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 183507 674116 183573 674117
rect 183507 674052 183508 674116
rect 183572 674052 183573 674116
rect 183507 674051 183573 674052
rect 183510 673845 183570 674051
rect 183507 673844 183573 673845
rect 183507 673780 183508 673844
rect 183572 673780 183573 673844
rect 183507 673779 183573 673780
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 543000 181404 577898
rect 184404 654054 185004 689498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 654247 188604 657098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 654247 192204 660698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 654247 199404 667898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 654247 203004 671498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 654247 206604 675098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 654247 210204 678698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 654247 217404 685898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654247 221004 689498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 654247 224604 657098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 654247 228204 660698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 654247 235404 667898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 654247 239004 671498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 654247 242604 675098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 654247 246204 678698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 654247 253404 685898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654247 257004 689498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 654247 260604 657098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 654247 264204 660698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 259131 652900 259197 652901
rect 259131 652836 259132 652900
rect 259196 652836 259197 652900
rect 259131 652835 259197 652836
rect 263731 652900 263797 652901
rect 263731 652836 263732 652900
rect 263796 652836 263797 652900
rect 263731 652835 263797 652836
rect 259134 651130 259194 652835
rect 263734 651130 263794 652835
rect 258608 651070 259194 651130
rect 263603 651070 263794 651130
rect 266938 643254 267262 643276
rect 266938 643018 266982 643254
rect 267218 643018 267262 643254
rect 266938 642934 267262 643018
rect 266938 642698 266982 642934
rect 267218 642698 267262 642934
rect 266938 642676 267262 642698
rect 266938 639654 267262 639676
rect 266938 639418 266982 639654
rect 267218 639418 267262 639654
rect 266938 639334 267262 639418
rect 266938 639098 266982 639334
rect 267218 639098 267262 639334
rect 266938 639076 267262 639098
rect 266938 636054 267262 636076
rect 266938 635818 266982 636054
rect 267218 635818 267262 636054
rect 266938 635734 267262 635818
rect 266938 635498 266982 635734
rect 267218 635498 267262 635734
rect 266938 635476 267262 635498
rect 266938 632454 267262 632476
rect 266938 632218 266982 632454
rect 267218 632218 267262 632454
rect 266938 632134 267262 632218
rect 266938 631898 266982 632134
rect 267218 631898 267262 632134
rect 266938 631876 267262 631898
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 266494 625254 266814 625276
rect 266494 625018 266536 625254
rect 266772 625018 266814 625254
rect 266494 624934 266814 625018
rect 266494 624698 266536 624934
rect 266772 624698 266814 624934
rect 266494 624676 266814 624698
rect 266494 621654 266814 621676
rect 266494 621418 266536 621654
rect 266772 621418 266814 621654
rect 266494 621334 266814 621418
rect 266494 621098 266536 621334
rect 266772 621098 266814 621334
rect 266494 621076 266814 621098
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 266494 618054 266814 618076
rect 266494 617818 266536 618054
rect 266772 617818 266814 618054
rect 266494 617734 266814 617818
rect 266494 617498 266536 617734
rect 266772 617498 266814 617734
rect 266494 617476 266814 617498
rect 266494 614454 266814 614476
rect 266494 614218 266536 614454
rect 266772 614218 266814 614454
rect 266494 614134 266814 614218
rect 266494 613898 266536 614134
rect 266772 613898 266814 614134
rect 266494 613876 266814 613898
rect 266938 607254 267262 607276
rect 266938 607018 266982 607254
rect 267218 607018 267262 607254
rect 266938 606934 267262 607018
rect 266938 606698 266982 606934
rect 267218 606698 267262 606934
rect 266938 606676 267262 606698
rect 266938 603654 267262 603676
rect 266938 603418 266982 603654
rect 267218 603418 267262 603654
rect 266938 603334 267262 603418
rect 266938 603098 266982 603334
rect 267218 603098 267262 603334
rect 266938 603076 267262 603098
rect 266938 600054 267262 600076
rect 266938 599818 266982 600054
rect 267218 599818 267262 600054
rect 266938 599734 267262 599818
rect 266938 599498 266982 599734
rect 267218 599498 267262 599734
rect 266938 599476 267262 599498
rect 266938 596454 267262 596476
rect 266938 596218 266982 596454
rect 267218 596218 267262 596454
rect 266938 596134 267262 596218
rect 266938 595898 266982 596134
rect 267218 595898 267262 596134
rect 266938 595876 267262 595898
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 266494 589254 266814 589276
rect 266494 589018 266536 589254
rect 266772 589018 266814 589254
rect 266494 588934 266814 589018
rect 266494 588698 266536 588934
rect 266772 588698 266814 588934
rect 266494 588676 266814 588698
rect 266494 585654 266814 585676
rect 266494 585418 266536 585654
rect 266772 585418 266814 585654
rect 266494 585334 266814 585418
rect 266494 585098 266536 585334
rect 266772 585098 266814 585334
rect 266494 585076 266814 585098
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 266494 582054 266814 582076
rect 266494 581818 266536 582054
rect 266772 581818 266814 582054
rect 266494 581734 266814 581818
rect 266494 581498 266536 581734
rect 266772 581498 266814 581734
rect 266494 581476 266814 581498
rect 266494 578454 266814 578476
rect 266494 578218 266536 578454
rect 266772 578218 266814 578454
rect 266494 578134 266814 578218
rect 266494 577898 266536 578134
rect 266772 577898 266814 578134
rect 266494 577876 266814 577898
rect 266938 571254 267262 571276
rect 266938 571018 266982 571254
rect 267218 571018 267262 571254
rect 266938 570934 267262 571018
rect 266938 570698 266982 570934
rect 267218 570698 267262 570934
rect 266938 570676 267262 570698
rect 266938 567654 267262 567676
rect 266938 567418 266982 567654
rect 267218 567418 267262 567654
rect 266938 567334 267262 567418
rect 266938 567098 266982 567334
rect 267218 567098 267262 567334
rect 266938 567076 267262 567098
rect 266938 564054 267262 564076
rect 266938 563818 266982 564054
rect 267218 563818 267262 564054
rect 266938 563734 267262 563818
rect 266938 563498 266982 563734
rect 267218 563498 267262 563734
rect 266938 563476 267262 563498
rect 201504 560430 201786 560490
rect 193814 558925 193874 560350
rect 196206 560290 196832 560350
rect 197494 560290 198000 560350
rect 198782 560290 199168 560350
rect 200254 560290 200336 560350
rect 193811 558924 193877 558925
rect 193811 558860 193812 558924
rect 193876 558860 193877 558924
rect 193811 558859 193877 558860
rect 196206 558789 196266 560290
rect 196203 558788 196269 558789
rect 196203 558724 196204 558788
rect 196268 558724 196269 558788
rect 196203 558723 196269 558724
rect 197494 558653 197554 560290
rect 197491 558652 197557 558653
rect 197491 558588 197492 558652
rect 197556 558588 197557 558652
rect 197491 558587 197557 558588
rect 198782 558517 198842 560290
rect 200254 558517 200314 560290
rect 201726 558789 201786 560430
rect 207062 560430 207344 560490
rect 210558 560430 210848 560490
rect 221046 560430 221360 560490
rect 270804 560454 271404 595898
rect 202462 560290 202672 560350
rect 202462 558789 202522 560290
rect 202766 559330 202826 560320
rect 202646 559270 202826 559330
rect 203750 560290 203840 560350
rect 202646 558925 202706 559270
rect 202643 558924 202709 558925
rect 202643 558860 202644 558924
rect 202708 558860 202709 558924
rect 202643 558859 202709 558860
rect 201723 558788 201789 558789
rect 201723 558724 201724 558788
rect 201788 558724 201789 558788
rect 201723 558723 201789 558724
rect 202459 558788 202525 558789
rect 202459 558724 202460 558788
rect 202524 558724 202525 558788
rect 202459 558723 202525 558724
rect 203750 558653 203810 560290
rect 203934 558925 203994 560320
rect 204854 560290 205008 560350
rect 205132 560290 205466 560350
rect 203931 558924 203997 558925
rect 203931 558860 203932 558924
rect 203996 558860 203997 558924
rect 203931 558859 203997 558860
rect 204854 558789 204914 560290
rect 205406 558925 205466 560290
rect 205403 558924 205469 558925
rect 205403 558860 205404 558924
rect 205468 558860 205469 558924
rect 205403 558859 205469 558860
rect 204851 558788 204917 558789
rect 204851 558724 204852 558788
rect 204916 558724 204917 558788
rect 204851 558723 204917 558724
rect 203747 558652 203813 558653
rect 203747 558588 203748 558652
rect 203812 558588 203813 558652
rect 203747 558587 203813 558588
rect 198779 558516 198845 558517
rect 198779 558452 198780 558516
rect 198844 558452 198845 558516
rect 198779 558451 198845 558452
rect 200251 558516 200317 558517
rect 200251 558452 200252 558516
rect 200316 558452 200317 558516
rect 200251 558451 200317 558452
rect 206142 558109 206202 560350
rect 206300 560290 206938 560350
rect 206139 558108 206205 558109
rect 206139 558044 206140 558108
rect 206204 558044 206205 558108
rect 206139 558043 206205 558044
rect 206878 557565 206938 560290
rect 207062 557701 207122 560430
rect 207468 560290 208042 560350
rect 207059 557700 207125 557701
rect 207059 557636 207060 557700
rect 207124 557636 207125 557700
rect 207059 557635 207125 557636
rect 207982 557565 208042 560290
rect 208350 560290 208512 560350
rect 208636 560290 209330 560350
rect 208350 557701 208410 560290
rect 208347 557700 208413 557701
rect 208347 557636 208348 557700
rect 208412 557636 208413 557700
rect 208347 557635 208413 557636
rect 209270 557565 209330 560290
rect 209638 558653 209698 560350
rect 209804 560290 210434 560350
rect 209635 558652 209701 558653
rect 209635 558588 209636 558652
rect 209700 558588 209701 558652
rect 209635 558587 209701 558588
rect 210374 557701 210434 560290
rect 210558 559877 210618 560430
rect 210942 560010 211002 560320
rect 211846 560290 212016 560350
rect 212140 560290 212458 560350
rect 211107 560012 211173 560013
rect 211107 560010 211108 560012
rect 210942 559950 211108 560010
rect 211107 559948 211108 559950
rect 211172 559948 211173 560012
rect 211107 559947 211173 559948
rect 210555 559876 210621 559877
rect 210555 559812 210556 559876
rect 210620 559812 210621 559876
rect 210555 559811 210621 559812
rect 211846 558925 211906 560290
rect 211843 558924 211909 558925
rect 211843 558860 211844 558924
rect 211908 558860 211909 558924
rect 211843 558859 211909 558860
rect 210371 557700 210437 557701
rect 210371 557636 210372 557700
rect 210436 557636 210437 557700
rect 210371 557635 210437 557636
rect 212398 557565 212458 560290
rect 213134 558925 213194 560350
rect 213308 560290 213562 560350
rect 213131 558924 213197 558925
rect 213131 558860 213132 558924
rect 213196 558860 213197 558924
rect 213131 558859 213197 558860
rect 213502 557565 213562 560290
rect 214054 560290 214352 560350
rect 214476 560290 214850 560350
rect 214054 558925 214114 560290
rect 214051 558924 214117 558925
rect 214051 558860 214052 558924
rect 214116 558860 214117 558924
rect 214051 558859 214117 558860
rect 214790 557565 214850 560290
rect 215342 560290 215520 560350
rect 215644 560290 216322 560350
rect 215342 558789 215402 560290
rect 216262 558925 216322 560290
rect 216259 558924 216325 558925
rect 216259 558860 216260 558924
rect 216324 558860 216325 558924
rect 216259 558859 216325 558860
rect 216630 558789 216690 560350
rect 216812 560290 217426 560350
rect 217366 558789 217426 560290
rect 217550 560290 217856 560350
rect 217550 558925 217610 560290
rect 217950 559330 218010 560320
rect 217918 559270 218010 559330
rect 218838 560290 219024 560350
rect 217918 558925 217978 559270
rect 218838 558925 218898 560290
rect 219118 560010 219178 560320
rect 220126 560290 220192 560350
rect 220316 560290 220738 560350
rect 219118 559950 219266 560010
rect 219206 558925 219266 559950
rect 220126 558925 220186 560290
rect 220678 558925 220738 560290
rect 221046 558925 221106 560430
rect 221484 560290 222026 560350
rect 221966 558925 222026 560290
rect 222334 560290 222528 560350
rect 222652 560290 223314 560350
rect 222334 558925 222394 560290
rect 223254 558925 223314 560290
rect 223622 560290 223696 560350
rect 223820 560290 224418 560350
rect 217547 558924 217613 558925
rect 217547 558860 217548 558924
rect 217612 558860 217613 558924
rect 217547 558859 217613 558860
rect 217915 558924 217981 558925
rect 217915 558860 217916 558924
rect 217980 558860 217981 558924
rect 217915 558859 217981 558860
rect 218835 558924 218901 558925
rect 218835 558860 218836 558924
rect 218900 558860 218901 558924
rect 218835 558859 218901 558860
rect 219203 558924 219269 558925
rect 219203 558860 219204 558924
rect 219268 558860 219269 558924
rect 219203 558859 219269 558860
rect 220123 558924 220189 558925
rect 220123 558860 220124 558924
rect 220188 558860 220189 558924
rect 220123 558859 220189 558860
rect 220675 558924 220741 558925
rect 220675 558860 220676 558924
rect 220740 558860 220741 558924
rect 220675 558859 220741 558860
rect 221043 558924 221109 558925
rect 221043 558860 221044 558924
rect 221108 558860 221109 558924
rect 221043 558859 221109 558860
rect 221963 558924 222029 558925
rect 221963 558860 221964 558924
rect 222028 558860 222029 558924
rect 221963 558859 222029 558860
rect 222331 558924 222397 558925
rect 222331 558860 222332 558924
rect 222396 558860 222397 558924
rect 222331 558859 222397 558860
rect 223251 558924 223317 558925
rect 223251 558860 223252 558924
rect 223316 558860 223317 558924
rect 223251 558859 223317 558860
rect 223622 558789 223682 560290
rect 224358 558925 224418 560290
rect 224542 560290 224864 560350
rect 224988 560290 225706 560350
rect 224355 558924 224421 558925
rect 224355 558860 224356 558924
rect 224420 558860 224421 558924
rect 224355 558859 224421 558860
rect 224542 558789 224602 560290
rect 225646 558789 225706 560290
rect 225830 560290 226032 560350
rect 225830 558925 225890 560290
rect 226126 560010 226186 560320
rect 227118 560290 227200 560350
rect 227324 560290 227546 560350
rect 226126 559950 226258 560010
rect 226198 558925 226258 559950
rect 227118 558925 227178 560290
rect 227486 558925 227546 560290
rect 227854 560290 228368 560350
rect 228492 560290 228834 560350
rect 225827 558924 225893 558925
rect 225827 558860 225828 558924
rect 225892 558860 225893 558924
rect 225827 558859 225893 558860
rect 226195 558924 226261 558925
rect 226195 558860 226196 558924
rect 226260 558860 226261 558924
rect 226195 558859 226261 558860
rect 227115 558924 227181 558925
rect 227115 558860 227116 558924
rect 227180 558860 227181 558924
rect 227115 558859 227181 558860
rect 227483 558924 227549 558925
rect 227483 558860 227484 558924
rect 227548 558860 227549 558924
rect 227483 558859 227549 558860
rect 227854 558789 227914 560290
rect 228774 558925 228834 560290
rect 229506 560010 229566 560320
rect 229660 560290 230306 560350
rect 229506 559950 229570 560010
rect 229510 558925 229570 559950
rect 230246 558925 230306 560290
rect 230614 560290 230704 560350
rect 228771 558924 228837 558925
rect 228771 558860 228772 558924
rect 228836 558860 228837 558924
rect 228771 558859 228837 558860
rect 229507 558924 229573 558925
rect 229507 558860 229508 558924
rect 229572 558860 229573 558924
rect 229507 558859 229573 558860
rect 230243 558924 230309 558925
rect 230243 558860 230244 558924
rect 230308 558860 230309 558924
rect 230243 558859 230309 558860
rect 215339 558788 215405 558789
rect 215339 558724 215340 558788
rect 215404 558724 215405 558788
rect 215339 558723 215405 558724
rect 216627 558788 216693 558789
rect 216627 558724 216628 558788
rect 216692 558724 216693 558788
rect 216627 558723 216693 558724
rect 217363 558788 217429 558789
rect 217363 558724 217364 558788
rect 217428 558724 217429 558788
rect 217363 558723 217429 558724
rect 223619 558788 223685 558789
rect 223619 558724 223620 558788
rect 223684 558724 223685 558788
rect 223619 558723 223685 558724
rect 224539 558788 224605 558789
rect 224539 558724 224540 558788
rect 224604 558724 224605 558788
rect 224539 558723 224605 558724
rect 225643 558788 225709 558789
rect 225643 558724 225644 558788
rect 225708 558724 225709 558788
rect 225643 558723 225709 558724
rect 227851 558788 227917 558789
rect 227851 558724 227852 558788
rect 227916 558724 227917 558788
rect 227851 558723 227917 558724
rect 230614 558653 230674 560290
rect 230798 558925 230858 560320
rect 231842 559330 231902 560320
rect 231996 560290 232698 560350
rect 231842 559270 231962 559330
rect 230795 558924 230861 558925
rect 230795 558860 230796 558924
rect 230860 558860 230861 558924
rect 230795 558859 230861 558860
rect 231902 558653 231962 559270
rect 232638 558789 232698 560290
rect 232822 560290 233040 560350
rect 232822 558925 232882 560290
rect 233134 559330 233194 560320
rect 233006 559270 233194 559330
rect 233558 560290 234208 560350
rect 234332 560290 234538 560350
rect 233006 558925 233066 559270
rect 232819 558924 232885 558925
rect 232819 558860 232820 558924
rect 232884 558860 232885 558924
rect 232819 558859 232885 558860
rect 233003 558924 233069 558925
rect 233003 558860 233004 558924
rect 233068 558860 233069 558924
rect 233003 558859 233069 558860
rect 233558 558789 233618 560290
rect 234478 558925 234538 560290
rect 234662 560290 235376 560350
rect 235500 560290 235826 560350
rect 234475 558924 234541 558925
rect 234475 558860 234476 558924
rect 234540 558860 234541 558924
rect 234475 558859 234541 558860
rect 232635 558788 232701 558789
rect 232635 558724 232636 558788
rect 232700 558724 232701 558788
rect 232635 558723 232701 558724
rect 233555 558788 233621 558789
rect 233555 558724 233556 558788
rect 233620 558724 233621 558788
rect 233555 558723 233621 558724
rect 234662 558653 234722 560290
rect 235766 558925 235826 560290
rect 236134 560290 236544 560350
rect 236668 560290 237298 560350
rect 235763 558924 235829 558925
rect 235763 558860 235764 558924
rect 235828 558860 235829 558924
rect 235763 558859 235829 558860
rect 236134 558789 236194 560290
rect 237238 558925 237298 560290
rect 237422 560290 237712 560350
rect 237836 560290 238402 560350
rect 237235 558924 237301 558925
rect 237235 558860 237236 558924
rect 237300 558860 237301 558924
rect 237235 558859 237301 558860
rect 236131 558788 236197 558789
rect 236131 558724 236132 558788
rect 236196 558724 236197 558788
rect 236131 558723 236197 558724
rect 230611 558652 230677 558653
rect 230611 558588 230612 558652
rect 230676 558588 230677 558652
rect 230611 558587 230677 558588
rect 231899 558652 231965 558653
rect 231899 558588 231900 558652
rect 231964 558588 231965 558652
rect 231899 558587 231965 558588
rect 234659 558652 234725 558653
rect 234659 558588 234660 558652
rect 234724 558588 234725 558652
rect 234659 558587 234725 558588
rect 237422 558517 237482 560290
rect 237419 558516 237485 558517
rect 237419 558452 237420 558516
rect 237484 558452 237485 558516
rect 237419 558451 237485 558452
rect 238342 558109 238402 560290
rect 238710 560290 238880 560350
rect 239004 560290 239690 560350
rect 238710 558517 238770 560290
rect 239630 558925 239690 560290
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 239627 558924 239693 558925
rect 239627 558860 239628 558924
rect 239692 558860 239693 558924
rect 239627 558859 239693 558860
rect 238707 558516 238773 558517
rect 238707 558452 238708 558516
rect 238772 558452 238773 558516
rect 238707 558451 238773 558452
rect 238339 558108 238405 558109
rect 238339 558044 238340 558108
rect 238404 558044 238405 558108
rect 238339 558043 238405 558044
rect 206875 557564 206941 557565
rect 206875 557500 206876 557564
rect 206940 557500 206941 557564
rect 206875 557499 206941 557500
rect 207979 557564 208045 557565
rect 207979 557500 207980 557564
rect 208044 557500 208045 557564
rect 207979 557499 208045 557500
rect 209267 557564 209333 557565
rect 209267 557500 209268 557564
rect 209332 557500 209333 557564
rect 209267 557499 209333 557500
rect 212395 557564 212461 557565
rect 212395 557500 212396 557564
rect 212460 557500 212461 557564
rect 212395 557499 212461 557500
rect 213499 557564 213565 557565
rect 213499 557500 213500 557564
rect 213564 557500 213565 557564
rect 213499 557499 213565 557500
rect 214787 557564 214853 557565
rect 214787 557500 214788 557564
rect 214852 557500 214853 557564
rect 214787 557499 214853 557500
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 543000 185004 545498
rect 188004 549654 188604 557000
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 543000 188604 549098
rect 191604 553254 192204 557000
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 543000 192204 552698
rect 198804 543000 199404 557000
rect 202404 543000 203004 557000
rect 206004 543000 206604 557000
rect 209604 543000 210204 557000
rect 216804 543000 217404 557000
rect 220404 546054 221004 557000
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 543000 221004 545498
rect 224004 549654 224604 557000
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 543000 224604 549098
rect 227604 553254 228204 557000
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 543000 228204 552698
rect 234804 543000 235404 557000
rect 238404 543000 239004 557000
rect 242004 543000 242604 557000
rect 245604 543000 246204 557000
rect 252804 543000 253404 557000
rect 256404 546054 257004 557000
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 543000 257004 545498
rect 260004 549654 260604 557000
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 543000 260604 549098
rect 263604 553254 264204 557000
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 543000 264204 552698
rect 270804 543000 271404 559898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 543000 275004 563498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 543000 278604 567098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 543000 282204 570698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 79568 535254 79888 535276
rect 79568 535018 79610 535254
rect 79846 535018 79888 535254
rect 79568 534934 79888 535018
rect 79568 534698 79610 534934
rect 79846 534698 79888 534934
rect 79568 534676 79888 534698
rect 79568 531654 79888 531676
rect 79568 531418 79610 531654
rect 79846 531418 79888 531654
rect 79568 531334 79888 531418
rect 79568 531098 79610 531334
rect 79846 531098 79888 531334
rect 79568 531076 79888 531098
rect 79568 528054 79888 528076
rect 79568 527818 79610 528054
rect 79846 527818 79888 528054
rect 79568 527734 79888 527818
rect 79568 527498 79610 527734
rect 79846 527498 79888 527734
rect 79568 527476 79888 527498
rect 79568 524454 79888 524476
rect 79568 524218 79610 524454
rect 79846 524218 79888 524454
rect 79568 524134 79888 524218
rect 79568 523898 79610 524134
rect 79846 523898 79888 524134
rect 79568 523876 79888 523898
rect 64208 517254 64528 517276
rect 64208 517018 64250 517254
rect 64486 517018 64528 517254
rect 64208 516934 64528 517018
rect 64208 516698 64250 516934
rect 64486 516698 64528 516934
rect 64208 516676 64528 516698
rect 64208 513654 64528 513676
rect 64208 513418 64250 513654
rect 64486 513418 64528 513654
rect 64208 513334 64528 513418
rect 64208 513098 64250 513334
rect 64486 513098 64528 513334
rect 64208 513076 64528 513098
rect 64208 510054 64528 510076
rect 64208 509818 64250 510054
rect 64486 509818 64528 510054
rect 64208 509734 64528 509818
rect 64208 509498 64250 509734
rect 64486 509498 64528 509734
rect 64208 509476 64528 509498
rect 64208 506454 64528 506476
rect 64208 506218 64250 506454
rect 64486 506218 64528 506454
rect 64208 506134 64528 506218
rect 64208 505898 64250 506134
rect 64486 505898 64528 506134
rect 64208 505876 64528 505898
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 79568 499254 79888 499276
rect 79568 499018 79610 499254
rect 79846 499018 79888 499254
rect 79568 498934 79888 499018
rect 79568 498698 79610 498934
rect 79846 498698 79888 498934
rect 79568 498676 79888 498698
rect 79568 495654 79888 495676
rect 79568 495418 79610 495654
rect 79846 495418 79888 495654
rect 79568 495334 79888 495418
rect 79568 495098 79610 495334
rect 79846 495098 79888 495334
rect 79568 495076 79888 495098
rect 79568 492054 79888 492076
rect 79568 491818 79610 492054
rect 79846 491818 79888 492054
rect 79568 491734 79888 491818
rect 79568 491498 79610 491734
rect 79846 491498 79888 491734
rect 79568 491476 79888 491498
rect 79568 488454 79888 488476
rect 79568 488218 79610 488454
rect 79846 488218 79888 488454
rect 79568 488134 79888 488218
rect 79568 487898 79610 488134
rect 79846 487898 79888 488134
rect 79568 487876 79888 487898
rect 64208 481254 64528 481276
rect 64208 481018 64250 481254
rect 64486 481018 64528 481254
rect 64208 480934 64528 481018
rect 64208 480698 64250 480934
rect 64486 480698 64528 480934
rect 64208 480676 64528 480698
rect 64208 477654 64528 477676
rect 64208 477418 64250 477654
rect 64486 477418 64528 477654
rect 64208 477334 64528 477418
rect 64208 477098 64250 477334
rect 64486 477098 64528 477334
rect 64208 477076 64528 477098
rect 64208 474054 64528 474076
rect 64208 473818 64250 474054
rect 64486 473818 64528 474054
rect 64208 473734 64528 473818
rect 64208 473498 64250 473734
rect 64486 473498 64528 473734
rect 64208 473476 64528 473498
rect 64208 470454 64528 470476
rect 64208 470218 64250 470454
rect 64486 470218 64528 470454
rect 64208 470134 64528 470218
rect 64208 469898 64250 470134
rect 64486 469898 64528 470134
rect 64208 469876 64528 469898
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 79568 463254 79888 463276
rect 79568 463018 79610 463254
rect 79846 463018 79888 463254
rect 79568 462934 79888 463018
rect 79568 462698 79610 462934
rect 79846 462698 79888 462934
rect 79568 462676 79888 462698
rect 79568 459654 79888 459676
rect 79568 459418 79610 459654
rect 79846 459418 79888 459654
rect 79568 459334 79888 459418
rect 79568 459098 79610 459334
rect 79846 459098 79888 459334
rect 79568 459076 79888 459098
rect 79568 456054 79888 456076
rect 79568 455818 79610 456054
rect 79846 455818 79888 456054
rect 79568 455734 79888 455818
rect 79568 455498 79610 455734
rect 79846 455498 79888 455734
rect 79568 455476 79888 455498
rect 79568 452454 79888 452476
rect 79568 452218 79610 452454
rect 79846 452218 79888 452454
rect 79568 452134 79888 452218
rect 79568 451898 79610 452134
rect 79846 451898 79888 452134
rect 79568 451876 79888 451898
rect 64208 445254 64528 445276
rect 64208 445018 64250 445254
rect 64486 445018 64528 445254
rect 64208 444934 64528 445018
rect 64208 444698 64250 444934
rect 64486 444698 64528 444934
rect 64208 444676 64528 444698
rect 64208 441654 64528 441676
rect 64208 441418 64250 441654
rect 64486 441418 64528 441654
rect 64208 441334 64528 441418
rect 64208 441098 64250 441334
rect 64486 441098 64528 441334
rect 64208 441076 64528 441098
rect 64208 438054 64528 438076
rect 64208 437818 64250 438054
rect 64486 437818 64528 438054
rect 64208 437734 64528 437818
rect 64208 437498 64250 437734
rect 64486 437498 64528 437734
rect 64208 437476 64528 437498
rect 64208 434454 64528 434476
rect 64208 434218 64250 434454
rect 64486 434218 64528 434454
rect 64208 434134 64528 434218
rect 64208 433898 64250 434134
rect 64486 433898 64528 434134
rect 64208 433876 64528 433898
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 79568 427254 79888 427276
rect 79568 427018 79610 427254
rect 79846 427018 79888 427254
rect 79568 426934 79888 427018
rect 79568 426698 79610 426934
rect 79846 426698 79888 426934
rect 79568 426676 79888 426698
rect 79568 423654 79888 423676
rect 79568 423418 79610 423654
rect 79846 423418 79888 423654
rect 79568 423334 79888 423418
rect 79568 423098 79610 423334
rect 79846 423098 79888 423334
rect 79568 423076 79888 423098
rect 79568 420054 79888 420076
rect 79568 419818 79610 420054
rect 79846 419818 79888 420054
rect 79568 419734 79888 419818
rect 79568 419498 79610 419734
rect 79846 419498 79888 419734
rect 79568 419476 79888 419498
rect 79568 416454 79888 416476
rect 79568 416218 79610 416454
rect 79846 416218 79888 416454
rect 79568 416134 79888 416218
rect 79568 415898 79610 416134
rect 79846 415898 79888 416134
rect 79568 415876 79888 415898
rect 64208 409254 64528 409276
rect 64208 409018 64250 409254
rect 64486 409018 64528 409254
rect 64208 408934 64528 409018
rect 64208 408698 64250 408934
rect 64486 408698 64528 408934
rect 64208 408676 64528 408698
rect 64208 405654 64528 405676
rect 64208 405418 64250 405654
rect 64486 405418 64528 405654
rect 64208 405334 64528 405418
rect 64208 405098 64250 405334
rect 64486 405098 64528 405334
rect 64208 405076 64528 405098
rect 64208 402054 64528 402076
rect 64208 401818 64250 402054
rect 64486 401818 64528 402054
rect 64208 401734 64528 401818
rect 64208 401498 64250 401734
rect 64486 401498 64528 401734
rect 64208 401476 64528 401498
rect 64208 398454 64528 398476
rect 64208 398218 64250 398454
rect 64486 398218 64528 398454
rect 64208 398134 64528 398218
rect 64208 397898 64250 398134
rect 64486 397898 64528 398134
rect 64208 397876 64528 397898
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 79568 391254 79888 391276
rect 79568 391018 79610 391254
rect 79846 391018 79888 391254
rect 79568 390934 79888 391018
rect 79568 390698 79610 390934
rect 79846 390698 79888 390934
rect 79568 390676 79888 390698
rect 79568 387654 79888 387676
rect 79568 387418 79610 387654
rect 79846 387418 79888 387654
rect 79568 387334 79888 387418
rect 79568 387098 79610 387334
rect 79846 387098 79888 387334
rect 79568 387076 79888 387098
rect 79568 384054 79888 384076
rect 79568 383818 79610 384054
rect 79846 383818 79888 384054
rect 79568 383734 79888 383818
rect 79568 383498 79610 383734
rect 79846 383498 79888 383734
rect 79568 383476 79888 383498
rect 79568 380454 79888 380476
rect 79568 380218 79610 380454
rect 79846 380218 79888 380454
rect 79568 380134 79888 380218
rect 79568 379898 79610 380134
rect 79846 379898 79888 380134
rect 79568 379876 79888 379898
rect 64208 373254 64528 373276
rect 64208 373018 64250 373254
rect 64486 373018 64528 373254
rect 64208 372934 64528 373018
rect 64208 372698 64250 372934
rect 64486 372698 64528 372934
rect 64208 372676 64528 372698
rect 64208 369654 64528 369676
rect 64208 369418 64250 369654
rect 64486 369418 64528 369654
rect 64208 369334 64528 369418
rect 64208 369098 64250 369334
rect 64486 369098 64528 369334
rect 64208 369076 64528 369098
rect 64208 366054 64528 366076
rect 64208 365818 64250 366054
rect 64486 365818 64528 366054
rect 64208 365734 64528 365818
rect 64208 365498 64250 365734
rect 64486 365498 64528 365734
rect 64208 365476 64528 365498
rect 64208 362454 64528 362476
rect 64208 362218 64250 362454
rect 64486 362218 64528 362454
rect 64208 362134 64528 362218
rect 64208 361898 64250 362134
rect 64486 361898 64528 362134
rect 64208 361876 64528 361898
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 79568 355254 79888 355276
rect 79568 355018 79610 355254
rect 79846 355018 79888 355254
rect 79568 354934 79888 355018
rect 79568 354698 79610 354934
rect 79846 354698 79888 354934
rect 79568 354676 79888 354698
rect 79568 351654 79888 351676
rect 79568 351418 79610 351654
rect 79846 351418 79888 351654
rect 79568 351334 79888 351418
rect 79568 351098 79610 351334
rect 79846 351098 79888 351334
rect 79568 351076 79888 351098
rect 79568 348054 79888 348076
rect 79568 347818 79610 348054
rect 79846 347818 79888 348054
rect 79568 347734 79888 347818
rect 79568 347498 79610 347734
rect 79846 347498 79888 347734
rect 79568 347476 79888 347498
rect 79568 344454 79888 344476
rect 79568 344218 79610 344454
rect 79846 344218 79888 344454
rect 79568 344134 79888 344218
rect 79568 343898 79610 344134
rect 79846 343898 79888 344134
rect 79568 343876 79888 343898
rect 64208 337254 64528 337276
rect 64208 337018 64250 337254
rect 64486 337018 64528 337254
rect 64208 336934 64528 337018
rect 64208 336698 64250 336934
rect 64486 336698 64528 336934
rect 64208 336676 64528 336698
rect 64208 333654 64528 333676
rect 64208 333418 64250 333654
rect 64486 333418 64528 333654
rect 64208 333334 64528 333418
rect 64208 333098 64250 333334
rect 64486 333098 64528 333334
rect 64208 333076 64528 333098
rect 64208 330054 64528 330076
rect 64208 329818 64250 330054
rect 64486 329818 64528 330054
rect 64208 329734 64528 329818
rect 64208 329498 64250 329734
rect 64486 329498 64528 329734
rect 64208 329476 64528 329498
rect 64208 326454 64528 326476
rect 64208 326218 64250 326454
rect 64486 326218 64528 326454
rect 64208 326134 64528 326218
rect 64208 325898 64250 326134
rect 64486 325898 64528 326134
rect 64208 325876 64528 325898
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 79568 319254 79888 319276
rect 79568 319018 79610 319254
rect 79846 319018 79888 319254
rect 79568 318934 79888 319018
rect 79568 318698 79610 318934
rect 79846 318698 79888 318934
rect 79568 318676 79888 318698
rect 79568 315654 79888 315676
rect 79568 315418 79610 315654
rect 79846 315418 79888 315654
rect 79568 315334 79888 315418
rect 79568 315098 79610 315334
rect 79846 315098 79888 315334
rect 79568 315076 79888 315098
rect 79568 312054 79888 312076
rect 79568 311818 79610 312054
rect 79846 311818 79888 312054
rect 79568 311734 79888 311818
rect 79568 311498 79610 311734
rect 79846 311498 79888 311734
rect 79568 311476 79888 311498
rect 79568 308454 79888 308476
rect 79568 308218 79610 308454
rect 79846 308218 79888 308454
rect 79568 308134 79888 308218
rect 79568 307898 79610 308134
rect 79846 307898 79888 308134
rect 79568 307876 79888 307898
rect 61147 300660 61213 300661
rect 61147 300596 61148 300660
rect 61212 300596 61213 300660
rect 61147 300595 61213 300596
rect 61699 300660 61765 300661
rect 61699 300596 61700 300660
rect 61764 300596 61765 300660
rect 61699 300595 61765 300596
rect 61150 299573 61210 300595
rect 61147 299572 61213 299573
rect 61147 299508 61148 299572
rect 61212 299508 61213 299572
rect 61147 299507 61213 299508
rect 58404 276054 59004 297000
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 57835 29340 57901 29341
rect 57835 29276 57836 29340
rect 57900 29276 57901 29340
rect 57835 29275 57901 29276
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 279654 62604 297000
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 283254 66204 297000
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 72804 290454 73404 297000
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 67403 177308 67469 177309
rect 67403 177244 67404 177308
rect 67468 177244 67469 177308
rect 67403 177243 67469 177244
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 67406 164253 67466 177243
rect 67403 164252 67469 164253
rect 67403 164188 67404 164252
rect 67468 164188 67469 164252
rect 67403 164187 67469 164188
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 67403 126036 67469 126037
rect 67403 125972 67404 126036
rect 67468 125972 67469 126036
rect 67403 125971 67469 125972
rect 67406 125629 67466 125971
rect 67403 125628 67469 125629
rect 67403 125564 67404 125628
rect 67468 125564 67469 125628
rect 67403 125563 67469 125564
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 67587 76124 67653 76125
rect 67587 76060 67588 76124
rect 67652 76060 67653 76124
rect 67587 76059 67653 76060
rect 67590 75853 67650 76059
rect 67587 75852 67653 75853
rect 67587 75788 67588 75852
rect 67652 75788 67653 75852
rect 67587 75787 67653 75788
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 67587 40220 67653 40221
rect 67587 40156 67588 40220
rect 67652 40156 67653 40220
rect 67587 40155 67653 40156
rect 67590 39949 67650 40155
rect 67587 39948 67653 39949
rect 67587 39884 67588 39948
rect 67652 39884 67653 39948
rect 67587 39883 67653 39884
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 294054 77004 297000
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 261654 80604 297000
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 265254 84204 297000
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 90804 272454 91404 297000
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 86907 29612 86973 29613
rect 86907 29548 86908 29612
rect 86972 29548 86973 29612
rect 86907 29547 86973 29548
rect 86910 29205 86970 29547
rect 86907 29204 86973 29205
rect 86907 29140 86908 29204
rect 86972 29140 86973 29204
rect 86907 29139 86973 29140
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 276054 95004 297000
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 279654 98604 297000
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 283254 102204 297000
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 290454 109404 297000
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 294054 113004 297000
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 116004 261654 116604 297000
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 115795 76396 115861 76397
rect 115795 76332 115796 76396
rect 115860 76332 115861 76396
rect 115795 76331 115861 76332
rect 115798 75989 115858 76331
rect 115795 75988 115861 75989
rect 115795 75924 115796 75988
rect 115860 75924 115861 75988
rect 115795 75923 115861 75924
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 115795 40492 115861 40493
rect 115795 40428 115796 40492
rect 115860 40428 115861 40492
rect 115795 40427 115861 40428
rect 115798 40085 115858 40427
rect 115795 40084 115861 40085
rect 115795 40020 115796 40084
rect 115860 40020 115861 40084
rect 115795 40019 115861 40020
rect 115795 29476 115861 29477
rect 115795 29412 115796 29476
rect 115860 29412 115861 29476
rect 115795 29411 115861 29412
rect 115798 29069 115858 29411
rect 115795 29068 115861 29069
rect 115795 29004 115796 29068
rect 115860 29004 115861 29068
rect 115795 29003 115861 29004
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 265254 120204 297000
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 126804 272454 127404 297000
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 125547 76532 125613 76533
rect 125547 76468 125548 76532
rect 125612 76468 125613 76532
rect 125547 76467 125613 76468
rect 125550 76261 125610 76467
rect 125547 76260 125613 76261
rect 125547 76196 125548 76260
rect 125612 76196 125613 76260
rect 125547 76195 125613 76196
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 125547 40628 125613 40629
rect 125547 40564 125548 40628
rect 125612 40564 125613 40628
rect 125547 40563 125613 40564
rect 125550 40357 125610 40563
rect 125547 40356 125613 40357
rect 125547 40292 125548 40356
rect 125612 40292 125613 40356
rect 125547 40291 125613 40292
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 276054 131004 297000
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 134004 279654 134604 297000
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 133827 29476 133893 29477
rect 133827 29412 133828 29476
rect 133892 29412 133893 29476
rect 133827 29411 133893 29412
rect 133830 29205 133890 29411
rect 133827 29204 133893 29205
rect 133827 29140 133828 29204
rect 133892 29140 133893 29204
rect 133827 29139 133893 29140
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 283254 138204 297000
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 290454 145404 297000
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 294054 149004 297000
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 261654 152604 297000
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 265254 156204 297000
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 272454 163404 297000
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 276054 167004 297000
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 279654 170604 297000
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 283254 174204 297000
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 290454 181404 297000
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 294054 185004 297000
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 261654 188604 297000
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 265254 192204 297000
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 272454 199404 297000
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 276054 203004 297000
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 279654 206604 297000
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 283254 210204 297000
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 290454 217404 297000
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 294054 221004 297000
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 261654 224604 297000
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 265254 228204 297000
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 272454 235404 297000
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 276054 239004 297000
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 279654 242604 297000
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 283254 246204 297000
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 290454 253404 297000
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 294054 257004 297000
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 261654 260604 297000
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 265254 264204 297000
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 272454 271404 297000
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 276054 275004 297000
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 279654 278604 297000
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 283254 282204 297000
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299427 686220 299493 686221
rect 299427 686156 299428 686220
rect 299492 686156 299493 686220
rect 299427 686155 299493 686156
rect 299430 685949 299490 686155
rect 299427 685948 299493 685949
rect 299427 685884 299428 685948
rect 299492 685884 299493 685948
rect 299427 685883 299493 685884
rect 299427 673844 299493 673845
rect 299427 673780 299428 673844
rect 299492 673780 299493 673844
rect 299427 673779 299493 673780
rect 299430 673573 299490 673779
rect 299427 673572 299493 673573
rect 299427 673508 299428 673572
rect 299492 673508 299493 673572
rect 299427 673507 299493 673508
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 654247 307404 667898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 654247 311004 671498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 654247 314604 675098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 654247 318204 678698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 654247 325404 685898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654247 329004 689498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 654247 332604 657098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 654247 336204 660698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 654247 343404 667898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 654247 347004 671498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 654247 350604 675098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 357387 686356 357453 686357
rect 357387 686292 357388 686356
rect 357452 686292 357453 686356
rect 357387 686291 357453 686292
rect 357390 685949 357450 686291
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 357387 685948 357453 685949
rect 357387 685884 357388 685948
rect 357452 685884 357453 685948
rect 357387 685883 357453 685884
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 654247 354204 678698
rect 357387 673980 357453 673981
rect 357387 673916 357388 673980
rect 357452 673916 357453 673980
rect 357387 673915 357453 673916
rect 357390 673573 357450 673915
rect 357387 673572 357453 673573
rect 357387 673508 357388 673572
rect 357452 673508 357453 673572
rect 357387 673507 357453 673508
rect 360804 654247 361404 685898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654247 365004 689498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 654247 368604 657098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 376707 686492 376773 686493
rect 376707 686428 376708 686492
rect 376772 686428 376773 686492
rect 376707 686427 376773 686428
rect 376710 686221 376770 686427
rect 376707 686220 376773 686221
rect 376707 686156 376708 686220
rect 376772 686156 376773 686220
rect 376707 686155 376773 686156
rect 376707 674116 376773 674117
rect 376707 674052 376708 674116
rect 376772 674052 376773 674116
rect 376707 674051 376773 674052
rect 376710 673845 376770 674051
rect 376707 673844 376773 673845
rect 376707 673780 376708 673844
rect 376772 673780 376773 673844
rect 376707 673779 376773 673780
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 654247 372204 660698
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 654247 379404 667898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 654247 383004 671498
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 654247 386604 675098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 654247 390204 678698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 378547 652900 378613 652901
rect 378547 652836 378548 652900
rect 378612 652836 378613 652900
rect 378547 652835 378613 652836
rect 383515 652900 383581 652901
rect 383515 652836 383516 652900
rect 383580 652836 383581 652900
rect 383515 652835 383581 652836
rect 378550 651070 378610 652835
rect 383518 651130 383578 652835
rect 383518 651070 383603 651130
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 386938 643254 387262 643276
rect 386938 643018 386982 643254
rect 387218 643018 387262 643254
rect 386938 642934 387262 643018
rect 386938 642698 386982 642934
rect 387218 642698 387262 642934
rect 386938 642676 387262 642698
rect 386938 639654 387262 639676
rect 386938 639418 386982 639654
rect 387218 639418 387262 639654
rect 386938 639334 387262 639418
rect 386938 639098 386982 639334
rect 387218 639098 387262 639334
rect 386938 639076 387262 639098
rect 386938 636054 387262 636076
rect 386938 635818 386982 636054
rect 387218 635818 387262 636054
rect 386938 635734 387262 635818
rect 386938 635498 386982 635734
rect 387218 635498 387262 635734
rect 386938 635476 387262 635498
rect 386938 632454 387262 632476
rect 386938 632218 386982 632454
rect 387218 632218 387262 632454
rect 386938 632134 387262 632218
rect 386938 631898 386982 632134
rect 387218 631898 387262 632134
rect 386938 631876 387262 631898
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 386494 625254 386814 625276
rect 386494 625018 386536 625254
rect 386772 625018 386814 625254
rect 386494 624934 386814 625018
rect 386494 624698 386536 624934
rect 386772 624698 386814 624934
rect 386494 624676 386814 624698
rect 386494 621654 386814 621676
rect 386494 621418 386536 621654
rect 386772 621418 386814 621654
rect 386494 621334 386814 621418
rect 386494 621098 386536 621334
rect 386772 621098 386814 621334
rect 386494 621076 386814 621098
rect 386494 618054 386814 618076
rect 386494 617818 386536 618054
rect 386772 617818 386814 618054
rect 386494 617734 386814 617818
rect 386494 617498 386536 617734
rect 386772 617498 386814 617734
rect 386494 617476 386814 617498
rect 386494 614454 386814 614476
rect 386494 614218 386536 614454
rect 386772 614218 386814 614454
rect 386494 614134 386814 614218
rect 386494 613898 386536 614134
rect 386772 613898 386814 614134
rect 386494 613876 386814 613898
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 386938 607254 387262 607276
rect 386938 607018 386982 607254
rect 387218 607018 387262 607254
rect 386938 606934 387262 607018
rect 386938 606698 386982 606934
rect 387218 606698 387262 606934
rect 386938 606676 387262 606698
rect 386938 603654 387262 603676
rect 386938 603418 386982 603654
rect 387218 603418 387262 603654
rect 386938 603334 387262 603418
rect 386938 603098 386982 603334
rect 387218 603098 387262 603334
rect 386938 603076 387262 603098
rect 386938 600054 387262 600076
rect 386938 599818 386982 600054
rect 387218 599818 387262 600054
rect 386938 599734 387262 599818
rect 386938 599498 386982 599734
rect 387218 599498 387262 599734
rect 386938 599476 387262 599498
rect 386938 596454 387262 596476
rect 386938 596218 386982 596454
rect 387218 596218 387262 596454
rect 386938 596134 387262 596218
rect 386938 595898 386982 596134
rect 387218 595898 387262 596134
rect 386938 595876 387262 595898
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 386494 589254 386814 589276
rect 386494 589018 386536 589254
rect 386772 589018 386814 589254
rect 386494 588934 386814 589018
rect 386494 588698 386536 588934
rect 386772 588698 386814 588934
rect 386494 588676 386814 588698
rect 386494 585654 386814 585676
rect 386494 585418 386536 585654
rect 386772 585418 386814 585654
rect 386494 585334 386814 585418
rect 386494 585098 386536 585334
rect 386772 585098 386814 585334
rect 386494 585076 386814 585098
rect 386494 582054 386814 582076
rect 386494 581818 386536 582054
rect 386772 581818 386814 582054
rect 386494 581734 386814 581818
rect 386494 581498 386536 581734
rect 386772 581498 386814 581734
rect 386494 581476 386814 581498
rect 386494 578454 386814 578476
rect 386494 578218 386536 578454
rect 386772 578218 386814 578454
rect 386494 578134 386814 578218
rect 386494 577898 386536 578134
rect 386772 577898 386814 578134
rect 386494 577876 386814 577898
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 386938 571254 387262 571276
rect 386938 571018 386982 571254
rect 387218 571018 387262 571254
rect 386938 570934 387262 571018
rect 386938 570698 386982 570934
rect 387218 570698 387262 570934
rect 386938 570676 387262 570698
rect 386938 567654 387262 567676
rect 386938 567418 386982 567654
rect 387218 567418 387262 567654
rect 386938 567334 387262 567418
rect 386938 567098 386982 567334
rect 387218 567098 387262 567334
rect 386938 567076 387262 567098
rect 386938 564054 387262 564076
rect 386938 563818 386982 564054
rect 387218 563818 387262 564054
rect 386938 563734 387262 563818
rect 386938 563498 386982 563734
rect 387218 563498 387262 563734
rect 386938 563476 387262 563498
rect 323534 560430 323840 560490
rect 327030 560430 327344 560490
rect 328636 560430 328930 560490
rect 313782 558925 313842 560350
rect 316174 560290 316832 560350
rect 317462 560290 318000 560350
rect 318934 560290 319168 560350
rect 316174 558925 316234 560290
rect 313779 558924 313845 558925
rect 313779 558860 313780 558924
rect 313844 558860 313845 558924
rect 313779 558859 313845 558860
rect 316171 558924 316237 558925
rect 316171 558860 316172 558924
rect 316236 558860 316237 558924
rect 316171 558859 316237 558860
rect 317462 558517 317522 560290
rect 318934 558925 318994 560290
rect 320306 560010 320366 560320
rect 320222 559950 320366 560010
rect 320958 560290 321504 560350
rect 322430 560290 322672 560350
rect 322796 560290 322858 560350
rect 318931 558924 318997 558925
rect 318931 558860 318932 558924
rect 318996 558860 318997 558924
rect 318931 558859 318997 558860
rect 317459 558516 317525 558517
rect 317459 558452 317460 558516
rect 317524 558452 317525 558516
rect 317459 558451 317525 558452
rect 320222 557837 320282 559950
rect 320958 558925 321018 560290
rect 320955 558924 321021 558925
rect 320955 558860 320956 558924
rect 321020 558860 321021 558924
rect 320955 558859 321021 558860
rect 322430 558789 322490 560290
rect 322798 558925 322858 560290
rect 322795 558924 322861 558925
rect 322795 558860 322796 558924
rect 322860 558860 322861 558924
rect 322795 558859 322861 558860
rect 322427 558788 322493 558789
rect 322427 558724 322428 558788
rect 322492 558724 322493 558788
rect 322427 558723 322493 558724
rect 323534 558653 323594 560430
rect 323964 560290 324146 560350
rect 323531 558652 323597 558653
rect 323531 558588 323532 558652
rect 323596 558588 323597 558652
rect 323531 558587 323597 558588
rect 324086 557973 324146 560290
rect 324822 560290 325008 560350
rect 324822 558653 324882 560290
rect 325102 560010 325162 560320
rect 326110 560290 326176 560350
rect 325102 559950 325250 560010
rect 325190 558925 325250 559950
rect 325187 558924 325253 558925
rect 325187 558860 325188 558924
rect 325252 558860 325253 558924
rect 325187 558859 325253 558860
rect 326110 558653 326170 560290
rect 326294 558925 326354 560350
rect 326291 558924 326357 558925
rect 326291 558860 326292 558924
rect 326356 558860 326357 558924
rect 326291 558859 326357 558860
rect 327030 558789 327090 560430
rect 327468 560290 327642 560350
rect 327582 558925 327642 560290
rect 328482 559330 328542 560320
rect 328482 559270 328562 559330
rect 327579 558924 327645 558925
rect 327579 558860 327580 558924
rect 327644 558860 327645 558924
rect 327579 558859 327645 558860
rect 328502 558789 328562 559270
rect 327027 558788 327093 558789
rect 327027 558724 327028 558788
rect 327092 558724 327093 558788
rect 327027 558723 327093 558724
rect 328499 558788 328565 558789
rect 328499 558724 328500 558788
rect 328564 558724 328565 558788
rect 328499 558723 328565 558724
rect 324819 558652 324885 558653
rect 324819 558588 324820 558652
rect 324884 558588 324885 558652
rect 324819 558587 324885 558588
rect 326107 558652 326173 558653
rect 326107 558588 326108 558652
rect 326172 558588 326173 558652
rect 326107 558587 326173 558588
rect 328870 558245 328930 560430
rect 330526 560430 330848 560490
rect 332140 560430 332426 560490
rect 329606 560290 329680 560350
rect 329606 558653 329666 560290
rect 329603 558652 329669 558653
rect 329603 558588 329604 558652
rect 329668 558588 329669 558652
rect 329603 558587 329669 558588
rect 329790 558381 329850 560350
rect 330526 558653 330586 560430
rect 330972 560290 331138 560350
rect 331078 558925 331138 560290
rect 331814 560290 332016 560350
rect 331814 558925 331874 560290
rect 331075 558924 331141 558925
rect 331075 558860 331076 558924
rect 331140 558860 331141 558924
rect 331075 558859 331141 558860
rect 331811 558924 331877 558925
rect 331811 558860 331812 558924
rect 331876 558860 331877 558924
rect 331811 558859 331877 558860
rect 330523 558652 330589 558653
rect 330523 558588 330524 558652
rect 330588 558588 330589 558652
rect 330523 558587 330589 558588
rect 329787 558380 329853 558381
rect 329787 558316 329788 558380
rect 329852 558316 329853 558380
rect 329787 558315 329853 558316
rect 332366 558245 332426 560430
rect 334022 560430 334352 560490
rect 335644 560430 335922 560490
rect 332734 560290 333184 560350
rect 332734 558789 332794 560290
rect 333286 558925 333346 560350
rect 333283 558924 333349 558925
rect 333283 558860 333284 558924
rect 333348 558860 333349 558924
rect 333283 558859 333349 558860
rect 334022 558789 334082 560430
rect 334476 560290 334634 560350
rect 334574 558925 334634 560290
rect 335490 560010 335550 560320
rect 335490 559950 335554 560010
rect 334571 558924 334637 558925
rect 334571 558860 334572 558924
rect 334636 558860 334637 558924
rect 334571 558859 334637 558860
rect 335494 558789 335554 559950
rect 335862 558925 335922 560430
rect 339910 560430 340192 560490
rect 341484 560430 341810 560490
rect 336598 560290 336688 560350
rect 335859 558924 335925 558925
rect 335859 558860 335860 558924
rect 335924 558860 335925 558924
rect 335859 558859 335925 558860
rect 336598 558789 336658 560290
rect 336782 558925 336842 560320
rect 337702 560290 337856 560350
rect 337702 558925 337762 560290
rect 337950 559330 338010 560320
rect 337886 559270 338010 559330
rect 336779 558924 336845 558925
rect 336779 558860 336780 558924
rect 336844 558860 336845 558924
rect 336779 558859 336845 558860
rect 337699 558924 337765 558925
rect 337699 558860 337700 558924
rect 337764 558860 337765 558924
rect 337699 558859 337765 558860
rect 332731 558788 332797 558789
rect 332731 558724 332732 558788
rect 332796 558724 332797 558788
rect 332731 558723 332797 558724
rect 334019 558788 334085 558789
rect 334019 558724 334020 558788
rect 334084 558724 334085 558788
rect 334019 558723 334085 558724
rect 335491 558788 335557 558789
rect 335491 558724 335492 558788
rect 335556 558724 335557 558788
rect 335491 558723 335557 558724
rect 336595 558788 336661 558789
rect 336595 558724 336596 558788
rect 336660 558724 336661 558788
rect 336595 558723 336661 558724
rect 337886 558517 337946 559270
rect 338990 558789 339050 560350
rect 339148 560290 339234 560350
rect 339174 558925 339234 560290
rect 339171 558924 339237 558925
rect 339171 558860 339172 558924
rect 339236 558860 339237 558924
rect 339171 558859 339237 558860
rect 339910 558789 339970 560430
rect 340316 560290 340522 560350
rect 340462 558925 340522 560290
rect 341014 560290 341360 560350
rect 340459 558924 340525 558925
rect 340459 558860 340460 558924
rect 340524 558860 340525 558924
rect 340459 558859 340525 558860
rect 341014 558789 341074 560290
rect 341750 558925 341810 560430
rect 346902 560430 347200 560490
rect 348492 560430 348802 560490
rect 351996 560430 352298 560490
rect 359004 560430 359290 560490
rect 341747 558924 341813 558925
rect 341747 558860 341748 558924
rect 341812 558860 341813 558924
rect 341747 558859 341813 558860
rect 342486 558789 342546 560350
rect 342652 560290 342730 560350
rect 342670 558925 342730 560290
rect 343666 560010 343726 560320
rect 343820 560290 344018 560350
rect 343590 559950 343726 560010
rect 342667 558924 342733 558925
rect 342667 558860 342668 558924
rect 342732 558860 342733 558924
rect 342667 558859 342733 558860
rect 343590 558789 343650 559950
rect 343958 558925 344018 560290
rect 344326 560290 344864 560350
rect 344326 558925 344386 560290
rect 344958 559330 345018 560320
rect 344878 559270 345018 559330
rect 343955 558924 344021 558925
rect 343955 558860 343956 558924
rect 344020 558860 344021 558924
rect 343955 558859 344021 558860
rect 344323 558924 344389 558925
rect 344323 558860 344324 558924
rect 344388 558860 344389 558924
rect 344323 558859 344389 558860
rect 338987 558788 339053 558789
rect 338987 558724 338988 558788
rect 339052 558724 339053 558788
rect 338987 558723 339053 558724
rect 339907 558788 339973 558789
rect 339907 558724 339908 558788
rect 339972 558724 339973 558788
rect 339907 558723 339973 558724
rect 341011 558788 341077 558789
rect 341011 558724 341012 558788
rect 341076 558724 341077 558788
rect 341011 558723 341077 558724
rect 342483 558788 342549 558789
rect 342483 558724 342484 558788
rect 342548 558724 342549 558788
rect 342483 558723 342549 558724
rect 343587 558788 343653 558789
rect 343587 558724 343588 558788
rect 343652 558724 343653 558788
rect 343587 558723 343653 558724
rect 337883 558516 337949 558517
rect 337883 558452 337884 558516
rect 337948 558452 337949 558516
rect 337883 558451 337949 558452
rect 328867 558244 328933 558245
rect 328867 558180 328868 558244
rect 328932 558180 328933 558244
rect 328867 558179 328933 558180
rect 332363 558244 332429 558245
rect 332363 558180 332364 558244
rect 332428 558180 332429 558244
rect 332363 558179 332429 558180
rect 324083 557972 324149 557973
rect 324083 557908 324084 557972
rect 324148 557908 324149 557972
rect 324083 557907 324149 557908
rect 320219 557836 320285 557837
rect 320219 557772 320220 557836
rect 320284 557772 320285 557836
rect 320219 557771 320285 557772
rect 344878 557701 344938 559270
rect 345982 558789 346042 560350
rect 346156 560290 346226 560350
rect 346166 558925 346226 560290
rect 346163 558924 346229 558925
rect 346163 558860 346164 558924
rect 346228 558860 346229 558924
rect 346163 558859 346229 558860
rect 346902 558789 346962 560430
rect 347324 560290 347514 560350
rect 347454 558925 347514 560290
rect 348190 560290 348368 560350
rect 347451 558924 347517 558925
rect 347451 558860 347452 558924
rect 347516 558860 347517 558924
rect 347451 558859 347517 558860
rect 348190 558789 348250 560290
rect 348742 558925 348802 560430
rect 348739 558924 348805 558925
rect 348739 558860 348740 558924
rect 348804 558860 348805 558924
rect 348739 558859 348805 558860
rect 349478 558789 349538 560350
rect 349660 560290 349722 560350
rect 349662 558925 349722 560290
rect 350674 560010 350734 560320
rect 350828 560290 351010 560350
rect 350582 559950 350734 560010
rect 349659 558924 349725 558925
rect 349659 558860 349660 558924
rect 349724 558860 349725 558924
rect 349659 558859 349725 558860
rect 345979 558788 346045 558789
rect 345979 558724 345980 558788
rect 346044 558724 346045 558788
rect 345979 558723 346045 558724
rect 346899 558788 346965 558789
rect 346899 558724 346900 558788
rect 346964 558724 346965 558788
rect 346899 558723 346965 558724
rect 348187 558788 348253 558789
rect 348187 558724 348188 558788
rect 348252 558724 348253 558788
rect 348187 558723 348253 558724
rect 349475 558788 349541 558789
rect 349475 558724 349476 558788
rect 349540 558724 349541 558788
rect 349475 558723 349541 558724
rect 350582 558517 350642 559950
rect 350579 558516 350645 558517
rect 350579 558452 350580 558516
rect 350644 558452 350645 558516
rect 350579 558451 350645 558452
rect 344875 557700 344941 557701
rect 344875 557636 344876 557700
rect 344940 557636 344941 557700
rect 344875 557635 344941 557636
rect 350950 557565 351010 560290
rect 351842 559333 351902 560320
rect 351842 559332 351933 559333
rect 351842 559270 351868 559332
rect 351867 559268 351868 559270
rect 351932 559268 351933 559332
rect 351867 559267 351933 559268
rect 350947 557564 351013 557565
rect 350947 557500 350948 557564
rect 351012 557500 351013 557564
rect 350947 557499 351013 557500
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 524454 307404 557000
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 528054 311004 557000
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 531654 314604 557000
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 535254 318204 557000
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 542454 325404 557000
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 546054 329004 557000
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 549654 332604 557000
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 553254 336204 557000
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 524454 343404 557000
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 528054 347004 557000
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 531654 350604 557000
rect 352238 555525 352298 560430
rect 352422 560290 353040 560350
rect 352422 558925 352482 560290
rect 352419 558924 352485 558925
rect 352419 558860 352420 558924
rect 352484 558860 352485 558924
rect 352419 558859 352485 558860
rect 353158 557701 353218 560350
rect 353526 560290 354208 560350
rect 354332 560290 354506 560350
rect 353526 558789 353586 560290
rect 353523 558788 353589 558789
rect 353523 558724 353524 558788
rect 353588 558724 353589 558788
rect 353523 558723 353589 558724
rect 353155 557700 353221 557701
rect 353155 557636 353156 557700
rect 353220 557636 353221 557700
rect 353155 557635 353221 557636
rect 354446 557565 354506 560290
rect 354814 560290 355376 560350
rect 354814 558381 354874 560290
rect 355470 560010 355530 560320
rect 356102 560290 356544 560350
rect 355470 559950 355610 560010
rect 354811 558380 354877 558381
rect 354811 558316 354812 558380
rect 354876 558316 354877 558380
rect 354811 558315 354877 558316
rect 355550 557565 355610 559950
rect 356102 558653 356162 560290
rect 356099 558652 356165 558653
rect 356099 558588 356100 558652
rect 356164 558588 356165 558652
rect 356099 558587 356165 558588
rect 356654 557565 356714 560350
rect 357682 560010 357742 560320
rect 357836 560290 358002 560350
rect 357574 559950 357742 560010
rect 357574 558789 357634 559950
rect 357571 558788 357637 558789
rect 357571 558724 357572 558788
rect 357636 558724 357637 558788
rect 357571 558723 357637 558724
rect 357942 557565 358002 560290
rect 358850 559333 358910 560320
rect 358850 559332 358925 559333
rect 358850 559270 358860 559332
rect 358859 559268 358860 559270
rect 358924 559268 358925 559332
rect 358859 559267 358925 559268
rect 354443 557564 354509 557565
rect 354443 557500 354444 557564
rect 354508 557500 354509 557564
rect 354443 557499 354509 557500
rect 355547 557564 355613 557565
rect 355547 557500 355548 557564
rect 355612 557500 355613 557564
rect 355547 557499 355613 557500
rect 356651 557564 356717 557565
rect 356651 557500 356652 557564
rect 356716 557500 356717 557564
rect 356651 557499 356717 557500
rect 357939 557564 358005 557565
rect 357939 557500 357940 557564
rect 358004 557500 358005 557564
rect 357939 557499 358005 557500
rect 352235 555524 352301 555525
rect 352235 555460 352236 555524
rect 352300 555460 352301 555524
rect 352235 555459 352301 555460
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 535254 354204 557000
rect 359230 555525 359290 560430
rect 359227 555524 359293 555525
rect 359227 555460 359228 555524
rect 359292 555460 359293 555524
rect 359227 555459 359293 555460
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 542454 361404 557000
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 546054 365004 557000
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 549654 368604 557000
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 553254 372204 557000
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 524454 379404 557000
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 528054 383004 557000
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 531654 386604 557000
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 535254 390204 557000
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 434667 686492 434733 686493
rect 434667 686428 434668 686492
rect 434732 686428 434733 686492
rect 434667 686427 434733 686428
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 434670 686085 434730 686427
rect 434667 686084 434733 686085
rect 434667 686020 434668 686084
rect 434732 686020 434733 686084
rect 434667 686019 434733 686020
rect 432804 650454 433404 685898
rect 436404 654247 437004 689498
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 654247 440604 657098
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 654247 444204 660698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 654247 451404 667898
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 654247 455004 671498
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 654247 458604 675098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 654247 462204 678698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 654247 469404 685898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654247 473004 689498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 654247 476604 657098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 654247 480204 660698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 654247 487404 667898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 654247 491004 671498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 654247 494604 675098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 654247 498204 678698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 654247 505404 685898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654247 509004 689498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 654247 512604 657098
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 654247 516204 660698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 507899 652900 507965 652901
rect 507899 652836 507900 652900
rect 507964 652836 507965 652900
rect 507899 652835 507965 652836
rect 513419 652900 513485 652901
rect 513419 652836 513420 652900
rect 513484 652836 513485 652900
rect 513419 652835 513485 652836
rect 507902 651130 507962 652835
rect 513422 651130 513482 652835
rect 507902 651070 508608 651130
rect 513422 651070 513603 651130
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 516938 643254 517262 643276
rect 516938 643018 516982 643254
rect 517218 643018 517262 643254
rect 516938 642934 517262 643018
rect 516938 642698 516982 642934
rect 517218 642698 517262 642934
rect 516938 642676 517262 642698
rect 516938 639654 517262 639676
rect 516938 639418 516982 639654
rect 517218 639418 517262 639654
rect 516938 639334 517262 639418
rect 516938 639098 516982 639334
rect 517218 639098 517262 639334
rect 516938 639076 517262 639098
rect 516938 636054 517262 636076
rect 516938 635818 516982 636054
rect 517218 635818 517262 636054
rect 516938 635734 517262 635818
rect 516938 635498 516982 635734
rect 517218 635498 517262 635734
rect 516938 635476 517262 635498
rect 516938 632454 517262 632476
rect 516938 632218 516982 632454
rect 517218 632218 517262 632454
rect 516938 632134 517262 632218
rect 516938 631898 516982 632134
rect 517218 631898 517262 632134
rect 516938 631876 517262 631898
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 516494 625254 516814 625276
rect 516494 625018 516536 625254
rect 516772 625018 516814 625254
rect 516494 624934 516814 625018
rect 516494 624698 516536 624934
rect 516772 624698 516814 624934
rect 516494 624676 516814 624698
rect 516494 621654 516814 621676
rect 516494 621418 516536 621654
rect 516772 621418 516814 621654
rect 516494 621334 516814 621418
rect 516494 621098 516536 621334
rect 516772 621098 516814 621334
rect 516494 621076 516814 621098
rect 516494 618054 516814 618076
rect 516494 617818 516536 618054
rect 516772 617818 516814 618054
rect 516494 617734 516814 617818
rect 516494 617498 516536 617734
rect 516772 617498 516814 617734
rect 516494 617476 516814 617498
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 516494 614454 516814 614476
rect 516494 614218 516536 614454
rect 516772 614218 516814 614454
rect 516494 614134 516814 614218
rect 516494 613898 516536 614134
rect 516772 613898 516814 614134
rect 516494 613876 516814 613898
rect 516938 607254 517262 607276
rect 516938 607018 516982 607254
rect 517218 607018 517262 607254
rect 516938 606934 517262 607018
rect 516938 606698 516982 606934
rect 517218 606698 517262 606934
rect 516938 606676 517262 606698
rect 516938 603654 517262 603676
rect 516938 603418 516982 603654
rect 517218 603418 517262 603654
rect 516938 603334 517262 603418
rect 516938 603098 516982 603334
rect 517218 603098 517262 603334
rect 516938 603076 517262 603098
rect 516938 600054 517262 600076
rect 516938 599818 516982 600054
rect 517218 599818 517262 600054
rect 516938 599734 517262 599818
rect 516938 599498 516982 599734
rect 517218 599498 517262 599734
rect 516938 599476 517262 599498
rect 516938 596454 517262 596476
rect 516938 596218 516982 596454
rect 517218 596218 517262 596454
rect 516938 596134 517262 596218
rect 516938 595898 516982 596134
rect 517218 595898 517262 596134
rect 516938 595876 517262 595898
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 516494 589254 516814 589276
rect 516494 589018 516536 589254
rect 516772 589018 516814 589254
rect 516494 588934 516814 589018
rect 516494 588698 516536 588934
rect 516772 588698 516814 588934
rect 516494 588676 516814 588698
rect 516494 585654 516814 585676
rect 516494 585418 516536 585654
rect 516772 585418 516814 585654
rect 516494 585334 516814 585418
rect 516494 585098 516536 585334
rect 516772 585098 516814 585334
rect 516494 585076 516814 585098
rect 516494 582054 516814 582076
rect 516494 581818 516536 582054
rect 516772 581818 516814 582054
rect 516494 581734 516814 581818
rect 516494 581498 516536 581734
rect 516772 581498 516814 581734
rect 516494 581476 516814 581498
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 516494 578454 516814 578476
rect 516494 578218 516536 578454
rect 516772 578218 516814 578454
rect 516494 578134 516814 578218
rect 516494 577898 516536 578134
rect 516772 577898 516814 578134
rect 516494 577876 516814 577898
rect 516938 571254 517262 571276
rect 516938 571018 516982 571254
rect 517218 571018 517262 571254
rect 516938 570934 517262 571018
rect 516938 570698 516982 570934
rect 517218 570698 517262 570934
rect 516938 570676 517262 570698
rect 516938 567654 517262 567676
rect 516938 567418 516982 567654
rect 517218 567418 517262 567654
rect 516938 567334 517262 567418
rect 516938 567098 516982 567334
rect 517218 567098 517262 567334
rect 516938 567076 517262 567098
rect 516938 564054 517262 564076
rect 516938 563818 516982 564054
rect 517218 563818 517262 564054
rect 516938 563734 517262 563818
rect 516938 563498 516982 563734
rect 517218 563498 517262 563734
rect 516938 563476 517262 563498
rect 454726 560430 455008 560490
rect 456300 560430 456626 560490
rect 443134 560290 443833 560350
rect 446262 560290 446832 560350
rect 447366 560290 448000 560350
rect 448470 560290 449168 560350
rect 449942 560290 450336 560350
rect 451414 560290 451504 560350
rect 443134 558925 443194 560290
rect 446262 558925 446322 560290
rect 447366 558925 447426 560290
rect 448470 558925 448530 560290
rect 449942 558925 450002 560290
rect 443131 558924 443197 558925
rect 443131 558860 443132 558924
rect 443196 558860 443197 558924
rect 443131 558859 443197 558860
rect 446259 558924 446325 558925
rect 446259 558860 446260 558924
rect 446324 558860 446325 558924
rect 446259 558859 446325 558860
rect 447363 558924 447429 558925
rect 447363 558860 447364 558924
rect 447428 558860 447429 558924
rect 447363 558859 447429 558860
rect 448467 558924 448533 558925
rect 448467 558860 448468 558924
rect 448532 558860 448533 558924
rect 448467 558859 448533 558860
rect 449939 558924 450005 558925
rect 449939 558860 449940 558924
rect 450004 558860 450005 558924
rect 449939 558859 450005 558860
rect 451414 557701 451474 560290
rect 452642 559330 452702 560320
rect 452796 560290 452946 560350
rect 452642 559270 452762 559330
rect 452702 558789 452762 559270
rect 452886 558925 452946 560290
rect 453622 560290 453840 560350
rect 453622 558925 453682 560290
rect 453934 559330 453994 560320
rect 453806 559270 453994 559330
rect 452883 558924 452949 558925
rect 452883 558860 452884 558924
rect 452948 558860 452949 558924
rect 452883 558859 452949 558860
rect 453619 558924 453685 558925
rect 453619 558860 453620 558924
rect 453684 558860 453685 558924
rect 453619 558859 453685 558860
rect 452699 558788 452765 558789
rect 452699 558724 452700 558788
rect 452764 558724 452765 558788
rect 452699 558723 452765 558724
rect 453806 558245 453866 559270
rect 454726 558925 454786 560430
rect 455132 560290 455338 560350
rect 454723 558924 454789 558925
rect 454723 558860 454724 558924
rect 454788 558860 454789 558924
rect 454723 558859 454789 558860
rect 455278 558381 455338 560290
rect 456014 560290 456176 560350
rect 456014 558653 456074 560290
rect 456011 558652 456077 558653
rect 456011 558588 456012 558652
rect 456076 558588 456077 558652
rect 456011 558587 456077 558588
rect 456566 558517 456626 560430
rect 461718 560430 462016 560490
rect 465214 560430 465520 560490
rect 472206 560430 472528 560490
rect 473820 560430 474106 560490
rect 457302 558653 457362 560350
rect 457468 560290 457546 560350
rect 457299 558652 457365 558653
rect 457299 558588 457300 558652
rect 457364 558588 457365 558652
rect 457299 558587 457365 558588
rect 456563 558516 456629 558517
rect 456563 558452 456564 558516
rect 456628 558452 456629 558516
rect 456563 558451 456629 558452
rect 457486 558381 457546 560290
rect 458482 560010 458542 560320
rect 458636 560290 458834 560350
rect 458406 559950 458542 560010
rect 458406 558925 458466 559950
rect 458403 558924 458469 558925
rect 458403 558860 458404 558924
rect 458468 558860 458469 558924
rect 458403 558859 458469 558860
rect 458774 558381 458834 560290
rect 459510 560290 459680 560350
rect 459510 558789 459570 560290
rect 459774 560010 459834 560320
rect 459774 559950 459938 560010
rect 459507 558788 459573 558789
rect 459507 558724 459508 558788
rect 459572 558724 459573 558788
rect 459507 558723 459573 558724
rect 455275 558380 455341 558381
rect 455275 558316 455276 558380
rect 455340 558316 455341 558380
rect 455275 558315 455341 558316
rect 457483 558380 457549 558381
rect 457483 558316 457484 558380
rect 457548 558316 457549 558380
rect 457483 558315 457549 558316
rect 458771 558380 458837 558381
rect 458771 558316 458772 558380
rect 458836 558316 458837 558380
rect 458771 558315 458837 558316
rect 459878 558245 459938 559950
rect 460798 558653 460858 560350
rect 460972 560290 461042 560350
rect 460982 558925 461042 560290
rect 461718 558925 461778 560430
rect 462110 559330 462170 560320
rect 462086 559270 462170 559330
rect 463006 560290 463184 560350
rect 460979 558924 461045 558925
rect 460979 558860 460980 558924
rect 461044 558860 461045 558924
rect 460979 558859 461045 558860
rect 461715 558924 461781 558925
rect 461715 558860 461716 558924
rect 461780 558860 461781 558924
rect 461715 558859 461781 558860
rect 462086 558789 462146 559270
rect 463006 558789 463066 560290
rect 463278 560010 463338 560320
rect 463278 559950 463434 560010
rect 463374 558925 463434 559950
rect 463371 558924 463437 558925
rect 463371 558860 463372 558924
rect 463436 558860 463437 558924
rect 463371 558859 463437 558860
rect 464294 558789 464354 560350
rect 464476 560290 464538 560350
rect 464478 558925 464538 560290
rect 464475 558924 464541 558925
rect 464475 558860 464476 558924
rect 464540 558860 464541 558924
rect 464475 558859 464541 558860
rect 465214 558789 465274 560430
rect 465644 560290 465826 560350
rect 465766 558925 465826 560290
rect 466502 560290 466688 560350
rect 465763 558924 465829 558925
rect 465763 558860 465764 558924
rect 465828 558860 465829 558924
rect 465763 558859 465829 558860
rect 462083 558788 462149 558789
rect 462083 558724 462084 558788
rect 462148 558724 462149 558788
rect 462083 558723 462149 558724
rect 463003 558788 463069 558789
rect 463003 558724 463004 558788
rect 463068 558724 463069 558788
rect 463003 558723 463069 558724
rect 464291 558788 464357 558789
rect 464291 558724 464292 558788
rect 464356 558724 464357 558788
rect 464291 558723 464357 558724
rect 465211 558788 465277 558789
rect 465211 558724 465212 558788
rect 465276 558724 465277 558788
rect 465211 558723 465277 558724
rect 466502 558653 466562 560290
rect 466782 560010 466842 560320
rect 467790 560290 467856 560350
rect 466782 559950 466930 560010
rect 466870 558925 466930 559950
rect 466867 558924 466933 558925
rect 466867 558860 466868 558924
rect 466932 558860 466933 558924
rect 466867 558859 466933 558860
rect 467790 558653 467850 560290
rect 467974 558925 468034 560350
rect 468710 560290 469024 560350
rect 468710 558925 468770 560290
rect 469118 559330 469178 560320
rect 469078 559270 469178 559330
rect 469998 560290 470192 560350
rect 467971 558924 468037 558925
rect 467971 558860 467972 558924
rect 468036 558860 468037 558924
rect 467971 558859 468037 558860
rect 468707 558924 468773 558925
rect 468707 558860 468708 558924
rect 468772 558860 468773 558924
rect 468707 558859 468773 558860
rect 469078 558789 469138 559270
rect 469998 558789 470058 560290
rect 470286 560010 470346 560320
rect 471286 560290 471360 560350
rect 470286 559950 470426 560010
rect 470366 558925 470426 559950
rect 470363 558924 470429 558925
rect 470363 558860 470364 558924
rect 470428 558860 470429 558924
rect 470363 558859 470429 558860
rect 471286 558789 471346 560290
rect 471470 558925 471530 560350
rect 471467 558924 471533 558925
rect 471467 558860 471468 558924
rect 471532 558860 471533 558924
rect 471467 558859 471533 558860
rect 472206 558789 472266 560430
rect 472652 560290 472818 560350
rect 472758 558925 472818 560290
rect 473494 560290 473696 560350
rect 472755 558924 472821 558925
rect 472755 558860 472756 558924
rect 472820 558860 472821 558924
rect 472755 558859 472821 558860
rect 473494 558789 473554 560290
rect 474046 558925 474106 560430
rect 481590 560430 481872 560490
rect 483164 560430 483490 560490
rect 486668 560430 486986 560490
rect 474782 560290 474864 560350
rect 474043 558924 474109 558925
rect 474043 558860 474044 558924
rect 474108 558860 474109 558924
rect 474043 558859 474109 558860
rect 474782 558789 474842 560290
rect 474966 558925 475026 560350
rect 475518 560290 476032 560350
rect 476156 560290 476314 560350
rect 474963 558924 475029 558925
rect 474963 558860 474964 558924
rect 475028 558860 475029 558924
rect 474963 558859 475029 558860
rect 475518 558789 475578 560290
rect 476254 558925 476314 560290
rect 477170 560010 477230 560320
rect 477294 560010 477354 560320
rect 478278 560290 478368 560350
rect 477170 559950 477234 560010
rect 477294 559950 477418 560010
rect 477174 558925 477234 559950
rect 476251 558924 476317 558925
rect 476251 558860 476252 558924
rect 476316 558860 476317 558924
rect 476251 558859 476317 558860
rect 477171 558924 477237 558925
rect 477171 558860 477172 558924
rect 477236 558860 477237 558924
rect 477171 558859 477237 558860
rect 469075 558788 469141 558789
rect 469075 558724 469076 558788
rect 469140 558724 469141 558788
rect 469075 558723 469141 558724
rect 469995 558788 470061 558789
rect 469995 558724 469996 558788
rect 470060 558724 470061 558788
rect 469995 558723 470061 558724
rect 471283 558788 471349 558789
rect 471283 558724 471284 558788
rect 471348 558724 471349 558788
rect 471283 558723 471349 558724
rect 472203 558788 472269 558789
rect 472203 558724 472204 558788
rect 472268 558724 472269 558788
rect 472203 558723 472269 558724
rect 473491 558788 473557 558789
rect 473491 558724 473492 558788
rect 473556 558724 473557 558788
rect 473491 558723 473557 558724
rect 474779 558788 474845 558789
rect 474779 558724 474780 558788
rect 474844 558724 474845 558788
rect 474779 558723 474845 558724
rect 475515 558788 475581 558789
rect 475515 558724 475516 558788
rect 475580 558724 475581 558788
rect 475515 558723 475581 558724
rect 460795 558652 460861 558653
rect 460795 558588 460796 558652
rect 460860 558588 460861 558652
rect 460795 558587 460861 558588
rect 466499 558652 466565 558653
rect 466499 558588 466500 558652
rect 466564 558588 466565 558652
rect 466499 558587 466565 558588
rect 467787 558652 467853 558653
rect 467787 558588 467788 558652
rect 467852 558588 467853 558652
rect 467787 558587 467853 558588
rect 453803 558244 453869 558245
rect 453803 558180 453804 558244
rect 453868 558180 453869 558244
rect 453803 558179 453869 558180
rect 459875 558244 459941 558245
rect 459875 558180 459876 558244
rect 459940 558180 459941 558244
rect 459875 558179 459941 558180
rect 475518 557701 475578 558723
rect 477358 558109 477418 559950
rect 478278 558925 478338 560290
rect 478275 558924 478341 558925
rect 478275 558860 478276 558924
rect 478340 558860 478341 558924
rect 478275 558859 478341 558860
rect 478462 558109 478522 560320
rect 479382 560290 479536 560350
rect 479660 560290 479810 560350
rect 479382 558925 479442 560290
rect 479379 558924 479445 558925
rect 479379 558860 479380 558924
rect 479444 558860 479445 558924
rect 479379 558859 479445 558860
rect 477355 558108 477421 558109
rect 477355 558044 477356 558108
rect 477420 558044 477421 558108
rect 477355 558043 477421 558044
rect 478459 558108 478525 558109
rect 478459 558044 478460 558108
rect 478524 558044 478525 558108
rect 478459 558043 478525 558044
rect 479750 557973 479810 560290
rect 480486 560290 480704 560350
rect 480828 560290 480914 560350
rect 480486 558789 480546 560290
rect 480854 558925 480914 560290
rect 480851 558924 480917 558925
rect 480851 558860 480852 558924
rect 480916 558860 480917 558924
rect 480851 558859 480917 558860
rect 480483 558788 480549 558789
rect 480483 558724 480484 558788
rect 480548 558724 480549 558788
rect 480483 558723 480549 558724
rect 481590 558517 481650 560430
rect 481996 560290 482202 560350
rect 481587 558516 481653 558517
rect 481587 558452 481588 558516
rect 481652 558452 481653 558516
rect 481587 558451 481653 558452
rect 479747 557972 479813 557973
rect 479747 557908 479748 557972
rect 479812 557908 479813 557972
rect 479747 557907 479813 557908
rect 482142 557837 482202 560290
rect 483010 559330 483070 560320
rect 483010 559270 483122 559330
rect 483062 558653 483122 559270
rect 483430 558925 483490 560430
rect 483614 560290 484208 560350
rect 483427 558924 483493 558925
rect 483427 558860 483428 558924
rect 483492 558860 483493 558924
rect 483427 558859 483493 558860
rect 483059 558652 483125 558653
rect 483059 558588 483060 558652
rect 483124 558588 483125 558652
rect 483059 558587 483125 558588
rect 482139 557836 482205 557837
rect 482139 557772 482140 557836
rect 482204 557772 482205 557836
rect 482139 557771 482205 557772
rect 483614 557701 483674 560290
rect 484302 559330 484362 560320
rect 484166 559270 484362 559330
rect 484718 560290 485376 560350
rect 485500 560290 485698 560350
rect 484166 558245 484226 559270
rect 484718 558789 484778 560290
rect 485638 558925 485698 560290
rect 486006 560290 486544 560350
rect 486006 558925 486066 560290
rect 485635 558924 485701 558925
rect 485635 558860 485636 558924
rect 485700 558860 485701 558924
rect 485635 558859 485701 558860
rect 486003 558924 486069 558925
rect 486003 558860 486004 558924
rect 486068 558860 486069 558924
rect 486003 558859 486069 558860
rect 484715 558788 484781 558789
rect 484715 558724 484716 558788
rect 484780 558724 484781 558788
rect 484715 558723 484781 558724
rect 486926 558245 486986 560430
rect 522804 560454 523404 595898
rect 487294 560290 487712 560350
rect 487836 560290 487906 560350
rect 487294 558517 487354 560290
rect 487291 558516 487357 558517
rect 487291 558452 487292 558516
rect 487356 558452 487357 558516
rect 487291 558451 487357 558452
rect 487846 558245 487906 560290
rect 488582 560290 488880 560350
rect 489004 560290 489194 560350
rect 488582 558653 488642 560290
rect 488579 558652 488645 558653
rect 488579 558588 488580 558652
rect 488644 558588 488645 558652
rect 488579 558587 488645 558588
rect 489134 558381 489194 560290
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 489131 558380 489197 558381
rect 489131 558316 489132 558380
rect 489196 558316 489197 558380
rect 489131 558315 489197 558316
rect 484163 558244 484229 558245
rect 484163 558180 484164 558244
rect 484228 558180 484229 558244
rect 484163 558179 484229 558180
rect 486923 558244 486989 558245
rect 486923 558180 486924 558244
rect 486988 558180 486989 558244
rect 486923 558179 486989 558180
rect 487843 558244 487909 558245
rect 487843 558180 487844 558244
rect 487908 558180 487909 558244
rect 487843 558179 487909 558180
rect 451411 557700 451477 557701
rect 451411 557636 451412 557700
rect 451476 557636 451477 557700
rect 451411 557635 451477 557636
rect 475515 557700 475581 557701
rect 475515 557636 475516 557700
rect 475580 557636 475581 557700
rect 475515 557635 475581 557636
rect 483611 557700 483677 557701
rect 483611 557636 483612 557700
rect 483676 557636 483677 557700
rect 483611 557635 483677 557636
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 546054 437004 557000
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 549654 440604 557000
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 553254 444204 557000
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 524454 451404 557000
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 528054 455004 557000
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 531654 458604 557000
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 535254 462204 557000
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 542454 469404 557000
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 546054 473004 557000
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 549654 476604 557000
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 553254 480204 557000
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 524454 487404 557000
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 528054 491004 557000
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 531654 494604 557000
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 535254 498204 557000
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 542454 505404 557000
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 546054 509004 557000
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 549654 512604 557000
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 553254 516204 557000
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 550587 697372 550653 697373
rect 550587 697308 550588 697372
rect 550652 697308 550653 697372
rect 550587 697307 550653 697308
rect 550590 696965 550650 697307
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 550587 696964 550653 696965
rect 550587 696900 550588 696964
rect 550652 696900 550653 696964
rect 550587 696899 550653 696900
rect 551604 696934 552204 697018
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 550587 686356 550653 686357
rect 550587 686292 550588 686356
rect 550652 686292 550653 686356
rect 550587 686291 550653 686292
rect 550590 685949 550650 686291
rect 550587 685948 550653 685949
rect 550587 685884 550588 685948
rect 550652 685884 550653 685948
rect 550587 685883 550653 685884
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 136982 643018 137218 643254
rect 136982 642698 137218 642934
rect 136982 639418 137218 639654
rect 136982 639098 137218 639334
rect 136982 635818 137218 636054
rect 136982 635498 137218 635734
rect 136982 632218 137218 632454
rect 136982 631898 137218 632134
rect 136536 625018 136772 625254
rect 136536 624698 136772 624934
rect 136536 621418 136772 621654
rect 136536 621098 136772 621334
rect 136536 617818 136772 618054
rect 136536 617498 136772 617734
rect 136536 614218 136772 614454
rect 136536 613898 136772 614134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 136982 607018 137218 607254
rect 136982 606698 137218 606934
rect 136982 603418 137218 603654
rect 136982 603098 137218 603334
rect 136982 599818 137218 600054
rect 136982 599498 137218 599734
rect 136982 596218 137218 596454
rect 136982 595898 137218 596134
rect 136536 589018 136772 589254
rect 136536 588698 136772 588934
rect 136536 585418 136772 585654
rect 136536 585098 136772 585334
rect 136536 581818 136772 582054
rect 136536 581498 136772 581734
rect 136536 578218 136772 578454
rect 136536 577898 136772 578134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 136982 571018 137218 571254
rect 136982 570698 137218 570934
rect 136982 567418 137218 567654
rect 136982 567098 137218 567334
rect 136982 563818 137218 564054
rect 136982 563498 137218 563734
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 266982 643018 267218 643254
rect 266982 642698 267218 642934
rect 266982 639418 267218 639654
rect 266982 639098 267218 639334
rect 266982 635818 267218 636054
rect 266982 635498 267218 635734
rect 266982 632218 267218 632454
rect 266982 631898 267218 632134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 266536 625018 266772 625254
rect 266536 624698 266772 624934
rect 266536 621418 266772 621654
rect 266536 621098 266772 621334
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 266536 617818 266772 618054
rect 266536 617498 266772 617734
rect 266536 614218 266772 614454
rect 266536 613898 266772 614134
rect 266982 607018 267218 607254
rect 266982 606698 267218 606934
rect 266982 603418 267218 603654
rect 266982 603098 267218 603334
rect 266982 599818 267218 600054
rect 266982 599498 267218 599734
rect 266982 596218 267218 596454
rect 266982 595898 267218 596134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 266536 589018 266772 589254
rect 266536 588698 266772 588934
rect 266536 585418 266772 585654
rect 266536 585098 266772 585334
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 266536 581818 266772 582054
rect 266536 581498 266772 581734
rect 266536 578218 266772 578454
rect 266536 577898 266772 578134
rect 266982 571018 267218 571254
rect 266982 570698 267218 570934
rect 266982 567418 267218 567654
rect 266982 567098 267218 567334
rect 266982 563818 267218 564054
rect 266982 563498 267218 563734
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 79610 535018 79846 535254
rect 79610 534698 79846 534934
rect 79610 531418 79846 531654
rect 79610 531098 79846 531334
rect 79610 527818 79846 528054
rect 79610 527498 79846 527734
rect 79610 524218 79846 524454
rect 79610 523898 79846 524134
rect 64250 517018 64486 517254
rect 64250 516698 64486 516934
rect 64250 513418 64486 513654
rect 64250 513098 64486 513334
rect 64250 509818 64486 510054
rect 64250 509498 64486 509734
rect 64250 506218 64486 506454
rect 64250 505898 64486 506134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 79610 499018 79846 499254
rect 79610 498698 79846 498934
rect 79610 495418 79846 495654
rect 79610 495098 79846 495334
rect 79610 491818 79846 492054
rect 79610 491498 79846 491734
rect 79610 488218 79846 488454
rect 79610 487898 79846 488134
rect 64250 481018 64486 481254
rect 64250 480698 64486 480934
rect 64250 477418 64486 477654
rect 64250 477098 64486 477334
rect 64250 473818 64486 474054
rect 64250 473498 64486 473734
rect 64250 470218 64486 470454
rect 64250 469898 64486 470134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 79610 463018 79846 463254
rect 79610 462698 79846 462934
rect 79610 459418 79846 459654
rect 79610 459098 79846 459334
rect 79610 455818 79846 456054
rect 79610 455498 79846 455734
rect 79610 452218 79846 452454
rect 79610 451898 79846 452134
rect 64250 445018 64486 445254
rect 64250 444698 64486 444934
rect 64250 441418 64486 441654
rect 64250 441098 64486 441334
rect 64250 437818 64486 438054
rect 64250 437498 64486 437734
rect 64250 434218 64486 434454
rect 64250 433898 64486 434134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 79610 427018 79846 427254
rect 79610 426698 79846 426934
rect 79610 423418 79846 423654
rect 79610 423098 79846 423334
rect 79610 419818 79846 420054
rect 79610 419498 79846 419734
rect 79610 416218 79846 416454
rect 79610 415898 79846 416134
rect 64250 409018 64486 409254
rect 64250 408698 64486 408934
rect 64250 405418 64486 405654
rect 64250 405098 64486 405334
rect 64250 401818 64486 402054
rect 64250 401498 64486 401734
rect 64250 398218 64486 398454
rect 64250 397898 64486 398134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 79610 391018 79846 391254
rect 79610 390698 79846 390934
rect 79610 387418 79846 387654
rect 79610 387098 79846 387334
rect 79610 383818 79846 384054
rect 79610 383498 79846 383734
rect 79610 380218 79846 380454
rect 79610 379898 79846 380134
rect 64250 373018 64486 373254
rect 64250 372698 64486 372934
rect 64250 369418 64486 369654
rect 64250 369098 64486 369334
rect 64250 365818 64486 366054
rect 64250 365498 64486 365734
rect 64250 362218 64486 362454
rect 64250 361898 64486 362134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 79610 355018 79846 355254
rect 79610 354698 79846 354934
rect 79610 351418 79846 351654
rect 79610 351098 79846 351334
rect 79610 347818 79846 348054
rect 79610 347498 79846 347734
rect 79610 344218 79846 344454
rect 79610 343898 79846 344134
rect 64250 337018 64486 337254
rect 64250 336698 64486 336934
rect 64250 333418 64486 333654
rect 64250 333098 64486 333334
rect 64250 329818 64486 330054
rect 64250 329498 64486 329734
rect 64250 326218 64486 326454
rect 64250 325898 64486 326134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 79610 319018 79846 319254
rect 79610 318698 79846 318934
rect 79610 315418 79846 315654
rect 79610 315098 79846 315334
rect 79610 311818 79846 312054
rect 79610 311498 79846 311734
rect 79610 308218 79846 308454
rect 79610 307898 79846 308134
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 386982 643018 387218 643254
rect 386982 642698 387218 642934
rect 386982 639418 387218 639654
rect 386982 639098 387218 639334
rect 386982 635818 387218 636054
rect 386982 635498 387218 635734
rect 386982 632218 387218 632454
rect 386982 631898 387218 632134
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 386536 625018 386772 625254
rect 386536 624698 386772 624934
rect 386536 621418 386772 621654
rect 386536 621098 386772 621334
rect 386536 617818 386772 618054
rect 386536 617498 386772 617734
rect 386536 614218 386772 614454
rect 386536 613898 386772 614134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 386982 607018 387218 607254
rect 386982 606698 387218 606934
rect 386982 603418 387218 603654
rect 386982 603098 387218 603334
rect 386982 599818 387218 600054
rect 386982 599498 387218 599734
rect 386982 596218 387218 596454
rect 386982 595898 387218 596134
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 386536 589018 386772 589254
rect 386536 588698 386772 588934
rect 386536 585418 386772 585654
rect 386536 585098 386772 585334
rect 386536 581818 386772 582054
rect 386536 581498 386772 581734
rect 386536 578218 386772 578454
rect 386536 577898 386772 578134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 386982 571018 387218 571254
rect 386982 570698 387218 570934
rect 386982 567418 387218 567654
rect 386982 567098 387218 567334
rect 386982 563818 387218 564054
rect 386982 563498 387218 563734
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 516982 643018 517218 643254
rect 516982 642698 517218 642934
rect 516982 639418 517218 639654
rect 516982 639098 517218 639334
rect 516982 635818 517218 636054
rect 516982 635498 517218 635734
rect 516982 632218 517218 632454
rect 516982 631898 517218 632134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 516536 625018 516772 625254
rect 516536 624698 516772 624934
rect 516536 621418 516772 621654
rect 516536 621098 516772 621334
rect 516536 617818 516772 618054
rect 516536 617498 516772 617734
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 516536 614218 516772 614454
rect 516536 613898 516772 614134
rect 516982 607018 517218 607254
rect 516982 606698 517218 606934
rect 516982 603418 517218 603654
rect 516982 603098 517218 603334
rect 516982 599818 517218 600054
rect 516982 599498 517218 599734
rect 516982 596218 517218 596454
rect 516982 595898 517218 596134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 516536 589018 516772 589254
rect 516536 588698 516772 588934
rect 516536 585418 516772 585654
rect 516536 585098 516772 585334
rect 516536 581818 516772 582054
rect 516536 581498 516772 581734
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 516536 578218 516772 578454
rect 516536 577898 516772 578134
rect 516982 571018 517218 571254
rect 516982 570698 517218 570934
rect 516982 567418 517218 567654
rect 516982 567098 517218 567334
rect 516982 563818 517218 564054
rect 516982 563498 517218 563734
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 551786 696698 552022 696934
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 292404 654076 293004 654078
rect 400404 654076 401004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 292586 654054
rect 292822 653818 400586 654054
rect 400822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 292586 653734
rect 292822 653498 400586 653734
rect 400822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 292404 653474 293004 653476
rect 400404 653474 401004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 288804 650476 289404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 288986 650454
rect 289222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 288986 650134
rect 289222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 288804 649874 289404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 136938 643276 137262 643278
rect 173604 643276 174204 643278
rect 266938 643276 267262 643278
rect 281604 643276 282204 643278
rect 386938 643276 387262 643278
rect 425604 643276 426204 643278
rect 516938 643276 517262 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 136982 643254
rect 137218 643018 173786 643254
rect 174022 643018 266982 643254
rect 267218 643018 281786 643254
rect 282022 643018 386982 643254
rect 387218 643018 425786 643254
rect 426022 643018 516982 643254
rect 517218 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 136982 642934
rect 137218 642698 173786 642934
rect 174022 642698 266982 642934
rect 267218 642698 281786 642934
rect 282022 642698 386982 642934
rect 387218 642698 425786 642934
rect 426022 642698 516982 642934
rect 517218 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 136938 642674 137262 642676
rect 173604 642674 174204 642676
rect 266938 642674 267262 642676
rect 281604 642674 282204 642676
rect 386938 642674 387262 642676
rect 425604 642674 426204 642676
rect 516938 642674 517262 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 136938 639676 137262 639678
rect 170004 639676 170604 639678
rect 266938 639676 267262 639678
rect 278004 639676 278604 639678
rect 386938 639676 387262 639678
rect 422004 639676 422604 639678
rect 516938 639676 517262 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 136982 639654
rect 137218 639418 170186 639654
rect 170422 639418 266982 639654
rect 267218 639418 278186 639654
rect 278422 639418 386982 639654
rect 387218 639418 422186 639654
rect 422422 639418 516982 639654
rect 517218 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 136982 639334
rect 137218 639098 170186 639334
rect 170422 639098 266982 639334
rect 267218 639098 278186 639334
rect 278422 639098 386982 639334
rect 387218 639098 422186 639334
rect 422422 639098 516982 639334
rect 517218 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 136938 639074 137262 639076
rect 170004 639074 170604 639076
rect 266938 639074 267262 639076
rect 278004 639074 278604 639076
rect 386938 639074 387262 639076
rect 422004 639074 422604 639076
rect 516938 639074 517262 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 136938 636076 137262 636078
rect 166404 636076 167004 636078
rect 266938 636076 267262 636078
rect 274404 636076 275004 636078
rect 386938 636076 387262 636078
rect 418404 636076 419004 636078
rect 516938 636076 517262 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 136982 636054
rect 137218 635818 166586 636054
rect 166822 635818 266982 636054
rect 267218 635818 274586 636054
rect 274822 635818 386982 636054
rect 387218 635818 418586 636054
rect 418822 635818 516982 636054
rect 517218 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 136982 635734
rect 137218 635498 166586 635734
rect 166822 635498 266982 635734
rect 267218 635498 274586 635734
rect 274822 635498 386982 635734
rect 387218 635498 418586 635734
rect 418822 635498 516982 635734
rect 517218 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 136938 635474 137262 635476
rect 166404 635474 167004 635476
rect 266938 635474 267262 635476
rect 274404 635474 275004 635476
rect 386938 635474 387262 635476
rect 418404 635474 419004 635476
rect 516938 635474 517262 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 136938 632476 137262 632478
rect 162804 632476 163404 632478
rect 266938 632476 267262 632478
rect 270804 632476 271404 632478
rect 386938 632476 387262 632478
rect 414804 632476 415404 632478
rect 516938 632476 517262 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 136982 632454
rect 137218 632218 162986 632454
rect 163222 632218 266982 632454
rect 267218 632218 270986 632454
rect 271222 632218 386982 632454
rect 387218 632218 414986 632454
rect 415222 632218 516982 632454
rect 517218 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 136982 632134
rect 137218 631898 162986 632134
rect 163222 631898 266982 632134
rect 267218 631898 270986 632134
rect 271222 631898 386982 632134
rect 387218 631898 414986 632134
rect 415222 631898 516982 632134
rect 517218 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 136938 631874 137262 631876
rect 162804 631874 163404 631876
rect 266938 631874 267262 631876
rect 270804 631874 271404 631876
rect 386938 631874 387262 631876
rect 414804 631874 415404 631876
rect 516938 631874 517262 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 136494 625276 136814 625278
rect 155604 625276 156204 625278
rect 266494 625276 266814 625278
rect 299604 625276 300204 625278
rect 386494 625276 386814 625278
rect 407604 625276 408204 625278
rect 516494 625276 516814 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 136536 625254
rect 136772 625018 155786 625254
rect 156022 625018 266536 625254
rect 266772 625018 299786 625254
rect 300022 625018 386536 625254
rect 386772 625018 407786 625254
rect 408022 625018 516536 625254
rect 516772 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 136536 624934
rect 136772 624698 155786 624934
rect 156022 624698 266536 624934
rect 266772 624698 299786 624934
rect 300022 624698 386536 624934
rect 386772 624698 407786 624934
rect 408022 624698 516536 624934
rect 516772 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 136494 624674 136814 624676
rect 155604 624674 156204 624676
rect 266494 624674 266814 624676
rect 299604 624674 300204 624676
rect 386494 624674 386814 624676
rect 407604 624674 408204 624676
rect 516494 624674 516814 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 136494 621676 136814 621678
rect 152004 621676 152604 621678
rect 266494 621676 266814 621678
rect 296004 621676 296604 621678
rect 386494 621676 386814 621678
rect 404004 621676 404604 621678
rect 516494 621676 516814 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 136536 621654
rect 136772 621418 152186 621654
rect 152422 621418 266536 621654
rect 266772 621418 296186 621654
rect 296422 621418 386536 621654
rect 386772 621418 404186 621654
rect 404422 621418 516536 621654
rect 516772 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 136536 621334
rect 136772 621098 152186 621334
rect 152422 621098 266536 621334
rect 266772 621098 296186 621334
rect 296422 621098 386536 621334
rect 386772 621098 404186 621334
rect 404422 621098 516536 621334
rect 516772 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 136494 621074 136814 621076
rect 152004 621074 152604 621076
rect 266494 621074 266814 621076
rect 296004 621074 296604 621076
rect 386494 621074 386814 621076
rect 404004 621074 404604 621076
rect 516494 621074 516814 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 136494 618076 136814 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 266494 618076 266814 618078
rect 292404 618076 293004 618078
rect 386494 618076 386814 618078
rect 400404 618076 401004 618078
rect 516494 618076 516814 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 136536 618054
rect 136772 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 266536 618054
rect 266772 617818 292586 618054
rect 292822 617818 386536 618054
rect 386772 617818 400586 618054
rect 400822 617818 516536 618054
rect 516772 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 136536 617734
rect 136772 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 266536 617734
rect 266772 617498 292586 617734
rect 292822 617498 386536 617734
rect 386772 617498 400586 617734
rect 400822 617498 516536 617734
rect 516772 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 136494 617474 136814 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 266494 617474 266814 617476
rect 292404 617474 293004 617476
rect 386494 617474 386814 617476
rect 400404 617474 401004 617476
rect 516494 617474 516814 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 136494 614476 136814 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 266494 614476 266814 614478
rect 288804 614476 289404 614478
rect 386494 614476 386814 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 516494 614476 516814 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 136536 614454
rect 136772 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 266536 614454
rect 266772 614218 288986 614454
rect 289222 614218 386536 614454
rect 386772 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 516536 614454
rect 516772 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 136536 614134
rect 136772 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 266536 614134
rect 266772 613898 288986 614134
rect 289222 613898 386536 614134
rect 386772 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 516536 614134
rect 516772 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 136494 613874 136814 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 266494 613874 266814 613876
rect 288804 613874 289404 613876
rect 386494 613874 386814 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 516494 613874 516814 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 136938 607276 137262 607278
rect 173604 607276 174204 607278
rect 266938 607276 267262 607278
rect 281604 607276 282204 607278
rect 386938 607276 387262 607278
rect 425604 607276 426204 607278
rect 516938 607276 517262 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 136982 607254
rect 137218 607018 173786 607254
rect 174022 607018 266982 607254
rect 267218 607018 281786 607254
rect 282022 607018 386982 607254
rect 387218 607018 425786 607254
rect 426022 607018 516982 607254
rect 517218 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 136982 606934
rect 137218 606698 173786 606934
rect 174022 606698 266982 606934
rect 267218 606698 281786 606934
rect 282022 606698 386982 606934
rect 387218 606698 425786 606934
rect 426022 606698 516982 606934
rect 517218 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 136938 606674 137262 606676
rect 173604 606674 174204 606676
rect 266938 606674 267262 606676
rect 281604 606674 282204 606676
rect 386938 606674 387262 606676
rect 425604 606674 426204 606676
rect 516938 606674 517262 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 136938 603676 137262 603678
rect 170004 603676 170604 603678
rect 266938 603676 267262 603678
rect 278004 603676 278604 603678
rect 386938 603676 387262 603678
rect 422004 603676 422604 603678
rect 516938 603676 517262 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 136982 603654
rect 137218 603418 170186 603654
rect 170422 603418 266982 603654
rect 267218 603418 278186 603654
rect 278422 603418 386982 603654
rect 387218 603418 422186 603654
rect 422422 603418 516982 603654
rect 517218 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 136982 603334
rect 137218 603098 170186 603334
rect 170422 603098 266982 603334
rect 267218 603098 278186 603334
rect 278422 603098 386982 603334
rect 387218 603098 422186 603334
rect 422422 603098 516982 603334
rect 517218 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 136938 603074 137262 603076
rect 170004 603074 170604 603076
rect 266938 603074 267262 603076
rect 278004 603074 278604 603076
rect 386938 603074 387262 603076
rect 422004 603074 422604 603076
rect 516938 603074 517262 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 136938 600076 137262 600078
rect 166404 600076 167004 600078
rect 266938 600076 267262 600078
rect 274404 600076 275004 600078
rect 386938 600076 387262 600078
rect 418404 600076 419004 600078
rect 516938 600076 517262 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 136982 600054
rect 137218 599818 166586 600054
rect 166822 599818 266982 600054
rect 267218 599818 274586 600054
rect 274822 599818 386982 600054
rect 387218 599818 418586 600054
rect 418822 599818 516982 600054
rect 517218 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 136982 599734
rect 137218 599498 166586 599734
rect 166822 599498 266982 599734
rect 267218 599498 274586 599734
rect 274822 599498 386982 599734
rect 387218 599498 418586 599734
rect 418822 599498 516982 599734
rect 517218 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 136938 599474 137262 599476
rect 166404 599474 167004 599476
rect 266938 599474 267262 599476
rect 274404 599474 275004 599476
rect 386938 599474 387262 599476
rect 418404 599474 419004 599476
rect 516938 599474 517262 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 136938 596476 137262 596478
rect 162804 596476 163404 596478
rect 266938 596476 267262 596478
rect 270804 596476 271404 596478
rect 386938 596476 387262 596478
rect 414804 596476 415404 596478
rect 516938 596476 517262 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 136982 596454
rect 137218 596218 162986 596454
rect 163222 596218 266982 596454
rect 267218 596218 270986 596454
rect 271222 596218 386982 596454
rect 387218 596218 414986 596454
rect 415222 596218 516982 596454
rect 517218 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 136982 596134
rect 137218 595898 162986 596134
rect 163222 595898 266982 596134
rect 267218 595898 270986 596134
rect 271222 595898 386982 596134
rect 387218 595898 414986 596134
rect 415222 595898 516982 596134
rect 517218 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 136938 595874 137262 595876
rect 162804 595874 163404 595876
rect 266938 595874 267262 595876
rect 270804 595874 271404 595876
rect 386938 595874 387262 595876
rect 414804 595874 415404 595876
rect 516938 595874 517262 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 136494 589276 136814 589278
rect 155604 589276 156204 589278
rect 266494 589276 266814 589278
rect 299604 589276 300204 589278
rect 386494 589276 386814 589278
rect 407604 589276 408204 589278
rect 516494 589276 516814 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 136536 589254
rect 136772 589018 155786 589254
rect 156022 589018 266536 589254
rect 266772 589018 299786 589254
rect 300022 589018 386536 589254
rect 386772 589018 407786 589254
rect 408022 589018 516536 589254
rect 516772 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 136536 588934
rect 136772 588698 155786 588934
rect 156022 588698 266536 588934
rect 266772 588698 299786 588934
rect 300022 588698 386536 588934
rect 386772 588698 407786 588934
rect 408022 588698 516536 588934
rect 516772 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 136494 588674 136814 588676
rect 155604 588674 156204 588676
rect 266494 588674 266814 588676
rect 299604 588674 300204 588676
rect 386494 588674 386814 588676
rect 407604 588674 408204 588676
rect 516494 588674 516814 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 136494 585676 136814 585678
rect 152004 585676 152604 585678
rect 266494 585676 266814 585678
rect 296004 585676 296604 585678
rect 386494 585676 386814 585678
rect 404004 585676 404604 585678
rect 516494 585676 516814 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 136536 585654
rect 136772 585418 152186 585654
rect 152422 585418 266536 585654
rect 266772 585418 296186 585654
rect 296422 585418 386536 585654
rect 386772 585418 404186 585654
rect 404422 585418 516536 585654
rect 516772 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 136536 585334
rect 136772 585098 152186 585334
rect 152422 585098 266536 585334
rect 266772 585098 296186 585334
rect 296422 585098 386536 585334
rect 386772 585098 404186 585334
rect 404422 585098 516536 585334
rect 516772 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 136494 585074 136814 585076
rect 152004 585074 152604 585076
rect 266494 585074 266814 585076
rect 296004 585074 296604 585076
rect 386494 585074 386814 585076
rect 404004 585074 404604 585076
rect 516494 585074 516814 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 136494 582076 136814 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 266494 582076 266814 582078
rect 292404 582076 293004 582078
rect 386494 582076 386814 582078
rect 400404 582076 401004 582078
rect 516494 582076 516814 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 136536 582054
rect 136772 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 266536 582054
rect 266772 581818 292586 582054
rect 292822 581818 386536 582054
rect 386772 581818 400586 582054
rect 400822 581818 516536 582054
rect 516772 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 136536 581734
rect 136772 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 266536 581734
rect 266772 581498 292586 581734
rect 292822 581498 386536 581734
rect 386772 581498 400586 581734
rect 400822 581498 516536 581734
rect 516772 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 136494 581474 136814 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 266494 581474 266814 581476
rect 292404 581474 293004 581476
rect 386494 581474 386814 581476
rect 400404 581474 401004 581476
rect 516494 581474 516814 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 136494 578476 136814 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 266494 578476 266814 578478
rect 288804 578476 289404 578478
rect 386494 578476 386814 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 516494 578476 516814 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 136536 578454
rect 136772 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 266536 578454
rect 266772 578218 288986 578454
rect 289222 578218 386536 578454
rect 386772 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 516536 578454
rect 516772 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 136536 578134
rect 136772 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 266536 578134
rect 266772 577898 288986 578134
rect 289222 577898 386536 578134
rect 386772 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 516536 578134
rect 516772 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 136494 577874 136814 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 266494 577874 266814 577876
rect 288804 577874 289404 577876
rect 386494 577874 386814 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 516494 577874 516814 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 136938 571276 137262 571278
rect 173604 571276 174204 571278
rect 266938 571276 267262 571278
rect 281604 571276 282204 571278
rect 386938 571276 387262 571278
rect 425604 571276 426204 571278
rect 516938 571276 517262 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 136982 571254
rect 137218 571018 173786 571254
rect 174022 571018 266982 571254
rect 267218 571018 281786 571254
rect 282022 571018 386982 571254
rect 387218 571018 425786 571254
rect 426022 571018 516982 571254
rect 517218 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 136982 570934
rect 137218 570698 173786 570934
rect 174022 570698 266982 570934
rect 267218 570698 281786 570934
rect 282022 570698 386982 570934
rect 387218 570698 425786 570934
rect 426022 570698 516982 570934
rect 517218 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 136938 570674 137262 570676
rect 173604 570674 174204 570676
rect 266938 570674 267262 570676
rect 281604 570674 282204 570676
rect 386938 570674 387262 570676
rect 425604 570674 426204 570676
rect 516938 570674 517262 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 136938 567676 137262 567678
rect 170004 567676 170604 567678
rect 266938 567676 267262 567678
rect 278004 567676 278604 567678
rect 386938 567676 387262 567678
rect 422004 567676 422604 567678
rect 516938 567676 517262 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 136982 567654
rect 137218 567418 170186 567654
rect 170422 567418 266982 567654
rect 267218 567418 278186 567654
rect 278422 567418 386982 567654
rect 387218 567418 422186 567654
rect 422422 567418 516982 567654
rect 517218 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 136982 567334
rect 137218 567098 170186 567334
rect 170422 567098 266982 567334
rect 267218 567098 278186 567334
rect 278422 567098 386982 567334
rect 387218 567098 422186 567334
rect 422422 567098 516982 567334
rect 517218 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 136938 567074 137262 567076
rect 170004 567074 170604 567076
rect 266938 567074 267262 567076
rect 278004 567074 278604 567076
rect 386938 567074 387262 567076
rect 422004 567074 422604 567076
rect 516938 567074 517262 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 136938 564076 137262 564078
rect 166404 564076 167004 564078
rect 266938 564076 267262 564078
rect 274404 564076 275004 564078
rect 386938 564076 387262 564078
rect 418404 564076 419004 564078
rect 516938 564076 517262 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 136982 564054
rect 137218 563818 166586 564054
rect 166822 563818 266982 564054
rect 267218 563818 274586 564054
rect 274822 563818 386982 564054
rect 387218 563818 418586 564054
rect 418822 563818 516982 564054
rect 517218 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 136982 563734
rect 137218 563498 166586 563734
rect 166822 563498 266982 563734
rect 267218 563498 274586 563734
rect 274822 563498 386982 563734
rect 387218 563498 418586 563734
rect 418822 563498 516982 563734
rect 517218 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 136938 563474 137262 563476
rect 166404 563474 167004 563476
rect 266938 563474 267262 563476
rect 274404 563474 275004 563476
rect 386938 563474 387262 563476
rect 418404 563474 419004 563476
rect 516938 563474 517262 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 162804 560476 163404 560478
rect 270804 560476 271404 560478
rect 414804 560476 415404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 162986 560454
rect 163222 560218 270986 560454
rect 271222 560218 414986 560454
rect 415222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 162986 560134
rect 163222 559898 270986 560134
rect 271222 559898 414986 560134
rect 415222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 162804 559874 163404 559876
rect 270804 559874 271404 559876
rect 414804 559874 415404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 79568 535276 79888 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 79610 535254
rect 79846 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 79610 534934
rect 79846 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 79568 534674 79888 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 79568 531676 79888 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 79610 531654
rect 79846 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 79610 531334
rect 79846 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 79568 531074 79888 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 79568 528076 79888 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 79610 528054
rect 79846 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 79610 527734
rect 79846 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 79568 527474 79888 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 79568 524476 79888 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 79610 524454
rect 79846 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 79610 524134
rect 79846 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 79568 523874 79888 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 64208 517276 64528 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 64250 517254
rect 64486 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 64250 516934
rect 64486 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 64208 516674 64528 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 64208 513676 64528 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 64250 513654
rect 64486 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 64250 513334
rect 64486 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 64208 513074 64528 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 64208 510076 64528 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 64250 510054
rect 64486 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 64250 509734
rect 64486 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 64208 509474 64528 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 64208 506476 64528 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 64250 506454
rect 64486 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 64250 506134
rect 64486 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 64208 505874 64528 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 79568 499276 79888 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 79610 499254
rect 79846 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 79610 498934
rect 79846 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 79568 498674 79888 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 79568 495676 79888 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 79610 495654
rect 79846 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 79610 495334
rect 79846 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 79568 495074 79888 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 79568 492076 79888 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 79610 492054
rect 79846 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 79610 491734
rect 79846 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 79568 491474 79888 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 79568 488476 79888 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 79610 488454
rect 79846 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 79610 488134
rect 79846 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 79568 487874 79888 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 64208 481276 64528 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 64250 481254
rect 64486 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 64250 480934
rect 64486 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 64208 480674 64528 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 64208 477676 64528 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 64250 477654
rect 64486 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 64250 477334
rect 64486 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 64208 477074 64528 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 64208 474076 64528 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 64250 474054
rect 64486 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 64250 473734
rect 64486 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 64208 473474 64528 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 64208 470476 64528 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 64250 470454
rect 64486 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 64250 470134
rect 64486 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 64208 469874 64528 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 79568 463276 79888 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 79610 463254
rect 79846 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 79610 462934
rect 79846 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 79568 462674 79888 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 79568 459676 79888 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 79610 459654
rect 79846 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 79610 459334
rect 79846 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 79568 459074 79888 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 79568 456076 79888 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 79610 456054
rect 79846 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 79610 455734
rect 79846 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 79568 455474 79888 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 79568 452476 79888 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 79610 452454
rect 79846 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 79610 452134
rect 79846 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 79568 451874 79888 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 64208 445276 64528 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 64250 445254
rect 64486 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 64250 444934
rect 64486 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 64208 444674 64528 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 64208 441676 64528 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 64250 441654
rect 64486 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 64250 441334
rect 64486 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 64208 441074 64528 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 64208 438076 64528 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 64250 438054
rect 64486 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 64250 437734
rect 64486 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 64208 437474 64528 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 64208 434476 64528 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 64250 434454
rect 64486 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 64250 434134
rect 64486 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 64208 433874 64528 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 79568 427276 79888 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 79610 427254
rect 79846 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 79610 426934
rect 79846 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 79568 426674 79888 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 79568 423676 79888 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 79610 423654
rect 79846 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 79610 423334
rect 79846 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 79568 423074 79888 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 79568 420076 79888 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 79610 420054
rect 79846 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 79610 419734
rect 79846 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 79568 419474 79888 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 79568 416476 79888 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 79610 416454
rect 79846 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 79610 416134
rect 79846 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 79568 415874 79888 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 64208 409276 64528 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 64250 409254
rect 64486 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 64250 408934
rect 64486 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 64208 408674 64528 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 64208 405676 64528 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 64250 405654
rect 64486 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 64250 405334
rect 64486 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 64208 405074 64528 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 64208 402076 64528 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 64250 402054
rect 64486 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 64250 401734
rect 64486 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 64208 401474 64528 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 64208 398476 64528 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 64250 398454
rect 64486 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 64250 398134
rect 64486 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 64208 397874 64528 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 79568 391276 79888 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 79610 391254
rect 79846 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 79610 390934
rect 79846 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 79568 390674 79888 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 79568 387676 79888 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 79610 387654
rect 79846 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 79610 387334
rect 79846 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 79568 387074 79888 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 79568 384076 79888 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 79610 384054
rect 79846 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 79610 383734
rect 79846 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 79568 383474 79888 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 79568 380476 79888 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 79610 380454
rect 79846 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 79610 380134
rect 79846 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 79568 379874 79888 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 64208 373276 64528 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 64250 373254
rect 64486 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 64250 372934
rect 64486 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 64208 372674 64528 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 64208 369676 64528 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 64250 369654
rect 64486 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 64250 369334
rect 64486 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 64208 369074 64528 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 64208 366076 64528 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 64250 366054
rect 64486 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 64250 365734
rect 64486 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 64208 365474 64528 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 64208 362476 64528 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 64250 362454
rect 64486 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 64250 362134
rect 64486 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 64208 361874 64528 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 79568 355276 79888 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 79610 355254
rect 79846 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 79610 354934
rect 79846 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 79568 354674 79888 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 79568 351676 79888 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 79610 351654
rect 79846 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 79610 351334
rect 79846 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 79568 351074 79888 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 79568 348076 79888 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 79610 348054
rect 79846 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 79610 347734
rect 79846 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 79568 347474 79888 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 79568 344476 79888 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 79610 344454
rect 79846 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 79610 344134
rect 79846 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 79568 343874 79888 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 64208 337276 64528 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 64250 337254
rect 64486 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 64250 336934
rect 64486 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 64208 336674 64528 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 64208 333676 64528 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 64250 333654
rect 64486 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 64250 333334
rect 64486 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 64208 333074 64528 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 64208 330076 64528 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 64250 330054
rect 64486 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 64250 329734
rect 64486 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 64208 329474 64528 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 64208 326476 64528 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 64250 326454
rect 64486 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 64250 326134
rect 64486 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 64208 325874 64528 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 79568 319276 79888 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 79610 319254
rect 79846 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 79610 318934
rect 79846 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 79568 318674 79888 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 79568 315676 79888 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 79610 315654
rect 79846 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 79610 315334
rect 79846 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 79568 315074 79888 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 79568 312076 79888 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 79610 312054
rect 79846 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 79610 311734
rect 79846 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 79568 311474 79888 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 79568 308476 79888 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 79610 308454
rect 79846 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 79610 308134
rect 79846 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 79568 307874 79888 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use sram_1rw1r_32_256_8_sky130  sram3
timestamp 1608703685
transform 1 0 440000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram2
timestamp 1608703685
transform 1 0 310000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram1
timestamp 1608703685
transform 1 0 190000 0 1 560000
box 0 0 77296 91247
use sram_1rw1r_32_256_8_sky130  sram0
timestamp 1608703685
transform 1 0 60000 0 1 560000
box 0 0 77296 91247
use hs32_core1  core1
timestamp 1608703685
transform 1 0 60000 0 1 300000
box 0 0 220000 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
