VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1099.930 BY 1100.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 126.520 1099.930 127.120 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 228.520 1099.930 229.120 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 238.720 1099.930 239.320 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 248.920 1099.930 249.520 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 259.120 1099.930 259.720 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 269.320 1099.930 269.920 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 279.520 1099.930 280.120 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 136.720 1099.930 137.320 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 146.920 1099.930 147.520 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 157.120 1099.930 157.720 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 167.320 1099.930 167.920 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 177.520 1099.930 178.120 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 187.720 1099.930 188.320 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 197.920 1099.930 198.520 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 208.120 1099.930 208.720 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 218.320 1099.930 218.920 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.580 1096.000 108.860 1100.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.540 1096.000 212.820 1100.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.660 1096.000 222.940 1100.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 233.240 1096.000 233.520 1100.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.360 1096.000 243.640 1100.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.940 1096.000 254.220 1100.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 264.060 1096.000 264.340 1100.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.160 1096.000 119.440 1100.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.280 1096.000 129.560 1100.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.860 1096.000 140.140 1100.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.980 1096.000 150.260 1100.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 160.560 1096.000 160.840 1100.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 170.680 1096.000 170.960 1100.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.260 1096.000 181.540 1100.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.840 1096.000 192.120 1100.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.960 1096.000 202.240 1100.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 452.920 1099.930 453.520 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 554.920 1099.930 555.520 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 564.440 1099.930 565.040 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 574.640 1099.930 575.240 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 584.840 1099.930 585.440 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 595.040 1099.930 595.640 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 605.240 1099.930 605.840 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 615.440 1099.930 616.040 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 625.640 1099.930 626.240 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 635.840 1099.930 636.440 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 646.040 1099.930 646.640 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 463.120 1099.930 463.720 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 656.240 1099.930 656.840 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 666.440 1099.930 667.040 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 676.640 1099.930 677.240 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 686.840 1099.930 687.440 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 697.040 1099.930 697.640 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 707.240 1099.930 707.840 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 717.440 1099.930 718.040 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 727.640 1099.930 728.240 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 737.840 1099.930 738.440 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 748.040 1099.930 748.640 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 473.320 1099.930 473.920 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 758.240 1099.930 758.840 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 768.440 1099.930 769.040 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 483.520 1099.930 484.120 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 493.720 1099.930 494.320 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 503.920 1099.930 504.520 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 514.120 1099.930 514.720 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 524.320 1099.930 524.920 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 534.520 1099.930 535.120 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 544.720 1099.930 545.320 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 778.640 1099.930 779.240 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 880.640 1099.930 881.240 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 890.840 1099.930 891.440 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 901.040 1099.930 901.640 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 911.240 1099.930 911.840 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 921.440 1099.930 922.040 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 931.640 1099.930 932.240 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 941.840 1099.930 942.440 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 952.040 1099.930 952.640 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 962.240 1099.930 962.840 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 972.440 1099.930 973.040 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 788.840 1099.930 789.440 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 982.640 1099.930 983.240 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 992.840 1099.930 993.440 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1003.040 1099.930 1003.640 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1013.240 1099.930 1013.840 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1023.440 1099.930 1024.040 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1033.640 1099.930 1034.240 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1043.840 1099.930 1044.440 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1054.040 1099.930 1054.640 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1064.240 1099.930 1064.840 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1074.440 1099.930 1075.040 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 799.040 1099.930 799.640 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1084.640 1099.930 1085.240 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 1094.840 1099.930 1095.440 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 809.240 1099.930 809.840 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 819.440 1099.930 820.040 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 829.640 1099.930 830.240 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 839.840 1099.930 840.440 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 850.040 1099.930 850.640 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 860.240 1099.930 860.840 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1095.930 870.440 1099.930 871.040 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.700 1096.000 440.980 1100.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.200 1096.000 544.480 1100.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.780 1096.000 555.060 1100.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.360 1096.000 565.640 1100.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.480 1096.000 575.760 1100.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.060 1096.000 586.340 1100.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.180 1096.000 596.460 1100.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 606.760 1096.000 607.040 1100.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.880 1096.000 617.160 1100.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.460 1096.000 627.740 1100.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 637.580 1096.000 637.860 1100.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.820 1096.000 451.100 1100.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.160 1096.000 648.440 1100.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.740 1096.000 659.020 1100.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.860 1096.000 669.140 1100.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.440 1096.000 679.720 1100.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.560 1096.000 689.840 1100.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.140 1096.000 700.420 1100.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 710.260 1096.000 710.540 1100.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.840 1096.000 721.120 1100.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.960 1096.000 731.240 1100.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.540 1096.000 741.820 1100.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.400 1096.000 461.680 1100.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.120 1096.000 752.400 1100.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 762.240 1096.000 762.520 1100.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.980 1096.000 472.260 1100.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 482.100 1096.000 482.380 1100.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.680 1096.000 492.960 1100.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 502.800 1096.000 503.080 1100.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.380 1096.000 513.660 1100.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.500 1096.000 523.780 1100.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.080 1096.000 534.360 1100.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.820 1096.000 773.100 1100.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.320 1096.000 876.600 1100.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.900 1096.000 887.180 1100.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 897.020 1096.000 897.300 1100.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.600 1096.000 907.880 1100.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.720 1096.000 918.000 1100.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.300 1096.000 928.580 1100.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.880 1096.000 939.160 1100.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.000 1096.000 949.280 1100.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.580 1096.000 959.860 1100.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.700 1096.000 969.980 1100.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.940 1096.000 783.220 1100.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 980.280 1096.000 980.560 1100.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.400 1096.000 990.680 1100.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.980 1096.000 1001.260 1100.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.100 1096.000 1011.380 1100.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.680 1096.000 1021.960 1100.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.260 1096.000 1032.540 1100.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1042.380 1096.000 1042.660 1100.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.960 1096.000 1053.240 1100.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.080 1096.000 1063.360 1100.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.660 1096.000 1073.940 1100.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.520 1096.000 793.800 1100.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.780 1096.000 1084.060 1100.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.360 1096.000 1094.640 1100.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.640 1096.000 803.920 1100.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.220 1096.000 814.500 1100.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.340 1096.000 824.620 1100.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.920 1096.000 835.200 1100.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 845.500 1096.000 845.780 1100.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.620 1096.000 855.900 1100.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.200 1096.000 866.480 1100.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 289.720 1099.930 290.320 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 391.720 1099.930 392.320 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 401.920 1099.930 402.520 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 412.120 1099.930 412.720 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 422.320 1099.930 422.920 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 432.520 1099.930 433.120 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 442.720 1099.930 443.320 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 299.920 1099.930 300.520 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 310.120 1099.930 310.720 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 320.320 1099.930 320.920 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 330.520 1099.930 331.120 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 340.720 1099.930 341.320 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 350.920 1099.930 351.520 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 361.120 1099.930 361.720 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 371.320 1099.930 371.920 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 381.520 1099.930 382.120 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.640 1096.000 274.920 1100.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 378.600 1096.000 378.880 1100.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.720 1096.000 389.000 1100.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 399.300 1096.000 399.580 1100.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.420 1096.000 409.700 1100.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.000 1096.000 420.280 1100.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 430.120 1096.000 430.400 1100.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.220 1096.000 285.500 1100.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 295.340 1096.000 295.620 1100.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.920 1096.000 306.200 1100.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 316.040 1096.000 316.320 1100.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 326.620 1096.000 326.900 1100.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.740 1096.000 337.020 1100.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.320 1096.000 347.600 1100.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.440 1096.000 357.720 1100.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.020 1096.000 368.300 1100.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 24.520 1099.930 25.120 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 34.720 1099.930 35.320 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 44.920 1099.930 45.520 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 55.120 1099.930 55.720 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 65.320 1099.930 65.920 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 75.520 1099.930 76.120 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 85.720 1099.930 86.320 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 95.920 1099.930 96.520 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.080 1096.000 5.360 1100.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 15.200 1096.000 15.480 1100.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.780 1096.000 26.060 1100.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.900 1096.000 36.180 1100.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.480 1096.000 46.760 1100.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.600 1096.000 56.880 1100.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.180 1096.000 67.460 1100.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.300 1096.000 77.580 1100.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 106.120 1099.930 106.720 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 116.320 1099.930 116.920 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.880 1096.000 88.160 1100.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.460 1096.000 98.740 1100.000 ;
    END
  END cpu_wen_n[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.760 0.000 239.040 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.200 0.000 912.480 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.640 0.000 918.920 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.540 0.000 925.820 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.440 0.000 932.720 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.880 0.000 939.160 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.780 0.000 946.060 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 952.220 0.000 952.500 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.120 0.000 959.400 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 966.020 0.000 966.300 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.460 0.000 972.740 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.920 0.000 306.200 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.360 0.000 979.640 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 986.260 0.000 986.540 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 992.700 0.000 992.980 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 999.600 0.000 999.880 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.500 0.000 1006.780 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.940 0.000 1013.220 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.840 0.000 1020.120 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1026.280 0.000 1026.560 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1033.180 0.000 1033.460 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1040.080 0.000 1040.360 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.820 0.000 313.100 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.520 0.000 1046.800 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.420 0.000 1053.700 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.320 0.000 1060.600 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1066.760 0.000 1067.040 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.660 0.000 1073.940 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.560 0.000 1080.840 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.000 0.000 1087.280 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.900 0.000 1094.180 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.260 0.000 319.540 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 326.160 0.000 326.440 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.060 0.000 333.340 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.500 0.000 339.780 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 346.400 0.000 346.680 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.300 0.000 353.580 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.740 0.000 360.020 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 366.640 0.000 366.920 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 245.200 0.000 245.480 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 373.540 0.000 373.820 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.980 0.000 380.260 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.880 0.000 387.160 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 393.320 0.000 393.600 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.220 0.000 400.500 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.120 0.000 407.400 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.560 0.000 413.840 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.460 0.000 420.740 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 427.360 0.000 427.640 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.800 0.000 434.080 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.100 0.000 252.380 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 447.600 0.000 447.880 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.040 0.000 454.320 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.940 0.000 461.220 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 467.380 0.000 467.660 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.280 0.000 474.560 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.180 0.000 481.460 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.620 0.000 487.900 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.520 0.000 494.800 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.420 0.000 501.700 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.000 0.000 259.280 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.860 0.000 508.140 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.760 0.000 515.040 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 521.660 0.000 521.940 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 528.100 0.000 528.380 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.000 0.000 535.280 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 541.440 0.000 541.720 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 548.340 0.000 548.620 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 555.240 0.000 555.520 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.680 0.000 561.960 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.580 0.000 568.860 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.440 0.000 265.720 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.480 0.000 575.760 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.920 0.000 582.200 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.820 0.000 589.100 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 595.720 0.000 596.000 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.160 0.000 602.440 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.060 0.000 609.340 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 615.960 0.000 616.240 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.400 0.000 622.680 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 629.300 0.000 629.580 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.740 0.000 636.020 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.340 0.000 272.620 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 642.640 0.000 642.920 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 649.540 0.000 649.820 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.980 0.000 656.260 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.880 0.000 663.160 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.780 0.000 670.060 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 676.220 0.000 676.500 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 683.120 0.000 683.400 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.020 0.000 690.300 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 696.460 0.000 696.740 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 703.360 0.000 703.640 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.240 0.000 279.520 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.800 0.000 710.080 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.700 0.000 716.980 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.600 0.000 723.880 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.040 0.000 730.320 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.940 0.000 737.220 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 743.840 0.000 744.120 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 750.280 0.000 750.560 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.180 0.000 757.460 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 764.080 0.000 764.360 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 770.520 0.000 770.800 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.680 0.000 285.960 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 777.420 0.000 777.700 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.860 0.000 784.140 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 790.760 0.000 791.040 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 797.660 0.000 797.940 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 804.100 0.000 804.380 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.000 0.000 811.280 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.900 0.000 818.180 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.340 0.000 824.620 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.240 0.000 831.520 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 838.140 0.000 838.420 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 292.580 0.000 292.860 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.580 0.000 844.860 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.480 0.000 851.760 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.380 0.000 858.660 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.820 0.000 865.100 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.720 0.000 872.000 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 878.160 0.000 878.440 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 885.060 0.000 885.340 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.960 0.000 892.240 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.400 0.000 898.680 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 905.300 0.000 905.580 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.020 0.000 299.300 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 241.060 0.000 241.340 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 914.040 0.000 914.320 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 920.940 0.000 921.220 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 927.840 0.000 928.120 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 934.280 0.000 934.560 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 941.180 0.000 941.460 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 948.080 0.000 948.360 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 954.520 0.000 954.800 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.420 0.000 961.700 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 968.320 0.000 968.600 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.760 0.000 975.040 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 308.220 0.000 308.500 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 981.660 0.000 981.940 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 988.560 0.000 988.840 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.000 0.000 995.280 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1001.900 0.000 1002.180 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.340 0.000 1008.620 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1015.240 0.000 1015.520 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1022.140 0.000 1022.420 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1028.580 0.000 1028.860 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.480 0.000 1035.760 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1042.380 0.000 1042.660 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 315.120 0.000 315.400 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1048.820 0.000 1049.100 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.720 0.000 1056.000 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1062.620 0.000 1062.900 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.060 0.000 1069.340 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1075.960 0.000 1076.240 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.400 0.000 1082.680 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1089.300 0.000 1089.580 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1096.200 0.000 1096.480 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.560 0.000 321.840 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.460 0.000 328.740 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.360 0.000 335.640 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.800 0.000 342.080 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 348.700 0.000 348.980 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.140 0.000 355.420 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.040 0.000 362.320 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.940 0.000 369.220 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.500 0.000 247.780 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.380 0.000 375.660 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.280 0.000 382.560 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.180 0.000 389.460 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 395.620 0.000 395.900 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.520 0.000 402.800 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.420 0.000 409.700 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.860 0.000 416.140 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 422.760 0.000 423.040 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.660 0.000 429.940 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 436.100 0.000 436.380 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.400 0.000 254.680 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 443.000 0.000 443.280 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 449.440 0.000 449.720 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.340 0.000 456.620 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 463.240 0.000 463.520 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 469.680 0.000 469.960 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 476.580 0.000 476.860 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.480 0.000 483.760 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.920 0.000 490.200 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.820 0.000 497.100 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.720 0.000 504.000 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.300 0.000 261.580 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 510.160 0.000 510.440 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 517.060 0.000 517.340 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 523.500 0.000 523.780 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.400 0.000 530.680 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.300 0.000 537.580 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 543.740 0.000 544.020 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 550.640 0.000 550.920 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.540 0.000 557.820 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.980 0.000 564.260 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.880 0.000 571.160 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.740 0.000 268.020 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 577.780 0.000 578.060 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 584.220 0.000 584.500 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 591.120 0.000 591.400 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 597.560 0.000 597.840 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 604.460 0.000 604.740 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 611.360 0.000 611.640 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 617.800 0.000 618.080 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 624.700 0.000 624.980 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.600 0.000 631.880 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 638.040 0.000 638.320 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.640 0.000 274.920 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.940 0.000 645.220 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.840 0.000 652.120 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 658.280 0.000 658.560 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 665.180 0.000 665.460 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 671.620 0.000 671.900 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 678.520 0.000 678.800 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.420 0.000 685.700 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 691.860 0.000 692.140 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 698.760 0.000 699.040 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.660 0.000 705.940 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 281.080 0.000 281.360 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.100 0.000 712.380 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.000 0.000 719.280 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 725.900 0.000 726.180 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 732.340 0.000 732.620 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 739.240 0.000 739.520 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.140 0.000 746.420 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 752.580 0.000 752.860 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.480 0.000 759.760 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.920 0.000 766.200 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 772.820 0.000 773.100 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.980 0.000 288.260 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 779.720 0.000 780.000 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.160 0.000 786.440 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 793.060 0.000 793.340 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.960 0.000 800.240 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.400 0.000 806.680 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.300 0.000 813.580 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 820.200 0.000 820.480 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 826.640 0.000 826.920 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 833.540 0.000 833.820 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.980 0.000 840.260 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.880 0.000 295.160 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.880 0.000 847.160 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 853.780 0.000 854.060 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.220 0.000 860.500 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 867.120 0.000 867.400 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 874.020 0.000 874.300 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.460 0.000 880.740 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 887.360 0.000 887.640 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 894.260 0.000 894.540 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 900.700 0.000 900.980 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.600 0.000 907.880 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 301.320 0.000 301.600 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.900 0.000 243.180 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 916.340 0.000 916.620 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 923.240 0.000 923.520 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.140 0.000 930.420 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.580 0.000 936.860 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 943.480 0.000 943.760 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.380 0.000 950.660 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.820 0.000 957.100 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 963.720 0.000 964.000 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 970.160 0.000 970.440 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.060 0.000 977.340 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.520 0.000 310.800 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.960 0.000 984.240 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.400 0.000 990.680 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 997.300 0.000 997.580 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1004.200 0.000 1004.480 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.640 0.000 1010.920 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1017.540 0.000 1017.820 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.440 0.000 1024.720 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.880 0.000 1031.160 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.780 0.000 1038.060 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.680 0.000 1044.960 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 317.420 0.000 317.700 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1051.120 0.000 1051.400 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.020 0.000 1058.300 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.460 0.000 1064.740 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1071.360 0.000 1071.640 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1078.260 0.000 1078.540 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.700 0.000 1084.980 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1091.600 0.000 1091.880 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.500 0.000 1098.780 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 323.860 0.000 324.140 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.760 0.000 331.040 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.200 0.000 337.480 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.100 0.000 344.380 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.000 0.000 351.280 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.440 0.000 357.720 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 364.340 0.000 364.620 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.240 0.000 371.520 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.800 0.000 250.080 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.680 0.000 377.960 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.580 0.000 384.860 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.480 0.000 391.760 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.920 0.000 398.200 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 404.820 0.000 405.100 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 411.260 0.000 411.540 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.160 0.000 418.440 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.060 0.000 425.340 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.500 0.000 431.780 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.400 0.000 438.680 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.700 0.000 256.980 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 445.300 0.000 445.580 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.740 0.000 452.020 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 458.640 0.000 458.920 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.540 0.000 465.820 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.980 0.000 472.260 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.880 0.000 479.160 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 485.320 0.000 485.600 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.220 0.000 492.500 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.120 0.000 499.400 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 505.560 0.000 505.840 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.140 0.000 263.420 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 512.460 0.000 512.740 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 519.360 0.000 519.640 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.800 0.000 526.080 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 532.700 0.000 532.980 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 539.600 0.000 539.880 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.040 0.000 546.320 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.940 0.000 553.220 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 559.840 0.000 560.120 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 566.280 0.000 566.560 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.180 0.000 573.460 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.040 0.000 270.320 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.620 0.000 579.900 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 586.520 0.000 586.800 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 593.420 0.000 593.700 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.860 0.000 600.140 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 606.760 0.000 607.040 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 613.660 0.000 613.940 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.100 0.000 620.380 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.000 0.000 627.280 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 633.900 0.000 634.180 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.340 0.000 640.620 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.940 0.000 277.220 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 647.240 0.000 647.520 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.680 0.000 653.960 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 660.580 0.000 660.860 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 667.480 0.000 667.760 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.920 0.000 674.200 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.820 0.000 681.100 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.720 0.000 688.000 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 694.160 0.000 694.440 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 701.060 0.000 701.340 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.960 0.000 708.240 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.380 0.000 283.660 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.400 0.000 714.680 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 721.300 0.000 721.580 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.740 0.000 728.020 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.640 0.000 734.920 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 741.540 0.000 741.820 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 747.980 0.000 748.260 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.880 0.000 755.160 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.780 0.000 762.060 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 768.220 0.000 768.500 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.120 0.000 775.400 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.280 0.000 290.560 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.020 0.000 782.300 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.460 0.000 788.740 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 795.360 0.000 795.640 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 802.260 0.000 802.540 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 808.700 0.000 808.980 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 815.600 0.000 815.880 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.040 0.000 822.320 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 828.940 0.000 829.220 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.840 0.000 836.120 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 842.280 0.000 842.560 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 297.180 0.000 297.460 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 849.180 0.000 849.460 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 856.080 0.000 856.360 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.520 0.000 862.800 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.420 0.000 869.700 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.320 0.000 876.600 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.760 0.000 883.040 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 889.660 0.000 889.940 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.100 0.000 896.380 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.000 0.000 903.280 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 909.900 0.000 910.180 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.620 0.000 303.900 4.000 ;
    END
  END la_oen[9]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 14.320 1099.930 14.920 ;
    END
  END one
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.940 0.000 1.220 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.780 0.000 3.060 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.080 0.000 5.360 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.280 0.000 14.560 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.640 0.000 90.920 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.080 0.000 97.360 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.880 0.000 111.160 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.320 0.000 117.600 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.220 0.000 124.500 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.120 0.000 131.400 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.560 0.000 137.840 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.460 0.000 144.740 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.900 0.000 151.180 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.020 0.000 23.300 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.800 0.000 158.080 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.700 0.000 164.980 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.040 0.000 178.320 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.940 0.000 185.220 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.380 0.000 191.660 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.280 0.000 198.560 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 205.180 0.000 205.460 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.620 0.000 211.900 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.520 0.000 218.800 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.220 0.000 32.500 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.960 0.000 225.240 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.860 0.000 232.140 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.960 0.000 41.240 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.160 0.000 50.440 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.600 0.000 56.880 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.500 0.000 63.780 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.400 0.000 70.680 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.840 0.000 77.120 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.740 0.000 84.020 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.380 0.000 7.660 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.580 0.000 16.860 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.940 0.000 93.220 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.380 0.000 99.660 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.280 0.000 106.560 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.720 0.000 113.000 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.620 0.000 119.900 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.520 0.000 126.800 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.960 0.000 133.240 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.860 0.000 140.140 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 146.760 0.000 147.040 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.200 0.000 153.480 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 25.320 0.000 25.600 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.100 0.000 160.380 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 167.000 0.000 167.280 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.440 0.000 173.720 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.340 0.000 180.620 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.240 0.000 187.520 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.680 0.000 193.960 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.580 0.000 200.860 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.020 0.000 207.300 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.920 0.000 214.200 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.820 0.000 221.100 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.520 0.000 34.800 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.260 0.000 227.540 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 234.160 0.000 234.440 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.260 0.000 43.540 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.460 0.000 52.740 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.900 0.000 59.180 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.800 0.000 66.080 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.700 0.000 72.980 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.140 0.000 79.420 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 86.040 0.000 86.320 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.880 0.000 19.160 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.780 0.000 95.060 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.680 0.000 101.960 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.580 0.000 108.860 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.020 0.000 115.300 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.920 0.000 122.200 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.820 0.000 129.100 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 135.260 0.000 135.540 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.160 0.000 142.440 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.060 0.000 149.340 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.500 0.000 155.780 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.620 0.000 27.900 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.400 0.000 162.680 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.840 0.000 169.120 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.740 0.000 176.020 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 182.640 0.000 182.920 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 189.080 0.000 189.360 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.980 0.000 196.260 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 202.880 0.000 203.160 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 209.320 0.000 209.600 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 216.220 0.000 216.500 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 223.120 0.000 223.400 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.820 0.000 37.100 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.560 0.000 229.840 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 236.460 0.000 236.740 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.560 0.000 45.840 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 54.760 0.000 55.040 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.200 0.000 61.480 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.100 0.000 68.380 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.000 0.000 75.280 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.440 0.000 81.720 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.340 0.000 88.620 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 20.720 0.000 21.000 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.920 0.000 30.200 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 38.660 0.000 38.940 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.860 0.000 48.140 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.680 0.000 9.960 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 4.000 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1095.930 4.800 1099.930 5.400 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.970 10.640 22.570 1088.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.770 10.640 99.370 1088.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.450 10.795 1094.270 1088.085 ;
      LAYER met1 ;
        RECT 0.000 10.640 1096.500 1095.780 ;
      LAYER met2 ;
        RECT 0.030 1095.720 4.800 1096.000 ;
        RECT 5.640 1095.720 14.920 1096.000 ;
        RECT 15.760 1095.720 25.500 1096.000 ;
        RECT 26.340 1095.720 35.620 1096.000 ;
        RECT 36.460 1095.720 46.200 1096.000 ;
        RECT 47.040 1095.720 56.320 1096.000 ;
        RECT 57.160 1095.720 66.900 1096.000 ;
        RECT 67.740 1095.720 77.020 1096.000 ;
        RECT 77.860 1095.720 87.600 1096.000 ;
        RECT 88.440 1095.720 98.180 1096.000 ;
        RECT 99.020 1095.720 108.300 1096.000 ;
        RECT 109.140 1095.720 118.880 1096.000 ;
        RECT 119.720 1095.720 129.000 1096.000 ;
        RECT 129.840 1095.720 139.580 1096.000 ;
        RECT 140.420 1095.720 149.700 1096.000 ;
        RECT 150.540 1095.720 160.280 1096.000 ;
        RECT 161.120 1095.720 170.400 1096.000 ;
        RECT 171.240 1095.720 180.980 1096.000 ;
        RECT 181.820 1095.720 191.560 1096.000 ;
        RECT 192.400 1095.720 201.680 1096.000 ;
        RECT 202.520 1095.720 212.260 1096.000 ;
        RECT 213.100 1095.720 222.380 1096.000 ;
        RECT 223.220 1095.720 232.960 1096.000 ;
        RECT 233.800 1095.720 243.080 1096.000 ;
        RECT 243.920 1095.720 253.660 1096.000 ;
        RECT 254.500 1095.720 263.780 1096.000 ;
        RECT 264.620 1095.720 274.360 1096.000 ;
        RECT 275.200 1095.720 284.940 1096.000 ;
        RECT 285.780 1095.720 295.060 1096.000 ;
        RECT 295.900 1095.720 305.640 1096.000 ;
        RECT 306.480 1095.720 315.760 1096.000 ;
        RECT 316.600 1095.720 326.340 1096.000 ;
        RECT 327.180 1095.720 336.460 1096.000 ;
        RECT 337.300 1095.720 347.040 1096.000 ;
        RECT 347.880 1095.720 357.160 1096.000 ;
        RECT 358.000 1095.720 367.740 1096.000 ;
        RECT 368.580 1095.720 378.320 1096.000 ;
        RECT 379.160 1095.720 388.440 1096.000 ;
        RECT 389.280 1095.720 399.020 1096.000 ;
        RECT 399.860 1095.720 409.140 1096.000 ;
        RECT 409.980 1095.720 419.720 1096.000 ;
        RECT 420.560 1095.720 429.840 1096.000 ;
        RECT 430.680 1095.720 440.420 1096.000 ;
        RECT 441.260 1095.720 450.540 1096.000 ;
        RECT 451.380 1095.720 461.120 1096.000 ;
        RECT 461.960 1095.720 471.700 1096.000 ;
        RECT 472.540 1095.720 481.820 1096.000 ;
        RECT 482.660 1095.720 492.400 1096.000 ;
        RECT 493.240 1095.720 502.520 1096.000 ;
        RECT 503.360 1095.720 513.100 1096.000 ;
        RECT 513.940 1095.720 523.220 1096.000 ;
        RECT 524.060 1095.720 533.800 1096.000 ;
        RECT 534.640 1095.720 543.920 1096.000 ;
        RECT 544.760 1095.720 554.500 1096.000 ;
        RECT 555.340 1095.720 565.080 1096.000 ;
        RECT 565.920 1095.720 575.200 1096.000 ;
        RECT 576.040 1095.720 585.780 1096.000 ;
        RECT 586.620 1095.720 595.900 1096.000 ;
        RECT 596.740 1095.720 606.480 1096.000 ;
        RECT 607.320 1095.720 616.600 1096.000 ;
        RECT 617.440 1095.720 627.180 1096.000 ;
        RECT 628.020 1095.720 637.300 1096.000 ;
        RECT 638.140 1095.720 647.880 1096.000 ;
        RECT 648.720 1095.720 658.460 1096.000 ;
        RECT 659.300 1095.720 668.580 1096.000 ;
        RECT 669.420 1095.720 679.160 1096.000 ;
        RECT 680.000 1095.720 689.280 1096.000 ;
        RECT 690.120 1095.720 699.860 1096.000 ;
        RECT 700.700 1095.720 709.980 1096.000 ;
        RECT 710.820 1095.720 720.560 1096.000 ;
        RECT 721.400 1095.720 730.680 1096.000 ;
        RECT 731.520 1095.720 741.260 1096.000 ;
        RECT 742.100 1095.720 751.840 1096.000 ;
        RECT 752.680 1095.720 761.960 1096.000 ;
        RECT 762.800 1095.720 772.540 1096.000 ;
        RECT 773.380 1095.720 782.660 1096.000 ;
        RECT 783.500 1095.720 793.240 1096.000 ;
        RECT 794.080 1095.720 803.360 1096.000 ;
        RECT 804.200 1095.720 813.940 1096.000 ;
        RECT 814.780 1095.720 824.060 1096.000 ;
        RECT 824.900 1095.720 834.640 1096.000 ;
        RECT 835.480 1095.720 845.220 1096.000 ;
        RECT 846.060 1095.720 855.340 1096.000 ;
        RECT 856.180 1095.720 865.920 1096.000 ;
        RECT 866.760 1095.720 876.040 1096.000 ;
        RECT 876.880 1095.720 886.620 1096.000 ;
        RECT 887.460 1095.720 896.740 1096.000 ;
        RECT 897.580 1095.720 907.320 1096.000 ;
        RECT 908.160 1095.720 917.440 1096.000 ;
        RECT 918.280 1095.720 928.020 1096.000 ;
        RECT 928.860 1095.720 938.600 1096.000 ;
        RECT 939.440 1095.720 948.720 1096.000 ;
        RECT 949.560 1095.720 959.300 1096.000 ;
        RECT 960.140 1095.720 969.420 1096.000 ;
        RECT 970.260 1095.720 980.000 1096.000 ;
        RECT 980.840 1095.720 990.120 1096.000 ;
        RECT 990.960 1095.720 1000.700 1096.000 ;
        RECT 1001.540 1095.720 1010.820 1096.000 ;
        RECT 1011.660 1095.720 1021.400 1096.000 ;
        RECT 1022.240 1095.720 1031.980 1096.000 ;
        RECT 1032.820 1095.720 1042.100 1096.000 ;
        RECT 1042.940 1095.720 1052.680 1096.000 ;
        RECT 1053.520 1095.720 1062.800 1096.000 ;
        RECT 1063.640 1095.720 1073.380 1096.000 ;
        RECT 1074.220 1095.720 1083.500 1096.000 ;
        RECT 1084.340 1095.720 1094.080 1096.000 ;
        RECT 1094.920 1095.720 1096.470 1096.000 ;
        RECT 0.030 4.280 1096.470 1095.720 ;
        RECT 0.030 4.000 0.660 4.280 ;
        RECT 1.500 4.000 2.500 4.280 ;
        RECT 3.340 4.000 4.800 4.280 ;
        RECT 5.640 4.000 7.100 4.280 ;
        RECT 7.940 4.000 9.400 4.280 ;
        RECT 10.240 4.000 11.700 4.280 ;
        RECT 12.540 4.000 14.000 4.280 ;
        RECT 14.840 4.000 16.300 4.280 ;
        RECT 17.140 4.000 18.600 4.280 ;
        RECT 19.440 4.000 20.440 4.280 ;
        RECT 21.280 4.000 22.740 4.280 ;
        RECT 23.580 4.000 25.040 4.280 ;
        RECT 25.880 4.000 27.340 4.280 ;
        RECT 28.180 4.000 29.640 4.280 ;
        RECT 30.480 4.000 31.940 4.280 ;
        RECT 32.780 4.000 34.240 4.280 ;
        RECT 35.080 4.000 36.540 4.280 ;
        RECT 37.380 4.000 38.380 4.280 ;
        RECT 39.220 4.000 40.680 4.280 ;
        RECT 41.520 4.000 42.980 4.280 ;
        RECT 43.820 4.000 45.280 4.280 ;
        RECT 46.120 4.000 47.580 4.280 ;
        RECT 48.420 4.000 49.880 4.280 ;
        RECT 50.720 4.000 52.180 4.280 ;
        RECT 53.020 4.000 54.480 4.280 ;
        RECT 55.320 4.000 56.320 4.280 ;
        RECT 57.160 4.000 58.620 4.280 ;
        RECT 59.460 4.000 60.920 4.280 ;
        RECT 61.760 4.000 63.220 4.280 ;
        RECT 64.060 4.000 65.520 4.280 ;
        RECT 66.360 4.000 67.820 4.280 ;
        RECT 68.660 4.000 70.120 4.280 ;
        RECT 70.960 4.000 72.420 4.280 ;
        RECT 73.260 4.000 74.720 4.280 ;
        RECT 75.560 4.000 76.560 4.280 ;
        RECT 77.400 4.000 78.860 4.280 ;
        RECT 79.700 4.000 81.160 4.280 ;
        RECT 82.000 4.000 83.460 4.280 ;
        RECT 84.300 4.000 85.760 4.280 ;
        RECT 86.600 4.000 88.060 4.280 ;
        RECT 88.900 4.000 90.360 4.280 ;
        RECT 91.200 4.000 92.660 4.280 ;
        RECT 93.500 4.000 94.500 4.280 ;
        RECT 95.340 4.000 96.800 4.280 ;
        RECT 97.640 4.000 99.100 4.280 ;
        RECT 99.940 4.000 101.400 4.280 ;
        RECT 102.240 4.000 103.700 4.280 ;
        RECT 104.540 4.000 106.000 4.280 ;
        RECT 106.840 4.000 108.300 4.280 ;
        RECT 109.140 4.000 110.600 4.280 ;
        RECT 111.440 4.000 112.440 4.280 ;
        RECT 113.280 4.000 114.740 4.280 ;
        RECT 115.580 4.000 117.040 4.280 ;
        RECT 117.880 4.000 119.340 4.280 ;
        RECT 120.180 4.000 121.640 4.280 ;
        RECT 122.480 4.000 123.940 4.280 ;
        RECT 124.780 4.000 126.240 4.280 ;
        RECT 127.080 4.000 128.540 4.280 ;
        RECT 129.380 4.000 130.840 4.280 ;
        RECT 131.680 4.000 132.680 4.280 ;
        RECT 133.520 4.000 134.980 4.280 ;
        RECT 135.820 4.000 137.280 4.280 ;
        RECT 138.120 4.000 139.580 4.280 ;
        RECT 140.420 4.000 141.880 4.280 ;
        RECT 142.720 4.000 144.180 4.280 ;
        RECT 145.020 4.000 146.480 4.280 ;
        RECT 147.320 4.000 148.780 4.280 ;
        RECT 149.620 4.000 150.620 4.280 ;
        RECT 151.460 4.000 152.920 4.280 ;
        RECT 153.760 4.000 155.220 4.280 ;
        RECT 156.060 4.000 157.520 4.280 ;
        RECT 158.360 4.000 159.820 4.280 ;
        RECT 160.660 4.000 162.120 4.280 ;
        RECT 162.960 4.000 164.420 4.280 ;
        RECT 165.260 4.000 166.720 4.280 ;
        RECT 167.560 4.000 168.560 4.280 ;
        RECT 169.400 4.000 170.860 4.280 ;
        RECT 171.700 4.000 173.160 4.280 ;
        RECT 174.000 4.000 175.460 4.280 ;
        RECT 176.300 4.000 177.760 4.280 ;
        RECT 178.600 4.000 180.060 4.280 ;
        RECT 180.900 4.000 182.360 4.280 ;
        RECT 183.200 4.000 184.660 4.280 ;
        RECT 185.500 4.000 186.960 4.280 ;
        RECT 187.800 4.000 188.800 4.280 ;
        RECT 189.640 4.000 191.100 4.280 ;
        RECT 191.940 4.000 193.400 4.280 ;
        RECT 194.240 4.000 195.700 4.280 ;
        RECT 196.540 4.000 198.000 4.280 ;
        RECT 198.840 4.000 200.300 4.280 ;
        RECT 201.140 4.000 202.600 4.280 ;
        RECT 203.440 4.000 204.900 4.280 ;
        RECT 205.740 4.000 206.740 4.280 ;
        RECT 207.580 4.000 209.040 4.280 ;
        RECT 209.880 4.000 211.340 4.280 ;
        RECT 212.180 4.000 213.640 4.280 ;
        RECT 214.480 4.000 215.940 4.280 ;
        RECT 216.780 4.000 218.240 4.280 ;
        RECT 219.080 4.000 220.540 4.280 ;
        RECT 221.380 4.000 222.840 4.280 ;
        RECT 223.680 4.000 224.680 4.280 ;
        RECT 225.520 4.000 226.980 4.280 ;
        RECT 227.820 4.000 229.280 4.280 ;
        RECT 230.120 4.000 231.580 4.280 ;
        RECT 232.420 4.000 233.880 4.280 ;
        RECT 234.720 4.000 236.180 4.280 ;
        RECT 237.020 4.000 238.480 4.280 ;
        RECT 239.320 4.000 240.780 4.280 ;
        RECT 241.620 4.000 242.620 4.280 ;
        RECT 243.460 4.000 244.920 4.280 ;
        RECT 245.760 4.000 247.220 4.280 ;
        RECT 248.060 4.000 249.520 4.280 ;
        RECT 250.360 4.000 251.820 4.280 ;
        RECT 252.660 4.000 254.120 4.280 ;
        RECT 254.960 4.000 256.420 4.280 ;
        RECT 257.260 4.000 258.720 4.280 ;
        RECT 259.560 4.000 261.020 4.280 ;
        RECT 261.860 4.000 262.860 4.280 ;
        RECT 263.700 4.000 265.160 4.280 ;
        RECT 266.000 4.000 267.460 4.280 ;
        RECT 268.300 4.000 269.760 4.280 ;
        RECT 270.600 4.000 272.060 4.280 ;
        RECT 272.900 4.000 274.360 4.280 ;
        RECT 275.200 4.000 276.660 4.280 ;
        RECT 277.500 4.000 278.960 4.280 ;
        RECT 279.800 4.000 280.800 4.280 ;
        RECT 281.640 4.000 283.100 4.280 ;
        RECT 283.940 4.000 285.400 4.280 ;
        RECT 286.240 4.000 287.700 4.280 ;
        RECT 288.540 4.000 290.000 4.280 ;
        RECT 290.840 4.000 292.300 4.280 ;
        RECT 293.140 4.000 294.600 4.280 ;
        RECT 295.440 4.000 296.900 4.280 ;
        RECT 297.740 4.000 298.740 4.280 ;
        RECT 299.580 4.000 301.040 4.280 ;
        RECT 301.880 4.000 303.340 4.280 ;
        RECT 304.180 4.000 305.640 4.280 ;
        RECT 306.480 4.000 307.940 4.280 ;
        RECT 308.780 4.000 310.240 4.280 ;
        RECT 311.080 4.000 312.540 4.280 ;
        RECT 313.380 4.000 314.840 4.280 ;
        RECT 315.680 4.000 317.140 4.280 ;
        RECT 317.980 4.000 318.980 4.280 ;
        RECT 319.820 4.000 321.280 4.280 ;
        RECT 322.120 4.000 323.580 4.280 ;
        RECT 324.420 4.000 325.880 4.280 ;
        RECT 326.720 4.000 328.180 4.280 ;
        RECT 329.020 4.000 330.480 4.280 ;
        RECT 331.320 4.000 332.780 4.280 ;
        RECT 333.620 4.000 335.080 4.280 ;
        RECT 335.920 4.000 336.920 4.280 ;
        RECT 337.760 4.000 339.220 4.280 ;
        RECT 340.060 4.000 341.520 4.280 ;
        RECT 342.360 4.000 343.820 4.280 ;
        RECT 344.660 4.000 346.120 4.280 ;
        RECT 346.960 4.000 348.420 4.280 ;
        RECT 349.260 4.000 350.720 4.280 ;
        RECT 351.560 4.000 353.020 4.280 ;
        RECT 353.860 4.000 354.860 4.280 ;
        RECT 355.700 4.000 357.160 4.280 ;
        RECT 358.000 4.000 359.460 4.280 ;
        RECT 360.300 4.000 361.760 4.280 ;
        RECT 362.600 4.000 364.060 4.280 ;
        RECT 364.900 4.000 366.360 4.280 ;
        RECT 367.200 4.000 368.660 4.280 ;
        RECT 369.500 4.000 370.960 4.280 ;
        RECT 371.800 4.000 373.260 4.280 ;
        RECT 374.100 4.000 375.100 4.280 ;
        RECT 375.940 4.000 377.400 4.280 ;
        RECT 378.240 4.000 379.700 4.280 ;
        RECT 380.540 4.000 382.000 4.280 ;
        RECT 382.840 4.000 384.300 4.280 ;
        RECT 385.140 4.000 386.600 4.280 ;
        RECT 387.440 4.000 388.900 4.280 ;
        RECT 389.740 4.000 391.200 4.280 ;
        RECT 392.040 4.000 393.040 4.280 ;
        RECT 393.880 4.000 395.340 4.280 ;
        RECT 396.180 4.000 397.640 4.280 ;
        RECT 398.480 4.000 399.940 4.280 ;
        RECT 400.780 4.000 402.240 4.280 ;
        RECT 403.080 4.000 404.540 4.280 ;
        RECT 405.380 4.000 406.840 4.280 ;
        RECT 407.680 4.000 409.140 4.280 ;
        RECT 409.980 4.000 410.980 4.280 ;
        RECT 411.820 4.000 413.280 4.280 ;
        RECT 414.120 4.000 415.580 4.280 ;
        RECT 416.420 4.000 417.880 4.280 ;
        RECT 418.720 4.000 420.180 4.280 ;
        RECT 421.020 4.000 422.480 4.280 ;
        RECT 423.320 4.000 424.780 4.280 ;
        RECT 425.620 4.000 427.080 4.280 ;
        RECT 427.920 4.000 429.380 4.280 ;
        RECT 430.220 4.000 431.220 4.280 ;
        RECT 432.060 4.000 433.520 4.280 ;
        RECT 434.360 4.000 435.820 4.280 ;
        RECT 436.660 4.000 438.120 4.280 ;
        RECT 438.960 4.000 440.420 4.280 ;
        RECT 441.260 4.000 442.720 4.280 ;
        RECT 443.560 4.000 445.020 4.280 ;
        RECT 445.860 4.000 447.320 4.280 ;
        RECT 448.160 4.000 449.160 4.280 ;
        RECT 450.000 4.000 451.460 4.280 ;
        RECT 452.300 4.000 453.760 4.280 ;
        RECT 454.600 4.000 456.060 4.280 ;
        RECT 456.900 4.000 458.360 4.280 ;
        RECT 459.200 4.000 460.660 4.280 ;
        RECT 461.500 4.000 462.960 4.280 ;
        RECT 463.800 4.000 465.260 4.280 ;
        RECT 466.100 4.000 467.100 4.280 ;
        RECT 467.940 4.000 469.400 4.280 ;
        RECT 470.240 4.000 471.700 4.280 ;
        RECT 472.540 4.000 474.000 4.280 ;
        RECT 474.840 4.000 476.300 4.280 ;
        RECT 477.140 4.000 478.600 4.280 ;
        RECT 479.440 4.000 480.900 4.280 ;
        RECT 481.740 4.000 483.200 4.280 ;
        RECT 484.040 4.000 485.040 4.280 ;
        RECT 485.880 4.000 487.340 4.280 ;
        RECT 488.180 4.000 489.640 4.280 ;
        RECT 490.480 4.000 491.940 4.280 ;
        RECT 492.780 4.000 494.240 4.280 ;
        RECT 495.080 4.000 496.540 4.280 ;
        RECT 497.380 4.000 498.840 4.280 ;
        RECT 499.680 4.000 501.140 4.280 ;
        RECT 501.980 4.000 503.440 4.280 ;
        RECT 504.280 4.000 505.280 4.280 ;
        RECT 506.120 4.000 507.580 4.280 ;
        RECT 508.420 4.000 509.880 4.280 ;
        RECT 510.720 4.000 512.180 4.280 ;
        RECT 513.020 4.000 514.480 4.280 ;
        RECT 515.320 4.000 516.780 4.280 ;
        RECT 517.620 4.000 519.080 4.280 ;
        RECT 519.920 4.000 521.380 4.280 ;
        RECT 522.220 4.000 523.220 4.280 ;
        RECT 524.060 4.000 525.520 4.280 ;
        RECT 526.360 4.000 527.820 4.280 ;
        RECT 528.660 4.000 530.120 4.280 ;
        RECT 530.960 4.000 532.420 4.280 ;
        RECT 533.260 4.000 534.720 4.280 ;
        RECT 535.560 4.000 537.020 4.280 ;
        RECT 537.860 4.000 539.320 4.280 ;
        RECT 540.160 4.000 541.160 4.280 ;
        RECT 542.000 4.000 543.460 4.280 ;
        RECT 544.300 4.000 545.760 4.280 ;
        RECT 546.600 4.000 548.060 4.280 ;
        RECT 548.900 4.000 550.360 4.280 ;
        RECT 551.200 4.000 552.660 4.280 ;
        RECT 553.500 4.000 554.960 4.280 ;
        RECT 555.800 4.000 557.260 4.280 ;
        RECT 558.100 4.000 559.560 4.280 ;
        RECT 560.400 4.000 561.400 4.280 ;
        RECT 562.240 4.000 563.700 4.280 ;
        RECT 564.540 4.000 566.000 4.280 ;
        RECT 566.840 4.000 568.300 4.280 ;
        RECT 569.140 4.000 570.600 4.280 ;
        RECT 571.440 4.000 572.900 4.280 ;
        RECT 573.740 4.000 575.200 4.280 ;
        RECT 576.040 4.000 577.500 4.280 ;
        RECT 578.340 4.000 579.340 4.280 ;
        RECT 580.180 4.000 581.640 4.280 ;
        RECT 582.480 4.000 583.940 4.280 ;
        RECT 584.780 4.000 586.240 4.280 ;
        RECT 587.080 4.000 588.540 4.280 ;
        RECT 589.380 4.000 590.840 4.280 ;
        RECT 591.680 4.000 593.140 4.280 ;
        RECT 593.980 4.000 595.440 4.280 ;
        RECT 596.280 4.000 597.280 4.280 ;
        RECT 598.120 4.000 599.580 4.280 ;
        RECT 600.420 4.000 601.880 4.280 ;
        RECT 602.720 4.000 604.180 4.280 ;
        RECT 605.020 4.000 606.480 4.280 ;
        RECT 607.320 4.000 608.780 4.280 ;
        RECT 609.620 4.000 611.080 4.280 ;
        RECT 611.920 4.000 613.380 4.280 ;
        RECT 614.220 4.000 615.680 4.280 ;
        RECT 616.520 4.000 617.520 4.280 ;
        RECT 618.360 4.000 619.820 4.280 ;
        RECT 620.660 4.000 622.120 4.280 ;
        RECT 622.960 4.000 624.420 4.280 ;
        RECT 625.260 4.000 626.720 4.280 ;
        RECT 627.560 4.000 629.020 4.280 ;
        RECT 629.860 4.000 631.320 4.280 ;
        RECT 632.160 4.000 633.620 4.280 ;
        RECT 634.460 4.000 635.460 4.280 ;
        RECT 636.300 4.000 637.760 4.280 ;
        RECT 638.600 4.000 640.060 4.280 ;
        RECT 640.900 4.000 642.360 4.280 ;
        RECT 643.200 4.000 644.660 4.280 ;
        RECT 645.500 4.000 646.960 4.280 ;
        RECT 647.800 4.000 649.260 4.280 ;
        RECT 650.100 4.000 651.560 4.280 ;
        RECT 652.400 4.000 653.400 4.280 ;
        RECT 654.240 4.000 655.700 4.280 ;
        RECT 656.540 4.000 658.000 4.280 ;
        RECT 658.840 4.000 660.300 4.280 ;
        RECT 661.140 4.000 662.600 4.280 ;
        RECT 663.440 4.000 664.900 4.280 ;
        RECT 665.740 4.000 667.200 4.280 ;
        RECT 668.040 4.000 669.500 4.280 ;
        RECT 670.340 4.000 671.340 4.280 ;
        RECT 672.180 4.000 673.640 4.280 ;
        RECT 674.480 4.000 675.940 4.280 ;
        RECT 676.780 4.000 678.240 4.280 ;
        RECT 679.080 4.000 680.540 4.280 ;
        RECT 681.380 4.000 682.840 4.280 ;
        RECT 683.680 4.000 685.140 4.280 ;
        RECT 685.980 4.000 687.440 4.280 ;
        RECT 688.280 4.000 689.740 4.280 ;
        RECT 690.580 4.000 691.580 4.280 ;
        RECT 692.420 4.000 693.880 4.280 ;
        RECT 694.720 4.000 696.180 4.280 ;
        RECT 697.020 4.000 698.480 4.280 ;
        RECT 699.320 4.000 700.780 4.280 ;
        RECT 701.620 4.000 703.080 4.280 ;
        RECT 703.920 4.000 705.380 4.280 ;
        RECT 706.220 4.000 707.680 4.280 ;
        RECT 708.520 4.000 709.520 4.280 ;
        RECT 710.360 4.000 711.820 4.280 ;
        RECT 712.660 4.000 714.120 4.280 ;
        RECT 714.960 4.000 716.420 4.280 ;
        RECT 717.260 4.000 718.720 4.280 ;
        RECT 719.560 4.000 721.020 4.280 ;
        RECT 721.860 4.000 723.320 4.280 ;
        RECT 724.160 4.000 725.620 4.280 ;
        RECT 726.460 4.000 727.460 4.280 ;
        RECT 728.300 4.000 729.760 4.280 ;
        RECT 730.600 4.000 732.060 4.280 ;
        RECT 732.900 4.000 734.360 4.280 ;
        RECT 735.200 4.000 736.660 4.280 ;
        RECT 737.500 4.000 738.960 4.280 ;
        RECT 739.800 4.000 741.260 4.280 ;
        RECT 742.100 4.000 743.560 4.280 ;
        RECT 744.400 4.000 745.860 4.280 ;
        RECT 746.700 4.000 747.700 4.280 ;
        RECT 748.540 4.000 750.000 4.280 ;
        RECT 750.840 4.000 752.300 4.280 ;
        RECT 753.140 4.000 754.600 4.280 ;
        RECT 755.440 4.000 756.900 4.280 ;
        RECT 757.740 4.000 759.200 4.280 ;
        RECT 760.040 4.000 761.500 4.280 ;
        RECT 762.340 4.000 763.800 4.280 ;
        RECT 764.640 4.000 765.640 4.280 ;
        RECT 766.480 4.000 767.940 4.280 ;
        RECT 768.780 4.000 770.240 4.280 ;
        RECT 771.080 4.000 772.540 4.280 ;
        RECT 773.380 4.000 774.840 4.280 ;
        RECT 775.680 4.000 777.140 4.280 ;
        RECT 777.980 4.000 779.440 4.280 ;
        RECT 780.280 4.000 781.740 4.280 ;
        RECT 782.580 4.000 783.580 4.280 ;
        RECT 784.420 4.000 785.880 4.280 ;
        RECT 786.720 4.000 788.180 4.280 ;
        RECT 789.020 4.000 790.480 4.280 ;
        RECT 791.320 4.000 792.780 4.280 ;
        RECT 793.620 4.000 795.080 4.280 ;
        RECT 795.920 4.000 797.380 4.280 ;
        RECT 798.220 4.000 799.680 4.280 ;
        RECT 800.520 4.000 801.980 4.280 ;
        RECT 802.820 4.000 803.820 4.280 ;
        RECT 804.660 4.000 806.120 4.280 ;
        RECT 806.960 4.000 808.420 4.280 ;
        RECT 809.260 4.000 810.720 4.280 ;
        RECT 811.560 4.000 813.020 4.280 ;
        RECT 813.860 4.000 815.320 4.280 ;
        RECT 816.160 4.000 817.620 4.280 ;
        RECT 818.460 4.000 819.920 4.280 ;
        RECT 820.760 4.000 821.760 4.280 ;
        RECT 822.600 4.000 824.060 4.280 ;
        RECT 824.900 4.000 826.360 4.280 ;
        RECT 827.200 4.000 828.660 4.280 ;
        RECT 829.500 4.000 830.960 4.280 ;
        RECT 831.800 4.000 833.260 4.280 ;
        RECT 834.100 4.000 835.560 4.280 ;
        RECT 836.400 4.000 837.860 4.280 ;
        RECT 838.700 4.000 839.700 4.280 ;
        RECT 840.540 4.000 842.000 4.280 ;
        RECT 842.840 4.000 844.300 4.280 ;
        RECT 845.140 4.000 846.600 4.280 ;
        RECT 847.440 4.000 848.900 4.280 ;
        RECT 849.740 4.000 851.200 4.280 ;
        RECT 852.040 4.000 853.500 4.280 ;
        RECT 854.340 4.000 855.800 4.280 ;
        RECT 856.640 4.000 858.100 4.280 ;
        RECT 858.940 4.000 859.940 4.280 ;
        RECT 860.780 4.000 862.240 4.280 ;
        RECT 863.080 4.000 864.540 4.280 ;
        RECT 865.380 4.000 866.840 4.280 ;
        RECT 867.680 4.000 869.140 4.280 ;
        RECT 869.980 4.000 871.440 4.280 ;
        RECT 872.280 4.000 873.740 4.280 ;
        RECT 874.580 4.000 876.040 4.280 ;
        RECT 876.880 4.000 877.880 4.280 ;
        RECT 878.720 4.000 880.180 4.280 ;
        RECT 881.020 4.000 882.480 4.280 ;
        RECT 883.320 4.000 884.780 4.280 ;
        RECT 885.620 4.000 887.080 4.280 ;
        RECT 887.920 4.000 889.380 4.280 ;
        RECT 890.220 4.000 891.680 4.280 ;
        RECT 892.520 4.000 893.980 4.280 ;
        RECT 894.820 4.000 895.820 4.280 ;
        RECT 896.660 4.000 898.120 4.280 ;
        RECT 898.960 4.000 900.420 4.280 ;
        RECT 901.260 4.000 902.720 4.280 ;
        RECT 903.560 4.000 905.020 4.280 ;
        RECT 905.860 4.000 907.320 4.280 ;
        RECT 908.160 4.000 909.620 4.280 ;
        RECT 910.460 4.000 911.920 4.280 ;
        RECT 912.760 4.000 913.760 4.280 ;
        RECT 914.600 4.000 916.060 4.280 ;
        RECT 916.900 4.000 918.360 4.280 ;
        RECT 919.200 4.000 920.660 4.280 ;
        RECT 921.500 4.000 922.960 4.280 ;
        RECT 923.800 4.000 925.260 4.280 ;
        RECT 926.100 4.000 927.560 4.280 ;
        RECT 928.400 4.000 929.860 4.280 ;
        RECT 930.700 4.000 932.160 4.280 ;
        RECT 933.000 4.000 934.000 4.280 ;
        RECT 934.840 4.000 936.300 4.280 ;
        RECT 937.140 4.000 938.600 4.280 ;
        RECT 939.440 4.000 940.900 4.280 ;
        RECT 941.740 4.000 943.200 4.280 ;
        RECT 944.040 4.000 945.500 4.280 ;
        RECT 946.340 4.000 947.800 4.280 ;
        RECT 948.640 4.000 950.100 4.280 ;
        RECT 950.940 4.000 951.940 4.280 ;
        RECT 952.780 4.000 954.240 4.280 ;
        RECT 955.080 4.000 956.540 4.280 ;
        RECT 957.380 4.000 958.840 4.280 ;
        RECT 959.680 4.000 961.140 4.280 ;
        RECT 961.980 4.000 963.440 4.280 ;
        RECT 964.280 4.000 965.740 4.280 ;
        RECT 966.580 4.000 968.040 4.280 ;
        RECT 968.880 4.000 969.880 4.280 ;
        RECT 970.720 4.000 972.180 4.280 ;
        RECT 973.020 4.000 974.480 4.280 ;
        RECT 975.320 4.000 976.780 4.280 ;
        RECT 977.620 4.000 979.080 4.280 ;
        RECT 979.920 4.000 981.380 4.280 ;
        RECT 982.220 4.000 983.680 4.280 ;
        RECT 984.520 4.000 985.980 4.280 ;
        RECT 986.820 4.000 988.280 4.280 ;
        RECT 989.120 4.000 990.120 4.280 ;
        RECT 990.960 4.000 992.420 4.280 ;
        RECT 993.260 4.000 994.720 4.280 ;
        RECT 995.560 4.000 997.020 4.280 ;
        RECT 997.860 4.000 999.320 4.280 ;
        RECT 1000.160 4.000 1001.620 4.280 ;
        RECT 1002.460 4.000 1003.920 4.280 ;
        RECT 1004.760 4.000 1006.220 4.280 ;
        RECT 1007.060 4.000 1008.060 4.280 ;
        RECT 1008.900 4.000 1010.360 4.280 ;
        RECT 1011.200 4.000 1012.660 4.280 ;
        RECT 1013.500 4.000 1014.960 4.280 ;
        RECT 1015.800 4.000 1017.260 4.280 ;
        RECT 1018.100 4.000 1019.560 4.280 ;
        RECT 1020.400 4.000 1021.860 4.280 ;
        RECT 1022.700 4.000 1024.160 4.280 ;
        RECT 1025.000 4.000 1026.000 4.280 ;
        RECT 1026.840 4.000 1028.300 4.280 ;
        RECT 1029.140 4.000 1030.600 4.280 ;
        RECT 1031.440 4.000 1032.900 4.280 ;
        RECT 1033.740 4.000 1035.200 4.280 ;
        RECT 1036.040 4.000 1037.500 4.280 ;
        RECT 1038.340 4.000 1039.800 4.280 ;
        RECT 1040.640 4.000 1042.100 4.280 ;
        RECT 1042.940 4.000 1044.400 4.280 ;
        RECT 1045.240 4.000 1046.240 4.280 ;
        RECT 1047.080 4.000 1048.540 4.280 ;
        RECT 1049.380 4.000 1050.840 4.280 ;
        RECT 1051.680 4.000 1053.140 4.280 ;
        RECT 1053.980 4.000 1055.440 4.280 ;
        RECT 1056.280 4.000 1057.740 4.280 ;
        RECT 1058.580 4.000 1060.040 4.280 ;
        RECT 1060.880 4.000 1062.340 4.280 ;
        RECT 1063.180 4.000 1064.180 4.280 ;
        RECT 1065.020 4.000 1066.480 4.280 ;
        RECT 1067.320 4.000 1068.780 4.280 ;
        RECT 1069.620 4.000 1071.080 4.280 ;
        RECT 1071.920 4.000 1073.380 4.280 ;
        RECT 1074.220 4.000 1075.680 4.280 ;
        RECT 1076.520 4.000 1077.980 4.280 ;
        RECT 1078.820 4.000 1080.280 4.280 ;
        RECT 1081.120 4.000 1082.120 4.280 ;
        RECT 1082.960 4.000 1084.420 4.280 ;
        RECT 1085.260 4.000 1086.720 4.280 ;
        RECT 1087.560 4.000 1089.020 4.280 ;
        RECT 1089.860 4.000 1091.320 4.280 ;
        RECT 1092.160 4.000 1093.620 4.280 ;
        RECT 1094.460 4.000 1095.920 4.280 ;
      LAYER met3 ;
        RECT 0.915 1094.440 1095.530 1095.305 ;
        RECT 0.915 1085.640 1095.930 1094.440 ;
        RECT 0.915 1084.240 1095.530 1085.640 ;
        RECT 0.915 1075.440 1095.930 1084.240 ;
        RECT 0.915 1074.040 1095.530 1075.440 ;
        RECT 0.915 1065.240 1095.930 1074.040 ;
        RECT 0.915 1063.840 1095.530 1065.240 ;
        RECT 0.915 1055.040 1095.930 1063.840 ;
        RECT 0.915 1053.640 1095.530 1055.040 ;
        RECT 0.915 1044.840 1095.930 1053.640 ;
        RECT 0.915 1043.440 1095.530 1044.840 ;
        RECT 0.915 1034.640 1095.930 1043.440 ;
        RECT 0.915 1033.240 1095.530 1034.640 ;
        RECT 0.915 1024.440 1095.930 1033.240 ;
        RECT 0.915 1023.040 1095.530 1024.440 ;
        RECT 0.915 1014.240 1095.930 1023.040 ;
        RECT 0.915 1012.840 1095.530 1014.240 ;
        RECT 0.915 1004.040 1095.930 1012.840 ;
        RECT 0.915 1002.640 1095.530 1004.040 ;
        RECT 0.915 993.840 1095.930 1002.640 ;
        RECT 0.915 992.440 1095.530 993.840 ;
        RECT 0.915 983.640 1095.930 992.440 ;
        RECT 0.915 982.240 1095.530 983.640 ;
        RECT 0.915 973.440 1095.930 982.240 ;
        RECT 0.915 972.040 1095.530 973.440 ;
        RECT 0.915 963.240 1095.930 972.040 ;
        RECT 0.915 961.840 1095.530 963.240 ;
        RECT 0.915 953.040 1095.930 961.840 ;
        RECT 0.915 951.640 1095.530 953.040 ;
        RECT 0.915 942.840 1095.930 951.640 ;
        RECT 0.915 941.440 1095.530 942.840 ;
        RECT 0.915 932.640 1095.930 941.440 ;
        RECT 0.915 931.240 1095.530 932.640 ;
        RECT 0.915 922.440 1095.930 931.240 ;
        RECT 0.915 921.040 1095.530 922.440 ;
        RECT 0.915 912.240 1095.930 921.040 ;
        RECT 0.915 910.840 1095.530 912.240 ;
        RECT 0.915 902.040 1095.930 910.840 ;
        RECT 0.915 900.640 1095.530 902.040 ;
        RECT 0.915 891.840 1095.930 900.640 ;
        RECT 0.915 890.440 1095.530 891.840 ;
        RECT 0.915 881.640 1095.930 890.440 ;
        RECT 0.915 880.240 1095.530 881.640 ;
        RECT 0.915 871.440 1095.930 880.240 ;
        RECT 0.915 870.040 1095.530 871.440 ;
        RECT 0.915 861.240 1095.930 870.040 ;
        RECT 0.915 859.840 1095.530 861.240 ;
        RECT 0.915 851.040 1095.930 859.840 ;
        RECT 0.915 849.640 1095.530 851.040 ;
        RECT 0.915 840.840 1095.930 849.640 ;
        RECT 0.915 839.440 1095.530 840.840 ;
        RECT 0.915 830.640 1095.930 839.440 ;
        RECT 0.915 829.240 1095.530 830.640 ;
        RECT 0.915 820.440 1095.930 829.240 ;
        RECT 0.915 819.040 1095.530 820.440 ;
        RECT 0.915 810.240 1095.930 819.040 ;
        RECT 0.915 808.840 1095.530 810.240 ;
        RECT 0.915 800.040 1095.930 808.840 ;
        RECT 0.915 798.640 1095.530 800.040 ;
        RECT 0.915 789.840 1095.930 798.640 ;
        RECT 0.915 788.440 1095.530 789.840 ;
        RECT 0.915 779.640 1095.930 788.440 ;
        RECT 0.915 778.240 1095.530 779.640 ;
        RECT 0.915 769.440 1095.930 778.240 ;
        RECT 0.915 768.040 1095.530 769.440 ;
        RECT 0.915 759.240 1095.930 768.040 ;
        RECT 0.915 757.840 1095.530 759.240 ;
        RECT 0.915 749.040 1095.930 757.840 ;
        RECT 0.915 747.640 1095.530 749.040 ;
        RECT 0.915 738.840 1095.930 747.640 ;
        RECT 0.915 737.440 1095.530 738.840 ;
        RECT 0.915 728.640 1095.930 737.440 ;
        RECT 0.915 727.240 1095.530 728.640 ;
        RECT 0.915 718.440 1095.930 727.240 ;
        RECT 0.915 717.040 1095.530 718.440 ;
        RECT 0.915 708.240 1095.930 717.040 ;
        RECT 0.915 706.840 1095.530 708.240 ;
        RECT 0.915 698.040 1095.930 706.840 ;
        RECT 0.915 696.640 1095.530 698.040 ;
        RECT 0.915 687.840 1095.930 696.640 ;
        RECT 0.915 686.440 1095.530 687.840 ;
        RECT 0.915 677.640 1095.930 686.440 ;
        RECT 0.915 676.240 1095.530 677.640 ;
        RECT 0.915 667.440 1095.930 676.240 ;
        RECT 0.915 666.040 1095.530 667.440 ;
        RECT 0.915 657.240 1095.930 666.040 ;
        RECT 0.915 655.840 1095.530 657.240 ;
        RECT 0.915 647.040 1095.930 655.840 ;
        RECT 0.915 645.640 1095.530 647.040 ;
        RECT 0.915 636.840 1095.930 645.640 ;
        RECT 0.915 635.440 1095.530 636.840 ;
        RECT 0.915 626.640 1095.930 635.440 ;
        RECT 0.915 625.240 1095.530 626.640 ;
        RECT 0.915 616.440 1095.930 625.240 ;
        RECT 0.915 615.040 1095.530 616.440 ;
        RECT 0.915 606.240 1095.930 615.040 ;
        RECT 0.915 604.840 1095.530 606.240 ;
        RECT 0.915 596.040 1095.930 604.840 ;
        RECT 0.915 594.640 1095.530 596.040 ;
        RECT 0.915 585.840 1095.930 594.640 ;
        RECT 0.915 584.440 1095.530 585.840 ;
        RECT 0.915 575.640 1095.930 584.440 ;
        RECT 0.915 574.240 1095.530 575.640 ;
        RECT 0.915 565.440 1095.930 574.240 ;
        RECT 0.915 564.040 1095.530 565.440 ;
        RECT 0.915 555.920 1095.930 564.040 ;
        RECT 0.915 554.520 1095.530 555.920 ;
        RECT 0.915 545.720 1095.930 554.520 ;
        RECT 0.915 544.320 1095.530 545.720 ;
        RECT 0.915 535.520 1095.930 544.320 ;
        RECT 0.915 534.120 1095.530 535.520 ;
        RECT 0.915 525.320 1095.930 534.120 ;
        RECT 0.915 523.920 1095.530 525.320 ;
        RECT 0.915 515.120 1095.930 523.920 ;
        RECT 0.915 513.720 1095.530 515.120 ;
        RECT 0.915 504.920 1095.930 513.720 ;
        RECT 0.915 503.520 1095.530 504.920 ;
        RECT 0.915 494.720 1095.930 503.520 ;
        RECT 0.915 493.320 1095.530 494.720 ;
        RECT 0.915 484.520 1095.930 493.320 ;
        RECT 0.915 483.120 1095.530 484.520 ;
        RECT 0.915 474.320 1095.930 483.120 ;
        RECT 0.915 472.920 1095.530 474.320 ;
        RECT 0.915 464.120 1095.930 472.920 ;
        RECT 0.915 462.720 1095.530 464.120 ;
        RECT 0.915 453.920 1095.930 462.720 ;
        RECT 0.915 452.520 1095.530 453.920 ;
        RECT 0.915 443.720 1095.930 452.520 ;
        RECT 0.915 442.320 1095.530 443.720 ;
        RECT 0.915 433.520 1095.930 442.320 ;
        RECT 0.915 432.120 1095.530 433.520 ;
        RECT 0.915 423.320 1095.930 432.120 ;
        RECT 0.915 421.920 1095.530 423.320 ;
        RECT 0.915 413.120 1095.930 421.920 ;
        RECT 0.915 411.720 1095.530 413.120 ;
        RECT 0.915 402.920 1095.930 411.720 ;
        RECT 0.915 401.520 1095.530 402.920 ;
        RECT 0.915 392.720 1095.930 401.520 ;
        RECT 0.915 391.320 1095.530 392.720 ;
        RECT 0.915 382.520 1095.930 391.320 ;
        RECT 0.915 381.120 1095.530 382.520 ;
        RECT 0.915 372.320 1095.930 381.120 ;
        RECT 0.915 370.920 1095.530 372.320 ;
        RECT 0.915 362.120 1095.930 370.920 ;
        RECT 0.915 360.720 1095.530 362.120 ;
        RECT 0.915 351.920 1095.930 360.720 ;
        RECT 0.915 350.520 1095.530 351.920 ;
        RECT 0.915 341.720 1095.930 350.520 ;
        RECT 0.915 340.320 1095.530 341.720 ;
        RECT 0.915 331.520 1095.930 340.320 ;
        RECT 0.915 330.120 1095.530 331.520 ;
        RECT 0.915 321.320 1095.930 330.120 ;
        RECT 0.915 319.920 1095.530 321.320 ;
        RECT 0.915 311.120 1095.930 319.920 ;
        RECT 0.915 309.720 1095.530 311.120 ;
        RECT 0.915 300.920 1095.930 309.720 ;
        RECT 0.915 299.520 1095.530 300.920 ;
        RECT 0.915 290.720 1095.930 299.520 ;
        RECT 0.915 289.320 1095.530 290.720 ;
        RECT 0.915 280.520 1095.930 289.320 ;
        RECT 0.915 279.120 1095.530 280.520 ;
        RECT 0.915 270.320 1095.930 279.120 ;
        RECT 0.915 268.920 1095.530 270.320 ;
        RECT 0.915 260.120 1095.930 268.920 ;
        RECT 0.915 258.720 1095.530 260.120 ;
        RECT 0.915 249.920 1095.930 258.720 ;
        RECT 0.915 248.520 1095.530 249.920 ;
        RECT 0.915 239.720 1095.930 248.520 ;
        RECT 0.915 238.320 1095.530 239.720 ;
        RECT 0.915 229.520 1095.930 238.320 ;
        RECT 0.915 228.120 1095.530 229.520 ;
        RECT 0.915 219.320 1095.930 228.120 ;
        RECT 0.915 217.920 1095.530 219.320 ;
        RECT 0.915 209.120 1095.930 217.920 ;
        RECT 0.915 207.720 1095.530 209.120 ;
        RECT 0.915 198.920 1095.930 207.720 ;
        RECT 0.915 197.520 1095.530 198.920 ;
        RECT 0.915 188.720 1095.930 197.520 ;
        RECT 0.915 187.320 1095.530 188.720 ;
        RECT 0.915 178.520 1095.930 187.320 ;
        RECT 0.915 177.120 1095.530 178.520 ;
        RECT 0.915 168.320 1095.930 177.120 ;
        RECT 0.915 166.920 1095.530 168.320 ;
        RECT 0.915 158.120 1095.930 166.920 ;
        RECT 0.915 156.720 1095.530 158.120 ;
        RECT 0.915 147.920 1095.930 156.720 ;
        RECT 0.915 146.520 1095.530 147.920 ;
        RECT 0.915 137.720 1095.930 146.520 ;
        RECT 0.915 136.320 1095.530 137.720 ;
        RECT 0.915 127.520 1095.930 136.320 ;
        RECT 0.915 126.120 1095.530 127.520 ;
        RECT 0.915 117.320 1095.930 126.120 ;
        RECT 0.915 115.920 1095.530 117.320 ;
        RECT 0.915 107.120 1095.930 115.920 ;
        RECT 0.915 105.720 1095.530 107.120 ;
        RECT 0.915 96.920 1095.930 105.720 ;
        RECT 0.915 95.520 1095.530 96.920 ;
        RECT 0.915 86.720 1095.930 95.520 ;
        RECT 0.915 85.320 1095.530 86.720 ;
        RECT 0.915 76.520 1095.930 85.320 ;
        RECT 0.915 75.120 1095.530 76.520 ;
        RECT 0.915 66.320 1095.930 75.120 ;
        RECT 0.915 64.920 1095.530 66.320 ;
        RECT 0.915 56.120 1095.930 64.920 ;
        RECT 0.915 54.720 1095.530 56.120 ;
        RECT 0.915 45.920 1095.930 54.720 ;
        RECT 0.915 44.520 1095.530 45.920 ;
        RECT 0.915 35.720 1095.930 44.520 ;
        RECT 0.915 34.320 1095.530 35.720 ;
        RECT 0.915 25.520 1095.930 34.320 ;
        RECT 0.915 24.120 1095.530 25.520 ;
        RECT 0.915 15.320 1095.930 24.120 ;
        RECT 0.915 13.920 1095.530 15.320 ;
        RECT 0.915 5.800 1095.930 13.920 ;
        RECT 0.915 4.935 1095.530 5.800 ;
      LAYER met4 ;
        RECT 66.465 10.640 97.370 1088.240 ;
        RECT 99.770 10.640 1087.995 1088.240 ;
  END
END hs32_core1
END LIBRARY

