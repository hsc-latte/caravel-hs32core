VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 289.410 89.660 289.730 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 289.410 89.520 2899.310 89.660 ;
        RECT 289.410 89.460 289.730 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 289.440 89.460 289.700 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 289.430 1604.955 289.710 1605.325 ;
        RECT 289.500 89.750 289.640 1604.955 ;
        RECT 289.440 89.430 289.700 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 289.430 1605.000 289.710 1605.280 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 289.405 1605.290 289.735 1605.305 ;
        RECT 300.000 1605.290 304.000 1605.400 ;
        RECT 289.405 1604.990 304.000 1605.290 ;
        RECT 289.405 1604.975 289.735 1604.990 ;
        RECT 300.000 1604.800 304.000 1604.990 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 288.030 2698.480 288.350 2698.540 ;
        RECT 2902.670 2698.480 2902.990 2698.540 ;
        RECT 288.030 2698.340 2902.990 2698.480 ;
        RECT 288.030 2698.280 288.350 2698.340 ;
        RECT 2902.670 2698.280 2902.990 2698.340 ;
      LAYER via ;
        RECT 288.060 2698.280 288.320 2698.540 ;
        RECT 2902.700 2698.280 2902.960 2698.540 ;
      LAYER met2 ;
        RECT 288.060 2698.250 288.320 2698.570 ;
        RECT 2902.700 2698.250 2902.960 2698.570 ;
        RECT 288.120 1894.325 288.260 2698.250 ;
        RECT 2902.760 2434.245 2902.900 2698.250 ;
        RECT 2902.690 2433.875 2902.970 2434.245 ;
        RECT 288.050 1893.955 288.330 1894.325 ;
      LAYER via2 ;
        RECT 2902.690 2433.920 2902.970 2434.200 ;
        RECT 288.050 1894.000 288.330 1894.280 ;
      LAYER met3 ;
        RECT 2902.665 2434.210 2902.995 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2902.665 2433.910 2924.800 2434.210 ;
        RECT 2902.665 2433.895 2902.995 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 288.025 1894.290 288.355 1894.305 ;
        RECT 300.000 1894.290 304.000 1894.400 ;
        RECT 288.025 1893.990 304.000 1894.290 ;
        RECT 288.025 1893.975 288.355 1893.990 ;
        RECT 300.000 1893.800 304.000 1893.990 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 297.690 2698.820 298.010 2698.880 ;
        RECT 2904.510 2698.820 2904.830 2698.880 ;
        RECT 297.690 2698.680 2904.830 2698.820 ;
        RECT 297.690 2698.620 298.010 2698.680 ;
        RECT 2904.510 2698.620 2904.830 2698.680 ;
      LAYER via ;
        RECT 297.720 2698.620 297.980 2698.880 ;
        RECT 2904.540 2698.620 2904.800 2698.880 ;
      LAYER met2 ;
        RECT 297.720 2698.590 297.980 2698.910 ;
        RECT 2904.540 2698.590 2904.800 2698.910 ;
        RECT 297.780 1923.565 297.920 2698.590 ;
        RECT 2904.600 2669.525 2904.740 2698.590 ;
        RECT 2904.530 2669.155 2904.810 2669.525 ;
        RECT 297.710 1923.195 297.990 1923.565 ;
      LAYER via2 ;
        RECT 2904.530 2669.200 2904.810 2669.480 ;
        RECT 297.710 1923.240 297.990 1923.520 ;
      LAYER met3 ;
        RECT 2904.505 2669.490 2904.835 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2904.505 2669.190 2924.800 2669.490 ;
        RECT 2904.505 2669.175 2904.835 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 297.685 1923.530 298.015 1923.545 ;
        RECT 300.000 1923.530 304.000 1923.640 ;
        RECT 297.685 1923.230 304.000 1923.530 ;
        RECT 297.685 1923.215 298.015 1923.230 ;
        RECT 300.000 1923.040 304.000 1923.230 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 298.150 2701.880 298.470 2701.940 ;
        RECT 2903.590 2701.880 2903.910 2701.940 ;
        RECT 298.150 2701.740 2903.910 2701.880 ;
        RECT 298.150 2701.680 298.470 2701.740 ;
        RECT 2903.590 2701.680 2903.910 2701.740 ;
      LAYER via ;
        RECT 298.180 2701.680 298.440 2701.940 ;
        RECT 2903.620 2701.680 2903.880 2701.940 ;
      LAYER met2 ;
        RECT 2903.610 2903.755 2903.890 2904.125 ;
        RECT 2903.680 2701.970 2903.820 2903.755 ;
        RECT 298.180 2701.650 298.440 2701.970 ;
        RECT 2903.620 2701.650 2903.880 2701.970 ;
        RECT 298.240 1952.125 298.380 2701.650 ;
        RECT 298.170 1951.755 298.450 1952.125 ;
      LAYER via2 ;
        RECT 2903.610 2903.800 2903.890 2904.080 ;
        RECT 298.170 1951.800 298.450 1952.080 ;
      LAYER met3 ;
        RECT 2903.585 2904.090 2903.915 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2903.585 2903.790 2924.800 2904.090 ;
        RECT 2903.585 2903.775 2903.915 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 298.145 1952.090 298.475 1952.105 ;
        RECT 300.000 1952.090 304.000 1952.200 ;
        RECT 298.145 1951.790 304.000 1952.090 ;
        RECT 298.145 1951.775 298.475 1951.790 ;
        RECT 300.000 1951.600 304.000 1951.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 298.610 2702.220 298.930 2702.280 ;
        RECT 2901.750 2702.220 2902.070 2702.280 ;
        RECT 298.610 2702.080 2902.070 2702.220 ;
        RECT 298.610 2702.020 298.930 2702.080 ;
        RECT 2901.750 2702.020 2902.070 2702.080 ;
      LAYER via ;
        RECT 298.640 2702.020 298.900 2702.280 ;
        RECT 2901.780 2702.020 2902.040 2702.280 ;
      LAYER met2 ;
        RECT 2901.770 3138.355 2902.050 3138.725 ;
        RECT 2901.840 2702.310 2901.980 3138.355 ;
        RECT 298.640 2701.990 298.900 2702.310 ;
        RECT 2901.780 2701.990 2902.040 2702.310 ;
        RECT 298.700 1981.365 298.840 2701.990 ;
        RECT 298.630 1980.995 298.910 1981.365 ;
      LAYER via2 ;
        RECT 2901.770 3138.400 2902.050 3138.680 ;
        RECT 298.630 1981.040 298.910 1981.320 ;
      LAYER met3 ;
        RECT 2901.745 3138.690 2902.075 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2901.745 3138.390 2924.800 3138.690 ;
        RECT 2901.745 3138.375 2902.075 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 298.605 1981.330 298.935 1981.345 ;
        RECT 300.000 1981.330 304.000 1981.440 ;
        RECT 298.605 1981.030 304.000 1981.330 ;
        RECT 298.605 1981.015 298.935 1981.030 ;
        RECT 300.000 1980.840 304.000 1981.030 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.470 3369.640 869.790 3369.700 ;
        RECT 893.850 3369.640 894.170 3369.700 ;
        RECT 869.470 3369.500 894.170 3369.640 ;
        RECT 869.470 3369.440 869.790 3369.500 ;
        RECT 893.850 3369.440 894.170 3369.500 ;
        RECT 1835.470 3369.640 1835.790 3369.700 ;
        RECT 1859.850 3369.640 1860.170 3369.700 ;
        RECT 1835.470 3369.500 1860.170 3369.640 ;
        RECT 1835.470 3369.440 1835.790 3369.500 ;
        RECT 1859.850 3369.440 1860.170 3369.500 ;
        RECT 2801.470 3369.640 2801.790 3369.700 ;
        RECT 2825.850 3369.640 2826.170 3369.700 ;
        RECT 2801.470 3369.500 2826.170 3369.640 ;
        RECT 2801.470 3369.440 2801.790 3369.500 ;
        RECT 2825.850 3369.440 2826.170 3369.500 ;
        RECT 772.870 3368.960 773.190 3369.020 ;
        RECT 811.050 3368.960 811.370 3369.020 ;
        RECT 772.870 3368.820 811.370 3368.960 ;
        RECT 772.870 3368.760 773.190 3368.820 ;
        RECT 811.050 3368.760 811.370 3368.820 ;
        RECT 1449.070 3368.960 1449.390 3369.020 ;
        RECT 1463.330 3368.960 1463.650 3369.020 ;
        RECT 1449.070 3368.820 1463.650 3368.960 ;
        RECT 1449.070 3368.760 1449.390 3368.820 ;
        RECT 1463.330 3368.760 1463.650 3368.820 ;
        RECT 1738.870 3368.960 1739.190 3369.020 ;
        RECT 1777.050 3368.960 1777.370 3369.020 ;
        RECT 1738.870 3368.820 1777.370 3368.960 ;
        RECT 1738.870 3368.760 1739.190 3368.820 ;
        RECT 1777.050 3368.760 1777.370 3368.820 ;
        RECT 2704.870 3368.960 2705.190 3369.020 ;
        RECT 2743.050 3368.960 2743.370 3369.020 ;
        RECT 2704.870 3368.820 2743.370 3368.960 ;
        RECT 2704.870 3368.760 2705.190 3368.820 ;
        RECT 2743.050 3368.760 2743.370 3368.820 ;
      LAYER via ;
        RECT 869.500 3369.440 869.760 3369.700 ;
        RECT 893.880 3369.440 894.140 3369.700 ;
        RECT 1835.500 3369.440 1835.760 3369.700 ;
        RECT 1859.880 3369.440 1860.140 3369.700 ;
        RECT 2801.500 3369.440 2801.760 3369.700 ;
        RECT 2825.880 3369.440 2826.140 3369.700 ;
        RECT 772.900 3368.760 773.160 3369.020 ;
        RECT 811.080 3368.760 811.340 3369.020 ;
        RECT 1449.100 3368.760 1449.360 3369.020 ;
        RECT 1463.360 3368.760 1463.620 3369.020 ;
        RECT 1738.900 3368.760 1739.160 3369.020 ;
        RECT 1777.080 3368.760 1777.340 3369.020 ;
        RECT 2704.900 3368.760 2705.160 3369.020 ;
        RECT 2743.080 3368.760 2743.340 3369.020 ;
      LAYER met2 ;
        RECT 941.710 3370.235 941.990 3370.605 ;
        RECT 1897.590 3370.235 1897.870 3370.605 ;
        RECT 834.990 3369.555 835.270 3369.925 ;
        RECT 869.490 3369.555 869.770 3369.925 ;
        RECT 772.890 3368.875 773.170 3369.245 ;
        RECT 772.900 3368.730 773.160 3368.875 ;
        RECT 811.080 3368.730 811.340 3369.050 ;
        RECT 811.140 3367.885 811.280 3368.730 ;
        RECT 811.070 3367.515 811.350 3367.885 ;
        RECT 834.530 3367.770 834.810 3367.885 ;
        RECT 835.060 3367.770 835.200 3369.555 ;
        RECT 869.500 3369.410 869.760 3369.555 ;
        RECT 893.880 3369.410 894.140 3369.730 ;
        RECT 893.940 3369.245 894.080 3369.410 ;
        RECT 941.780 3369.245 941.920 3370.235 ;
        RECT 1800.530 3369.810 1800.810 3369.925 ;
        RECT 1801.450 3369.810 1801.730 3369.925 ;
        RECT 1800.530 3369.670 1801.730 3369.810 ;
        RECT 1800.530 3369.555 1800.810 3369.670 ;
        RECT 1801.450 3369.555 1801.730 3369.670 ;
        RECT 1835.490 3369.555 1835.770 3369.925 ;
        RECT 1835.500 3369.410 1835.760 3369.555 ;
        RECT 1859.880 3369.410 1860.140 3369.730 ;
        RECT 1859.940 3369.245 1860.080 3369.410 ;
        RECT 1897.660 3369.245 1897.800 3370.235 ;
        RECT 2766.990 3369.555 2767.270 3369.925 ;
        RECT 2801.490 3369.555 2801.770 3369.925 ;
        RECT 893.870 3368.875 894.150 3369.245 ;
        RECT 941.710 3368.875 941.990 3369.245 ;
        RECT 1449.090 3368.875 1449.370 3369.245 ;
        RECT 1449.100 3368.730 1449.360 3368.875 ;
        RECT 1463.360 3368.730 1463.620 3369.050 ;
        RECT 1738.890 3368.875 1739.170 3369.245 ;
        RECT 1738.900 3368.730 1739.160 3368.875 ;
        RECT 1777.080 3368.730 1777.340 3369.050 ;
        RECT 1859.870 3368.875 1860.150 3369.245 ;
        RECT 1897.590 3368.875 1897.870 3369.245 ;
        RECT 2704.890 3368.875 2705.170 3369.245 ;
        RECT 2704.900 3368.730 2705.160 3368.875 ;
        RECT 2743.080 3368.730 2743.340 3369.050 ;
        RECT 1463.420 3367.885 1463.560 3368.730 ;
        RECT 1777.140 3367.885 1777.280 3368.730 ;
        RECT 2743.140 3367.885 2743.280 3368.730 ;
        RECT 834.530 3367.630 835.200 3367.770 ;
        RECT 834.530 3367.515 834.810 3367.630 ;
        RECT 1463.350 3367.515 1463.630 3367.885 ;
        RECT 1777.070 3367.515 1777.350 3367.885 ;
        RECT 2743.070 3367.515 2743.350 3367.885 ;
        RECT 2766.530 3367.770 2766.810 3367.885 ;
        RECT 2767.060 3367.770 2767.200 3369.555 ;
        RECT 2801.500 3369.410 2801.760 3369.555 ;
        RECT 2825.880 3369.410 2826.140 3369.730 ;
        RECT 2825.940 3369.245 2826.080 3369.410 ;
        RECT 2825.870 3368.875 2826.150 3369.245 ;
        RECT 2863.590 3369.130 2863.870 3369.245 ;
        RECT 2863.200 3368.990 2863.870 3369.130 ;
        RECT 2863.200 3368.565 2863.340 3368.990 ;
        RECT 2863.590 3368.875 2863.870 3368.990 ;
        RECT 2863.130 3368.195 2863.410 3368.565 ;
        RECT 2766.530 3367.630 2767.200 3367.770 ;
        RECT 2766.530 3367.515 2766.810 3367.630 ;
      LAYER via2 ;
        RECT 941.710 3370.280 941.990 3370.560 ;
        RECT 1897.590 3370.280 1897.870 3370.560 ;
        RECT 834.990 3369.600 835.270 3369.880 ;
        RECT 869.490 3369.600 869.770 3369.880 ;
        RECT 772.890 3368.920 773.170 3369.200 ;
        RECT 811.070 3367.560 811.350 3367.840 ;
        RECT 834.530 3367.560 834.810 3367.840 ;
        RECT 1800.530 3369.600 1800.810 3369.880 ;
        RECT 1801.450 3369.600 1801.730 3369.880 ;
        RECT 1835.490 3369.600 1835.770 3369.880 ;
        RECT 2766.990 3369.600 2767.270 3369.880 ;
        RECT 2801.490 3369.600 2801.770 3369.880 ;
        RECT 893.870 3368.920 894.150 3369.200 ;
        RECT 941.710 3368.920 941.990 3369.200 ;
        RECT 1449.090 3368.920 1449.370 3369.200 ;
        RECT 1738.890 3368.920 1739.170 3369.200 ;
        RECT 1859.870 3368.920 1860.150 3369.200 ;
        RECT 1897.590 3368.920 1897.870 3369.200 ;
        RECT 2704.890 3368.920 2705.170 3369.200 ;
        RECT 1463.350 3367.560 1463.630 3367.840 ;
        RECT 1777.070 3367.560 1777.350 3367.840 ;
        RECT 2743.070 3367.560 2743.350 3367.840 ;
        RECT 2766.530 3367.560 2766.810 3367.840 ;
        RECT 2825.870 3368.920 2826.150 3369.200 ;
        RECT 2863.590 3368.920 2863.870 3369.200 ;
        RECT 2863.130 3368.240 2863.410 3368.520 ;
      LAYER met3 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2916.710 3372.990 2924.800 3373.290 ;
        RECT 917.510 3370.570 917.890 3370.580 ;
        RECT 941.685 3370.570 942.015 3370.585 ;
        RECT 917.510 3370.270 942.015 3370.570 ;
        RECT 917.510 3370.260 917.890 3370.270 ;
        RECT 941.685 3370.255 942.015 3370.270 ;
        RECT 1883.510 3370.570 1883.890 3370.580 ;
        RECT 1897.565 3370.570 1897.895 3370.585 ;
        RECT 1883.510 3370.270 1897.895 3370.570 ;
        RECT 1883.510 3370.260 1883.890 3370.270 ;
        RECT 1897.565 3370.255 1897.895 3370.270 ;
        RECT 834.965 3369.890 835.295 3369.905 ;
        RECT 869.465 3369.890 869.795 3369.905 ;
        RECT 834.965 3369.590 869.795 3369.890 ;
        RECT 834.965 3369.575 835.295 3369.590 ;
        RECT 869.465 3369.575 869.795 3369.590 ;
        RECT 1786.910 3369.890 1787.290 3369.900 ;
        RECT 1800.505 3369.890 1800.835 3369.905 ;
        RECT 1786.910 3369.590 1800.835 3369.890 ;
        RECT 1786.910 3369.580 1787.290 3369.590 ;
        RECT 1800.505 3369.575 1800.835 3369.590 ;
        RECT 1801.425 3369.890 1801.755 3369.905 ;
        RECT 1835.465 3369.890 1835.795 3369.905 ;
        RECT 1801.425 3369.590 1835.795 3369.890 ;
        RECT 1801.425 3369.575 1801.755 3369.590 ;
        RECT 1835.465 3369.575 1835.795 3369.590 ;
        RECT 2766.965 3369.890 2767.295 3369.905 ;
        RECT 2801.465 3369.890 2801.795 3369.905 ;
        RECT 2766.965 3369.590 2801.795 3369.890 ;
        RECT 2766.965 3369.575 2767.295 3369.590 ;
        RECT 2801.465 3369.575 2801.795 3369.590 ;
        RECT 296.510 3369.210 296.890 3369.220 ;
        RECT 772.865 3369.210 773.195 3369.225 ;
        RECT 296.510 3368.910 324.450 3369.210 ;
        RECT 296.510 3368.900 296.890 3368.910 ;
        RECT 324.150 3368.530 324.450 3368.910 ;
        RECT 372.910 3368.910 421.050 3369.210 ;
        RECT 324.150 3368.230 372.290 3368.530 ;
        RECT 371.990 3367.850 372.290 3368.230 ;
        RECT 372.910 3367.850 373.210 3368.910 ;
        RECT 420.750 3368.530 421.050 3368.910 ;
        RECT 469.510 3368.910 517.650 3369.210 ;
        RECT 420.750 3368.230 468.890 3368.530 ;
        RECT 371.990 3367.550 373.210 3367.850 ;
        RECT 468.590 3367.850 468.890 3368.230 ;
        RECT 469.510 3367.850 469.810 3368.910 ;
        RECT 517.350 3368.530 517.650 3368.910 ;
        RECT 566.110 3368.910 614.250 3369.210 ;
        RECT 517.350 3368.230 565.490 3368.530 ;
        RECT 468.590 3367.550 469.810 3367.850 ;
        RECT 565.190 3367.850 565.490 3368.230 ;
        RECT 566.110 3367.850 566.410 3368.910 ;
        RECT 613.950 3368.530 614.250 3368.910 ;
        RECT 662.710 3368.910 710.850 3369.210 ;
        RECT 613.950 3368.230 662.090 3368.530 ;
        RECT 565.190 3367.550 566.410 3367.850 ;
        RECT 661.790 3367.850 662.090 3368.230 ;
        RECT 662.710 3367.850 663.010 3368.910 ;
        RECT 710.550 3368.530 710.850 3368.910 ;
        RECT 759.310 3368.910 773.195 3369.210 ;
        RECT 710.550 3368.230 758.690 3368.530 ;
        RECT 661.790 3367.550 663.010 3367.850 ;
        RECT 758.390 3367.850 758.690 3368.230 ;
        RECT 759.310 3367.850 759.610 3368.910 ;
        RECT 772.865 3368.895 773.195 3368.910 ;
        RECT 893.845 3369.210 894.175 3369.225 ;
        RECT 917.510 3369.210 917.890 3369.220 ;
        RECT 893.845 3368.910 917.890 3369.210 ;
        RECT 893.845 3368.895 894.175 3368.910 ;
        RECT 917.510 3368.900 917.890 3368.910 ;
        RECT 941.685 3369.210 942.015 3369.225 ;
        RECT 1449.065 3369.210 1449.395 3369.225 ;
        RECT 941.685 3368.910 1000.650 3369.210 ;
        RECT 941.685 3368.895 942.015 3368.910 ;
        RECT 1000.350 3368.530 1000.650 3368.910 ;
        RECT 1049.110 3368.910 1097.250 3369.210 ;
        RECT 1000.350 3368.230 1048.490 3368.530 ;
        RECT 758.390 3367.550 759.610 3367.850 ;
        RECT 811.045 3367.850 811.375 3367.865 ;
        RECT 834.505 3367.850 834.835 3367.865 ;
        RECT 811.045 3367.550 834.835 3367.850 ;
        RECT 1048.190 3367.850 1048.490 3368.230 ;
        RECT 1049.110 3367.850 1049.410 3368.910 ;
        RECT 1096.950 3368.530 1097.250 3368.910 ;
        RECT 1145.710 3368.910 1193.850 3369.210 ;
        RECT 1096.950 3368.230 1145.090 3368.530 ;
        RECT 1048.190 3367.550 1049.410 3367.850 ;
        RECT 1144.790 3367.850 1145.090 3368.230 ;
        RECT 1145.710 3367.850 1146.010 3368.910 ;
        RECT 1193.550 3368.530 1193.850 3368.910 ;
        RECT 1242.310 3368.910 1290.450 3369.210 ;
        RECT 1193.550 3368.230 1241.690 3368.530 ;
        RECT 1144.790 3367.550 1146.010 3367.850 ;
        RECT 1241.390 3367.850 1241.690 3368.230 ;
        RECT 1242.310 3367.850 1242.610 3368.910 ;
        RECT 1290.150 3368.530 1290.450 3368.910 ;
        RECT 1338.910 3368.910 1387.050 3369.210 ;
        RECT 1290.150 3368.230 1338.290 3368.530 ;
        RECT 1241.390 3367.550 1242.610 3367.850 ;
        RECT 1337.990 3367.850 1338.290 3368.230 ;
        RECT 1338.910 3367.850 1339.210 3368.910 ;
        RECT 1386.750 3368.530 1387.050 3368.910 ;
        RECT 1435.510 3368.910 1449.395 3369.210 ;
        RECT 1386.750 3368.230 1434.890 3368.530 ;
        RECT 1337.990 3367.550 1339.210 3367.850 ;
        RECT 1434.590 3367.850 1434.890 3368.230 ;
        RECT 1435.510 3367.850 1435.810 3368.910 ;
        RECT 1449.065 3368.895 1449.395 3368.910 ;
        RECT 1497.110 3369.210 1497.490 3369.220 ;
        RECT 1738.865 3369.210 1739.195 3369.225 ;
        RECT 1497.110 3368.910 1580.250 3369.210 ;
        RECT 1497.110 3368.900 1497.490 3368.910 ;
        RECT 1579.950 3368.530 1580.250 3368.910 ;
        RECT 1628.710 3368.910 1676.850 3369.210 ;
        RECT 1579.950 3368.230 1628.090 3368.530 ;
        RECT 1434.590 3367.550 1435.810 3367.850 ;
        RECT 1463.325 3367.850 1463.655 3367.865 ;
        RECT 1497.110 3367.850 1497.490 3367.860 ;
        RECT 1463.325 3367.550 1497.490 3367.850 ;
        RECT 1627.790 3367.850 1628.090 3368.230 ;
        RECT 1628.710 3367.850 1629.010 3368.910 ;
        RECT 1676.550 3368.530 1676.850 3368.910 ;
        RECT 1725.310 3368.910 1739.195 3369.210 ;
        RECT 1676.550 3368.230 1724.690 3368.530 ;
        RECT 1627.790 3367.550 1629.010 3367.850 ;
        RECT 1724.390 3367.850 1724.690 3368.230 ;
        RECT 1725.310 3367.850 1725.610 3368.910 ;
        RECT 1738.865 3368.895 1739.195 3368.910 ;
        RECT 1859.845 3369.210 1860.175 3369.225 ;
        RECT 1883.510 3369.210 1883.890 3369.220 ;
        RECT 1859.845 3368.910 1883.890 3369.210 ;
        RECT 1859.845 3368.895 1860.175 3368.910 ;
        RECT 1883.510 3368.900 1883.890 3368.910 ;
        RECT 1897.565 3369.210 1897.895 3369.225 ;
        RECT 2704.865 3369.210 2705.195 3369.225 ;
        RECT 1897.565 3368.910 1966.650 3369.210 ;
        RECT 1897.565 3368.895 1897.895 3368.910 ;
        RECT 1966.350 3368.530 1966.650 3368.910 ;
        RECT 2015.110 3368.910 2063.250 3369.210 ;
        RECT 1966.350 3368.230 2014.490 3368.530 ;
        RECT 1724.390 3367.550 1725.610 3367.850 ;
        RECT 1777.045 3367.850 1777.375 3367.865 ;
        RECT 1786.910 3367.850 1787.290 3367.860 ;
        RECT 1777.045 3367.550 1787.290 3367.850 ;
        RECT 2014.190 3367.850 2014.490 3368.230 ;
        RECT 2015.110 3367.850 2015.410 3368.910 ;
        RECT 2062.950 3368.530 2063.250 3368.910 ;
        RECT 2159.550 3368.910 2207.690 3369.210 ;
        RECT 2062.950 3368.230 2111.090 3368.530 ;
        RECT 2014.190 3367.550 2015.410 3367.850 ;
        RECT 2110.790 3367.850 2111.090 3368.230 ;
        RECT 2159.550 3367.850 2159.850 3368.910 ;
        RECT 2110.790 3367.550 2159.850 3367.850 ;
        RECT 2207.390 3367.850 2207.690 3368.910 ;
        RECT 2208.310 3368.910 2256.450 3369.210 ;
        RECT 2208.310 3367.850 2208.610 3368.910 ;
        RECT 2256.150 3368.530 2256.450 3368.910 ;
        RECT 2304.910 3368.910 2353.050 3369.210 ;
        RECT 2256.150 3368.230 2304.290 3368.530 ;
        RECT 2207.390 3367.550 2208.610 3367.850 ;
        RECT 2303.990 3367.850 2304.290 3368.230 ;
        RECT 2304.910 3367.850 2305.210 3368.910 ;
        RECT 2352.750 3368.530 2353.050 3368.910 ;
        RECT 2401.510 3368.910 2449.650 3369.210 ;
        RECT 2352.750 3368.230 2400.890 3368.530 ;
        RECT 2303.990 3367.550 2305.210 3367.850 ;
        RECT 2400.590 3367.850 2400.890 3368.230 ;
        RECT 2401.510 3367.850 2401.810 3368.910 ;
        RECT 2449.350 3368.530 2449.650 3368.910 ;
        RECT 2498.110 3368.910 2546.250 3369.210 ;
        RECT 2449.350 3368.230 2497.490 3368.530 ;
        RECT 2400.590 3367.550 2401.810 3367.850 ;
        RECT 2497.190 3367.850 2497.490 3368.230 ;
        RECT 2498.110 3367.850 2498.410 3368.910 ;
        RECT 2545.950 3368.530 2546.250 3368.910 ;
        RECT 2594.710 3368.910 2642.850 3369.210 ;
        RECT 2545.950 3368.230 2594.090 3368.530 ;
        RECT 2497.190 3367.550 2498.410 3367.850 ;
        RECT 2593.790 3367.850 2594.090 3368.230 ;
        RECT 2594.710 3367.850 2595.010 3368.910 ;
        RECT 2642.550 3368.530 2642.850 3368.910 ;
        RECT 2691.310 3368.910 2705.195 3369.210 ;
        RECT 2642.550 3368.230 2690.690 3368.530 ;
        RECT 2593.790 3367.550 2595.010 3367.850 ;
        RECT 2690.390 3367.850 2690.690 3368.230 ;
        RECT 2691.310 3367.850 2691.610 3368.910 ;
        RECT 2704.865 3368.895 2705.195 3368.910 ;
        RECT 2825.845 3369.210 2826.175 3369.225 ;
        RECT 2863.565 3369.210 2863.895 3369.225 ;
        RECT 2825.845 3368.910 2849.850 3369.210 ;
        RECT 2825.845 3368.895 2826.175 3368.910 ;
        RECT 2849.550 3368.530 2849.850 3368.910 ;
        RECT 2863.565 3368.910 2884.810 3369.210 ;
        RECT 2863.565 3368.895 2863.895 3368.910 ;
        RECT 2863.105 3368.530 2863.435 3368.545 ;
        RECT 2849.550 3368.230 2863.435 3368.530 ;
        RECT 2884.510 3368.530 2884.810 3368.910 ;
        RECT 2916.710 3368.530 2917.010 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2884.510 3368.230 2917.010 3368.530 ;
        RECT 2863.105 3368.215 2863.435 3368.230 ;
        RECT 2690.390 3367.550 2691.610 3367.850 ;
        RECT 2743.045 3367.850 2743.375 3367.865 ;
        RECT 2766.505 3367.850 2766.835 3367.865 ;
        RECT 2743.045 3367.550 2766.835 3367.850 ;
        RECT 811.045 3367.535 811.375 3367.550 ;
        RECT 834.505 3367.535 834.835 3367.550 ;
        RECT 1463.325 3367.535 1463.655 3367.550 ;
        RECT 1497.110 3367.540 1497.490 3367.550 ;
        RECT 1777.045 3367.535 1777.375 3367.550 ;
        RECT 1786.910 3367.540 1787.290 3367.550 ;
        RECT 2743.045 3367.535 2743.375 3367.550 ;
        RECT 2766.505 3367.535 2766.835 3367.550 ;
        RECT 296.510 2010.570 296.890 2010.580 ;
        RECT 300.000 2010.570 304.000 2010.680 ;
        RECT 296.510 2010.270 304.000 2010.570 ;
        RECT 296.510 2010.260 296.890 2010.270 ;
        RECT 300.000 2010.080 304.000 2010.270 ;
      LAYER via3 ;
        RECT 917.540 3370.260 917.860 3370.580 ;
        RECT 1883.540 3370.260 1883.860 3370.580 ;
        RECT 1786.940 3369.580 1787.260 3369.900 ;
        RECT 296.540 3368.900 296.860 3369.220 ;
        RECT 917.540 3368.900 917.860 3369.220 ;
        RECT 1497.140 3368.900 1497.460 3369.220 ;
        RECT 1497.140 3367.540 1497.460 3367.860 ;
        RECT 1883.540 3368.900 1883.860 3369.220 ;
        RECT 1786.940 3367.540 1787.260 3367.860 ;
        RECT 296.540 2010.260 296.860 2010.580 ;
      LAYER met4 ;
        RECT 917.535 3370.255 917.865 3370.585 ;
        RECT 1883.535 3370.255 1883.865 3370.585 ;
        RECT 917.550 3369.225 917.850 3370.255 ;
        RECT 1786.935 3369.575 1787.265 3369.905 ;
        RECT 296.535 3368.895 296.865 3369.225 ;
        RECT 917.535 3368.895 917.865 3369.225 ;
        RECT 1497.135 3368.895 1497.465 3369.225 ;
        RECT 296.550 2010.585 296.850 3368.895 ;
        RECT 1497.150 3367.865 1497.450 3368.895 ;
        RECT 1786.950 3367.865 1787.250 3369.575 ;
        RECT 1883.550 3369.225 1883.850 3370.255 ;
        RECT 1883.535 3368.895 1883.865 3369.225 ;
        RECT 1497.135 3367.535 1497.465 3367.865 ;
        RECT 1786.935 3367.535 1787.265 3367.865 ;
        RECT 296.535 2010.255 296.865 2010.585 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2795.030 3422.680 2795.350 3422.740 ;
        RECT 2798.250 3422.680 2798.570 3422.740 ;
        RECT 2795.030 3422.540 2798.570 3422.680 ;
        RECT 2795.030 3422.480 2795.350 3422.540 ;
        RECT 2798.250 3422.480 2798.570 3422.540 ;
        RECT 2795.030 3374.400 2795.350 3374.460 ;
        RECT 2796.870 3374.400 2797.190 3374.460 ;
        RECT 2795.030 3374.260 2797.190 3374.400 ;
        RECT 2795.030 3374.200 2795.350 3374.260 ;
        RECT 2796.870 3374.200 2797.190 3374.260 ;
        RECT 2795.490 3308.780 2795.810 3308.840 ;
        RECT 2796.870 3308.780 2797.190 3308.840 ;
        RECT 2795.490 3308.640 2797.190 3308.780 ;
        RECT 2795.490 3308.580 2795.810 3308.640 ;
        RECT 2796.870 3308.580 2797.190 3308.640 ;
        RECT 2795.490 3284.640 2795.810 3284.700 ;
        RECT 2795.950 3284.640 2796.270 3284.700 ;
        RECT 2795.490 3284.500 2796.270 3284.640 ;
        RECT 2795.490 3284.440 2795.810 3284.500 ;
        RECT 2795.950 3284.440 2796.270 3284.500 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.030 3042.900 2795.350 3042.960 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.030 3042.760 2795.810 3042.900 ;
        RECT 2795.030 3042.700 2795.350 3042.760 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.030 3008.560 2795.350 3008.620 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.030 3008.420 2796.730 3008.560 ;
        RECT 2795.030 3008.360 2795.350 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2795.490 2994.620 2795.810 2994.680 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2795.490 2994.480 2796.730 2994.620 ;
        RECT 2795.490 2994.420 2795.810 2994.480 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2795.490 2946.680 2795.810 2946.740 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2795.490 2946.540 2797.190 2946.680 ;
        RECT 2795.490 2946.480 2795.810 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 2796.870 2912.340 2797.190 2912.400 ;
        RECT 2796.500 2912.200 2797.190 2912.340 ;
        RECT 2796.500 2911.720 2796.640 2912.200 ;
        RECT 2796.870 2912.140 2797.190 2912.200 ;
        RECT 2796.410 2911.460 2796.730 2911.720 ;
        RECT 2795.030 2801.500 2795.350 2801.560 ;
        RECT 2795.490 2801.500 2795.810 2801.560 ;
        RECT 2795.030 2801.360 2795.810 2801.500 ;
        RECT 2795.030 2801.300 2795.350 2801.360 ;
        RECT 2795.490 2801.300 2795.810 2801.360 ;
      LAYER via ;
        RECT 2795.060 3422.480 2795.320 3422.740 ;
        RECT 2798.280 3422.480 2798.540 3422.740 ;
        RECT 2795.060 3374.200 2795.320 3374.460 ;
        RECT 2796.900 3374.200 2797.160 3374.460 ;
        RECT 2795.520 3308.580 2795.780 3308.840 ;
        RECT 2796.900 3308.580 2797.160 3308.840 ;
        RECT 2795.520 3284.440 2795.780 3284.700 ;
        RECT 2795.980 3284.440 2796.240 3284.700 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.060 3042.700 2795.320 3042.960 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2795.060 3008.360 2795.320 3008.620 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2795.520 2994.420 2795.780 2994.680 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2795.520 2946.480 2795.780 2946.740 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 2796.900 2912.140 2797.160 2912.400 ;
        RECT 2796.440 2911.460 2796.700 2911.720 ;
        RECT 2795.060 2801.300 2795.320 2801.560 ;
        RECT 2795.520 2801.300 2795.780 2801.560 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3422.770 2798.480 3517.600 ;
        RECT 2795.060 3422.450 2795.320 3422.770 ;
        RECT 2798.280 3422.450 2798.540 3422.770 ;
        RECT 2795.120 3422.285 2795.260 3422.450 ;
        RECT 2795.050 3421.915 2795.330 3422.285 ;
        RECT 2795.050 3421.235 2795.330 3421.605 ;
        RECT 2795.120 3374.490 2795.260 3421.235 ;
        RECT 2795.060 3374.170 2795.320 3374.490 ;
        RECT 2796.900 3374.170 2797.160 3374.490 ;
        RECT 2796.960 3308.870 2797.100 3374.170 ;
        RECT 2795.520 3308.550 2795.780 3308.870 ;
        RECT 2796.900 3308.550 2797.160 3308.870 ;
        RECT 2795.580 3284.730 2795.720 3308.550 ;
        RECT 2795.520 3284.410 2795.780 3284.730 ;
        RECT 2795.980 3284.410 2796.240 3284.730 ;
        RECT 2796.040 3236.450 2796.180 3284.410 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.060 3042.670 2795.320 3042.990 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2795.120 3008.650 2795.260 3042.670 ;
        RECT 2795.060 3008.330 2795.320 3008.650 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2795.520 2994.390 2795.780 2994.710 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2795.580 2946.770 2795.720 2994.390 ;
        RECT 2795.520 2946.450 2795.780 2946.770 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2912.430 2797.100 2946.450 ;
        RECT 2796.900 2912.110 2797.160 2912.430 ;
        RECT 2796.440 2911.430 2796.700 2911.750 ;
        RECT 2796.500 2863.210 2796.640 2911.430 ;
        RECT 2795.580 2863.070 2796.640 2863.210 ;
        RECT 2795.580 2801.590 2795.720 2863.070 ;
        RECT 2795.060 2801.270 2795.320 2801.590 ;
        RECT 2795.520 2801.270 2795.780 2801.590 ;
        RECT 2795.120 2766.650 2795.260 2801.270 ;
        RECT 2795.120 2766.510 2795.720 2766.650 ;
        RECT 2795.580 2719.050 2795.720 2766.510 ;
        RECT 2795.580 2718.910 2796.180 2719.050 ;
        RECT 2796.040 2702.165 2796.180 2718.910 ;
        RECT 2795.970 2701.795 2796.250 2702.165 ;
      LAYER via2 ;
        RECT 2795.050 3421.960 2795.330 3422.240 ;
        RECT 2795.050 3421.280 2795.330 3421.560 ;
        RECT 2795.970 2701.840 2796.250 2702.120 ;
      LAYER met3 ;
        RECT 2795.025 3421.935 2795.355 3422.265 ;
        RECT 2795.040 3421.585 2795.340 3421.935 ;
        RECT 2795.025 3421.255 2795.355 3421.585 ;
        RECT 297.430 2702.130 297.810 2702.140 ;
        RECT 2795.945 2702.130 2796.275 2702.145 ;
        RECT 297.430 2701.830 2796.275 2702.130 ;
        RECT 297.430 2701.820 297.810 2701.830 ;
        RECT 2795.945 2701.815 2796.275 2701.830 ;
        RECT 297.430 2039.130 297.810 2039.140 ;
        RECT 300.000 2039.130 304.000 2039.240 ;
        RECT 297.430 2038.830 304.000 2039.130 ;
        RECT 297.430 2038.820 297.810 2038.830 ;
        RECT 300.000 2038.640 304.000 2038.830 ;
      LAYER via3 ;
        RECT 297.460 2701.820 297.780 2702.140 ;
        RECT 297.460 2038.820 297.780 2039.140 ;
      LAYER met4 ;
        RECT 297.455 2701.815 297.785 2702.145 ;
        RECT 297.470 2039.145 297.770 2701.815 ;
        RECT 297.455 2038.815 297.785 2039.145 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2470.270 3464.160 2470.590 3464.220 ;
        RECT 2474.410 3464.160 2474.730 3464.220 ;
        RECT 2470.270 3464.020 2474.730 3464.160 ;
        RECT 2470.270 3463.960 2470.590 3464.020 ;
        RECT 2474.410 3463.960 2474.730 3464.020 ;
        RECT 2470.270 3367.600 2470.590 3367.660 ;
        RECT 2471.190 3367.600 2471.510 3367.660 ;
        RECT 2470.270 3367.460 2471.510 3367.600 ;
        RECT 2470.270 3367.400 2470.590 3367.460 ;
        RECT 2471.190 3367.400 2471.510 3367.460 ;
        RECT 2470.270 3346.520 2470.590 3346.580 ;
        RECT 2471.190 3346.520 2471.510 3346.580 ;
        RECT 2470.270 3346.380 2471.510 3346.520 ;
        RECT 2470.270 3346.320 2470.590 3346.380 ;
        RECT 2471.190 3346.320 2471.510 3346.380 ;
        RECT 2469.810 3332.580 2470.130 3332.640 ;
        RECT 2471.190 3332.580 2471.510 3332.640 ;
        RECT 2469.810 3332.440 2471.510 3332.580 ;
        RECT 2469.810 3332.380 2470.130 3332.440 ;
        RECT 2471.190 3332.380 2471.510 3332.440 ;
        RECT 2469.810 3284.640 2470.130 3284.700 ;
        RECT 2470.730 3284.640 2471.050 3284.700 ;
        RECT 2469.810 3284.500 2471.050 3284.640 ;
        RECT 2469.810 3284.440 2470.130 3284.500 ;
        RECT 2470.730 3284.440 2471.050 3284.500 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 2469.350 2946.340 2469.670 2946.400 ;
        RECT 2470.730 2946.340 2471.050 2946.400 ;
        RECT 2469.350 2946.200 2471.050 2946.340 ;
        RECT 2469.350 2946.140 2469.670 2946.200 ;
        RECT 2470.730 2946.140 2471.050 2946.200 ;
        RECT 2469.350 2898.400 2469.670 2898.460 ;
        RECT 2470.270 2898.400 2470.590 2898.460 ;
        RECT 2469.350 2898.260 2470.590 2898.400 ;
        RECT 2469.350 2898.200 2469.670 2898.260 ;
        RECT 2470.270 2898.200 2470.590 2898.260 ;
        RECT 2470.730 2849.440 2471.050 2849.500 ;
        RECT 2471.650 2849.440 2471.970 2849.500 ;
        RECT 2470.730 2849.300 2471.970 2849.440 ;
        RECT 2470.730 2849.240 2471.050 2849.300 ;
        RECT 2471.650 2849.240 2471.970 2849.300 ;
        RECT 2471.650 2815.920 2471.970 2816.180 ;
        RECT 2471.740 2815.500 2471.880 2815.920 ;
        RECT 2471.650 2815.240 2471.970 2815.500 ;
        RECT 299.070 2702.560 299.390 2702.620 ;
        RECT 2458.770 2702.560 2459.090 2702.620 ;
        RECT 299.070 2702.420 2459.090 2702.560 ;
        RECT 299.070 2702.360 299.390 2702.420 ;
        RECT 2458.770 2702.360 2459.090 2702.420 ;
      LAYER via ;
        RECT 2470.300 3463.960 2470.560 3464.220 ;
        RECT 2474.440 3463.960 2474.700 3464.220 ;
        RECT 2470.300 3367.400 2470.560 3367.660 ;
        RECT 2471.220 3367.400 2471.480 3367.660 ;
        RECT 2470.300 3346.320 2470.560 3346.580 ;
        RECT 2471.220 3346.320 2471.480 3346.580 ;
        RECT 2469.840 3332.380 2470.100 3332.640 ;
        RECT 2471.220 3332.380 2471.480 3332.640 ;
        RECT 2469.840 3284.440 2470.100 3284.700 ;
        RECT 2470.760 3284.440 2471.020 3284.700 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 2469.380 2946.140 2469.640 2946.400 ;
        RECT 2470.760 2946.140 2471.020 2946.400 ;
        RECT 2469.380 2898.200 2469.640 2898.460 ;
        RECT 2470.300 2898.200 2470.560 2898.460 ;
        RECT 2470.760 2849.240 2471.020 2849.500 ;
        RECT 2471.680 2849.240 2471.940 2849.500 ;
        RECT 2471.680 2815.920 2471.940 2816.180 ;
        RECT 2471.680 2815.240 2471.940 2815.500 ;
        RECT 299.100 2702.360 299.360 2702.620 ;
        RECT 2458.800 2702.360 2459.060 2702.620 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3464.250 2474.640 3517.230 ;
        RECT 2470.300 3463.930 2470.560 3464.250 ;
        RECT 2474.440 3463.930 2474.700 3464.250 ;
        RECT 2470.360 3415.370 2470.500 3463.930 ;
        RECT 2470.360 3415.230 2471.420 3415.370 ;
        RECT 2471.280 3367.690 2471.420 3415.230 ;
        RECT 2470.300 3367.370 2470.560 3367.690 ;
        RECT 2471.220 3367.370 2471.480 3367.690 ;
        RECT 2470.360 3346.610 2470.500 3367.370 ;
        RECT 2470.300 3346.290 2470.560 3346.610 ;
        RECT 2471.220 3346.290 2471.480 3346.610 ;
        RECT 2471.280 3332.670 2471.420 3346.290 ;
        RECT 2469.840 3332.350 2470.100 3332.670 ;
        RECT 2471.220 3332.350 2471.480 3332.670 ;
        RECT 2469.900 3284.730 2470.040 3332.350 ;
        RECT 2469.840 3284.410 2470.100 3284.730 ;
        RECT 2470.760 3284.410 2471.020 3284.730 ;
        RECT 2470.820 3250.130 2470.960 3284.410 ;
        RECT 2470.360 3249.990 2470.960 3250.130 ;
        RECT 2470.360 3222.250 2470.500 3249.990 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2959.770 2471.420 2980.030 ;
        RECT 2470.820 2959.630 2471.420 2959.770 ;
        RECT 2470.820 2946.430 2470.960 2959.630 ;
        RECT 2469.380 2946.110 2469.640 2946.430 ;
        RECT 2470.760 2946.110 2471.020 2946.430 ;
        RECT 2469.440 2898.490 2469.580 2946.110 ;
        RECT 2469.380 2898.170 2469.640 2898.490 ;
        RECT 2470.300 2898.170 2470.560 2898.490 ;
        RECT 2470.360 2863.210 2470.500 2898.170 ;
        RECT 2470.360 2863.070 2470.960 2863.210 ;
        RECT 2470.820 2849.530 2470.960 2863.070 ;
        RECT 2470.760 2849.210 2471.020 2849.530 ;
        RECT 2471.680 2849.210 2471.940 2849.530 ;
        RECT 2471.740 2816.210 2471.880 2849.210 ;
        RECT 2471.680 2815.890 2471.940 2816.210 ;
        RECT 2471.680 2815.210 2471.940 2815.530 ;
        RECT 2471.740 2801.330 2471.880 2815.210 ;
        RECT 2471.740 2801.190 2472.800 2801.330 ;
        RECT 2472.660 2766.650 2472.800 2801.190 ;
        RECT 2472.200 2766.510 2472.800 2766.650 ;
        RECT 2472.200 2753.050 2472.340 2766.510 ;
        RECT 2472.200 2752.910 2473.260 2753.050 ;
        RECT 2473.120 2746.365 2473.260 2752.910 ;
        RECT 2458.790 2745.995 2459.070 2746.365 ;
        RECT 2473.050 2745.995 2473.330 2746.365 ;
        RECT 2458.860 2702.650 2459.000 2745.995 ;
        RECT 299.100 2702.330 299.360 2702.650 ;
        RECT 2458.800 2702.330 2459.060 2702.650 ;
        RECT 299.160 2068.405 299.300 2702.330 ;
        RECT 299.090 2068.035 299.370 2068.405 ;
      LAYER via2 ;
        RECT 2458.790 2746.040 2459.070 2746.320 ;
        RECT 2473.050 2746.040 2473.330 2746.320 ;
        RECT 299.090 2068.080 299.370 2068.360 ;
      LAYER met3 ;
        RECT 2458.765 2746.330 2459.095 2746.345 ;
        RECT 2473.025 2746.330 2473.355 2746.345 ;
        RECT 2458.765 2746.030 2473.355 2746.330 ;
        RECT 2458.765 2746.015 2459.095 2746.030 ;
        RECT 2473.025 2746.015 2473.355 2746.030 ;
        RECT 299.065 2068.370 299.395 2068.385 ;
        RECT 300.000 2068.370 304.000 2068.480 ;
        RECT 299.065 2068.070 304.000 2068.370 ;
        RECT 299.065 2068.055 299.395 2068.070 ;
        RECT 300.000 2067.880 304.000 2068.070 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.970 3464.160 2146.290 3464.220 ;
        RECT 2149.650 3464.160 2149.970 3464.220 ;
        RECT 2145.970 3464.020 2149.970 3464.160 ;
        RECT 2145.970 3463.960 2146.290 3464.020 ;
        RECT 2149.650 3463.960 2149.970 3464.020 ;
        RECT 2145.970 3367.260 2146.290 3367.320 ;
        RECT 2147.350 3367.260 2147.670 3367.320 ;
        RECT 2145.970 3367.120 2147.670 3367.260 ;
        RECT 2145.970 3367.060 2146.290 3367.120 ;
        RECT 2147.350 3367.060 2147.670 3367.120 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.430 3042.900 2146.750 3042.960 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.430 3042.760 2147.210 3042.900 ;
        RECT 2146.430 3042.700 2146.750 3042.760 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.430 3008.560 2146.750 3008.620 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.430 3008.420 2148.130 3008.560 ;
        RECT 2146.430 3008.360 2146.750 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2960.080 2148.130 2960.340 ;
        RECT 2147.900 2959.600 2148.040 2960.080 ;
        RECT 2148.270 2959.600 2148.590 2959.660 ;
        RECT 2147.900 2959.460 2148.590 2959.600 ;
        RECT 2148.270 2959.400 2148.590 2959.460 ;
        RECT 2146.430 2915.400 2146.750 2915.460 ;
        RECT 2147.810 2915.400 2148.130 2915.460 ;
        RECT 2146.430 2915.260 2148.130 2915.400 ;
        RECT 2146.430 2915.200 2146.750 2915.260 ;
        RECT 2147.810 2915.200 2148.130 2915.260 ;
        RECT 2146.430 2891.260 2146.750 2891.320 ;
        RECT 2146.890 2891.260 2147.210 2891.320 ;
        RECT 2146.430 2891.120 2147.210 2891.260 ;
        RECT 2146.430 2891.060 2146.750 2891.120 ;
        RECT 2146.890 2891.060 2147.210 2891.120 ;
        RECT 2146.890 2863.040 2147.210 2863.100 ;
        RECT 2148.270 2863.040 2148.590 2863.100 ;
        RECT 2146.890 2862.900 2148.590 2863.040 ;
        RECT 2146.890 2862.840 2147.210 2862.900 ;
        RECT 2148.270 2862.840 2148.590 2862.900 ;
        RECT 2147.350 2801.500 2147.670 2801.560 ;
        RECT 2148.270 2801.500 2148.590 2801.560 ;
        RECT 2147.350 2801.360 2148.590 2801.500 ;
        RECT 2147.350 2801.300 2147.670 2801.360 ;
        RECT 2148.270 2801.300 2148.590 2801.360 ;
        RECT 2146.890 2718.880 2147.210 2718.940 ;
        RECT 2146.890 2718.740 2147.580 2718.880 ;
        RECT 2146.890 2718.680 2147.210 2718.740 ;
        RECT 2147.440 2718.600 2147.580 2718.740 ;
        RECT 2147.350 2718.340 2147.670 2718.600 ;
        RECT 2146.890 2704.940 2147.210 2705.000 ;
        RECT 2147.350 2704.940 2147.670 2705.000 ;
        RECT 2146.890 2704.800 2147.670 2704.940 ;
        RECT 2146.890 2704.740 2147.210 2704.800 ;
        RECT 2147.350 2704.740 2147.670 2704.800 ;
        RECT 299.530 2703.240 299.850 2703.300 ;
        RECT 2146.890 2703.240 2147.210 2703.300 ;
        RECT 299.530 2703.100 2147.210 2703.240 ;
        RECT 299.530 2703.040 299.850 2703.100 ;
        RECT 2146.890 2703.040 2147.210 2703.100 ;
        RECT 297.230 2097.360 297.550 2097.420 ;
        RECT 299.530 2097.360 299.850 2097.420 ;
        RECT 297.230 2097.220 299.850 2097.360 ;
        RECT 297.230 2097.160 297.550 2097.220 ;
        RECT 299.530 2097.160 299.850 2097.220 ;
      LAYER via ;
        RECT 2146.000 3463.960 2146.260 3464.220 ;
        RECT 2149.680 3463.960 2149.940 3464.220 ;
        RECT 2146.000 3367.060 2146.260 3367.320 ;
        RECT 2147.380 3367.060 2147.640 3367.320 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.460 3042.700 2146.720 3042.960 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2146.460 3008.360 2146.720 3008.620 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2960.080 2148.100 2960.340 ;
        RECT 2148.300 2959.400 2148.560 2959.660 ;
        RECT 2146.460 2915.200 2146.720 2915.460 ;
        RECT 2147.840 2915.200 2148.100 2915.460 ;
        RECT 2146.460 2891.060 2146.720 2891.320 ;
        RECT 2146.920 2891.060 2147.180 2891.320 ;
        RECT 2146.920 2862.840 2147.180 2863.100 ;
        RECT 2148.300 2862.840 2148.560 2863.100 ;
        RECT 2147.380 2801.300 2147.640 2801.560 ;
        RECT 2148.300 2801.300 2148.560 2801.560 ;
        RECT 2146.920 2718.680 2147.180 2718.940 ;
        RECT 2147.380 2718.340 2147.640 2718.600 ;
        RECT 2146.920 2704.740 2147.180 2705.000 ;
        RECT 2147.380 2704.740 2147.640 2705.000 ;
        RECT 299.560 2703.040 299.820 2703.300 ;
        RECT 2146.920 2703.040 2147.180 2703.300 ;
        RECT 297.260 2097.160 297.520 2097.420 ;
        RECT 299.560 2097.160 299.820 2097.420 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3517.370 2149.420 3517.600 ;
        RECT 2149.280 3517.230 2149.880 3517.370 ;
        RECT 2149.740 3464.250 2149.880 3517.230 ;
        RECT 2146.000 3463.930 2146.260 3464.250 ;
        RECT 2149.680 3463.930 2149.940 3464.250 ;
        RECT 2146.060 3367.350 2146.200 3463.930 ;
        RECT 2146.000 3367.030 2146.260 3367.350 ;
        RECT 2147.380 3367.030 2147.640 3367.350 ;
        RECT 2147.440 3236.450 2147.580 3367.030 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.460 3042.670 2146.720 3042.990 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2146.520 3008.650 2146.660 3042.670 ;
        RECT 2146.460 3008.330 2146.720 3008.650 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2960.370 2148.040 3008.330 ;
        RECT 2147.840 2960.050 2148.100 2960.370 ;
        RECT 2148.300 2959.370 2148.560 2959.690 ;
        RECT 2148.360 2939.370 2148.500 2959.370 ;
        RECT 2147.900 2939.230 2148.500 2939.370 ;
        RECT 2147.900 2915.490 2148.040 2939.230 ;
        RECT 2146.460 2915.170 2146.720 2915.490 ;
        RECT 2147.840 2915.170 2148.100 2915.490 ;
        RECT 2146.520 2891.350 2146.660 2915.170 ;
        RECT 2146.460 2891.030 2146.720 2891.350 ;
        RECT 2146.920 2891.030 2147.180 2891.350 ;
        RECT 2146.980 2863.130 2147.120 2891.030 ;
        RECT 2146.920 2862.810 2147.180 2863.130 ;
        RECT 2148.300 2862.810 2148.560 2863.130 ;
        RECT 2148.360 2801.590 2148.500 2862.810 ;
        RECT 2147.380 2801.270 2147.640 2801.590 ;
        RECT 2148.300 2801.270 2148.560 2801.590 ;
        RECT 2147.440 2753.050 2147.580 2801.270 ;
        RECT 2146.980 2752.910 2147.580 2753.050 ;
        RECT 2146.980 2718.970 2147.120 2752.910 ;
        RECT 2146.920 2718.650 2147.180 2718.970 ;
        RECT 2147.380 2718.310 2147.640 2718.630 ;
        RECT 2147.440 2705.030 2147.580 2718.310 ;
        RECT 2146.920 2704.710 2147.180 2705.030 ;
        RECT 2147.380 2704.710 2147.640 2705.030 ;
        RECT 2146.980 2703.330 2147.120 2704.710 ;
        RECT 299.560 2703.010 299.820 2703.330 ;
        RECT 2146.920 2703.010 2147.180 2703.330 ;
        RECT 299.620 2097.450 299.760 2703.010 ;
        RECT 297.260 2097.130 297.520 2097.450 ;
        RECT 299.560 2097.130 299.820 2097.450 ;
        RECT 297.320 2096.965 297.460 2097.130 ;
        RECT 297.250 2096.595 297.530 2096.965 ;
      LAYER via2 ;
        RECT 297.250 2096.640 297.530 2096.920 ;
      LAYER met3 ;
        RECT 297.225 2096.930 297.555 2096.945 ;
        RECT 300.000 2096.930 304.000 2097.040 ;
        RECT 297.225 2096.630 304.000 2096.930 ;
        RECT 297.225 2096.615 297.555 2096.630 ;
        RECT 300.000 2096.440 304.000 2096.630 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1822.130 3491.360 1822.450 3491.420 ;
        RECT 1825.350 3491.360 1825.670 3491.420 ;
        RECT 1822.130 3491.220 1825.670 3491.360 ;
        RECT 1822.130 3491.160 1822.450 3491.220 ;
        RECT 1825.350 3491.160 1825.670 3491.220 ;
        RECT 1822.130 3347.000 1822.450 3347.260 ;
        RECT 1822.220 3346.580 1822.360 3347.000 ;
        RECT 1822.130 3346.320 1822.450 3346.580 ;
        RECT 297.230 3253.360 297.550 3253.420 ;
        RECT 1822.590 3253.360 1822.910 3253.420 ;
        RECT 297.230 3253.220 1822.910 3253.360 ;
        RECT 297.230 3253.160 297.550 3253.220 ;
        RECT 1822.590 3253.160 1822.910 3253.220 ;
      LAYER via ;
        RECT 1822.160 3491.160 1822.420 3491.420 ;
        RECT 1825.380 3491.160 1825.640 3491.420 ;
        RECT 1822.160 3347.000 1822.420 3347.260 ;
        RECT 1822.160 3346.320 1822.420 3346.580 ;
        RECT 297.260 3253.160 297.520 3253.420 ;
        RECT 1822.620 3253.160 1822.880 3253.420 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1825.580 3517.370 ;
        RECT 1825.440 3491.450 1825.580 3517.230 ;
        RECT 1822.160 3491.130 1822.420 3491.450 ;
        RECT 1825.380 3491.130 1825.640 3491.450 ;
        RECT 1822.220 3443.250 1822.360 3491.130 ;
        RECT 1821.760 3443.110 1822.360 3443.250 ;
        RECT 1821.760 3442.570 1821.900 3443.110 ;
        RECT 1821.760 3442.430 1822.360 3442.570 ;
        RECT 1822.220 3347.290 1822.360 3442.430 ;
        RECT 1822.160 3346.970 1822.420 3347.290 ;
        RECT 1822.160 3346.290 1822.420 3346.610 ;
        RECT 1822.220 3298.410 1822.360 3346.290 ;
        RECT 1822.220 3298.270 1822.820 3298.410 ;
        RECT 1822.680 3253.450 1822.820 3298.270 ;
        RECT 297.260 3253.130 297.520 3253.450 ;
        RECT 1822.620 3253.130 1822.880 3253.450 ;
        RECT 297.320 2126.205 297.460 3253.130 ;
        RECT 297.250 2125.835 297.530 2126.205 ;
      LAYER via2 ;
        RECT 297.250 2125.880 297.530 2126.160 ;
      LAYER met3 ;
        RECT 297.225 2126.170 297.555 2126.185 ;
        RECT 300.000 2126.170 304.000 2126.280 ;
        RECT 297.225 2125.870 304.000 2126.170 ;
        RECT 297.225 2125.855 297.555 2125.870 ;
        RECT 300.000 2125.680 304.000 2125.870 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.830 3429.480 1498.150 3429.540 ;
        RECT 1500.590 3429.480 1500.910 3429.540 ;
        RECT 1497.830 3429.340 1500.910 3429.480 ;
        RECT 1497.830 3429.280 1498.150 3429.340 ;
        RECT 1500.590 3429.280 1500.910 3429.340 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1498.290 3422.340 1498.610 3422.400 ;
        RECT 1497.830 3422.200 1498.610 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1498.290 3422.140 1498.610 3422.200 ;
        RECT 1498.290 3394.940 1498.610 3395.200 ;
        RECT 1498.380 3394.520 1498.520 3394.940 ;
        RECT 1498.290 3394.260 1498.610 3394.520 ;
        RECT 1498.290 3332.920 1498.610 3332.980 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1498.290 3332.780 1499.990 3332.920 ;
        RECT 1498.290 3332.720 1498.610 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1497.370 3284.300 1497.690 3284.360 ;
        RECT 1498.750 3284.300 1499.070 3284.360 ;
        RECT 1497.370 3284.160 1499.070 3284.300 ;
        RECT 1497.370 3284.100 1497.690 3284.160 ;
        RECT 1498.750 3284.100 1499.070 3284.160 ;
        RECT 1497.370 3236.360 1497.690 3236.420 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1497.370 3236.220 1498.610 3236.360 ;
        RECT 1497.370 3236.160 1497.690 3236.220 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.290 3153.740 1498.610 3153.800 ;
        RECT 1498.750 3153.740 1499.070 3153.800 ;
        RECT 1498.290 3153.600 1499.070 3153.740 ;
        RECT 1498.290 3153.540 1498.610 3153.600 ;
        RECT 1498.750 3153.540 1499.070 3153.600 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1497.830 3042.900 1498.150 3042.960 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1497.830 3042.760 1498.610 3042.900 ;
        RECT 1497.830 3042.700 1498.150 3042.760 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1497.830 3008.560 1498.150 3008.620 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1497.830 3008.420 1499.530 3008.560 ;
        RECT 1497.830 3008.360 1498.150 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1498.290 2994.620 1498.610 2994.680 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1498.290 2994.480 1499.530 2994.620 ;
        RECT 1498.290 2994.420 1498.610 2994.480 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 284.810 2703.580 285.130 2703.640 ;
        RECT 1498.750 2703.580 1499.070 2703.640 ;
        RECT 284.810 2703.440 1499.070 2703.580 ;
        RECT 284.810 2703.380 285.130 2703.440 ;
        RECT 1498.750 2703.380 1499.070 2703.440 ;
      LAYER via ;
        RECT 1497.860 3429.280 1498.120 3429.540 ;
        RECT 1500.620 3429.280 1500.880 3429.540 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1498.320 3422.140 1498.580 3422.400 ;
        RECT 1498.320 3394.940 1498.580 3395.200 ;
        RECT 1498.320 3394.260 1498.580 3394.520 ;
        RECT 1498.320 3332.720 1498.580 3332.980 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1497.400 3284.100 1497.660 3284.360 ;
        RECT 1498.780 3284.100 1499.040 3284.360 ;
        RECT 1497.400 3236.160 1497.660 3236.420 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.320 3153.540 1498.580 3153.800 ;
        RECT 1498.780 3153.540 1499.040 3153.800 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1497.860 3042.700 1498.120 3042.960 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1497.860 3008.360 1498.120 3008.620 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1498.320 2994.420 1498.580 2994.680 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 284.840 2703.380 285.100 2703.640 ;
        RECT 1498.780 2703.380 1499.040 2703.640 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3429.570 1500.820 3517.600 ;
        RECT 1497.860 3429.250 1498.120 3429.570 ;
        RECT 1500.620 3429.250 1500.880 3429.570 ;
        RECT 1497.920 3422.430 1498.060 3429.250 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1498.320 3422.110 1498.580 3422.430 ;
        RECT 1498.380 3395.230 1498.520 3422.110 ;
        RECT 1498.320 3394.910 1498.580 3395.230 ;
        RECT 1498.320 3394.230 1498.580 3394.550 ;
        RECT 1498.380 3333.010 1498.520 3394.230 ;
        RECT 1498.320 3332.690 1498.580 3333.010 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3284.390 1498.980 3298.270 ;
        RECT 1497.400 3284.070 1497.660 3284.390 ;
        RECT 1498.780 3284.070 1499.040 3284.390 ;
        RECT 1497.460 3236.450 1497.600 3284.070 ;
        RECT 1497.400 3236.130 1497.660 3236.450 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.380 3153.830 1498.520 3236.130 ;
        RECT 1498.320 3153.510 1498.580 3153.830 ;
        RECT 1498.780 3153.510 1499.040 3153.830 ;
        RECT 1498.840 3056.930 1498.980 3153.510 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1497.860 3042.670 1498.120 3042.990 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1497.920 3008.650 1498.060 3042.670 ;
        RECT 1497.860 3008.330 1498.120 3008.650 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1498.320 2994.390 1498.580 2994.710 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1498.380 2946.965 1498.520 2994.390 ;
        RECT 1498.310 2946.595 1498.590 2946.965 ;
        RECT 1499.690 2946.595 1499.970 2946.965 ;
        RECT 1499.760 2912.430 1499.900 2946.595 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2815.610 1498.520 2863.070 ;
        RECT 1497.920 2815.470 1498.520 2815.610 ;
        RECT 1497.920 2814.930 1498.060 2815.470 ;
        RECT 1497.920 2814.790 1498.520 2814.930 ;
        RECT 1498.380 2767.330 1498.520 2814.790 ;
        RECT 1498.380 2767.190 1498.980 2767.330 ;
        RECT 1498.840 2703.670 1498.980 2767.190 ;
        RECT 284.840 2703.350 285.100 2703.670 ;
        RECT 1498.780 2703.350 1499.040 2703.670 ;
        RECT 284.900 2155.445 285.040 2703.350 ;
        RECT 284.830 2155.075 285.110 2155.445 ;
      LAYER via2 ;
        RECT 1498.310 2946.640 1498.590 2946.920 ;
        RECT 1499.690 2946.640 1499.970 2946.920 ;
        RECT 284.830 2155.120 285.110 2155.400 ;
      LAYER met3 ;
        RECT 1498.285 2946.930 1498.615 2946.945 ;
        RECT 1499.665 2946.930 1499.995 2946.945 ;
        RECT 1498.285 2946.630 1499.995 2946.930 ;
        RECT 1498.285 2946.615 1498.615 2946.630 ;
        RECT 1499.665 2946.615 1499.995 2946.630 ;
        RECT 284.805 2155.410 285.135 2155.425 ;
        RECT 300.000 2155.410 304.000 2155.520 ;
        RECT 284.805 2155.110 304.000 2155.410 ;
        RECT 284.805 2155.095 285.135 2155.110 ;
        RECT 300.000 2154.920 304.000 2155.110 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.310 324.260 296.630 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 296.310 324.120 2899.310 324.260 ;
        RECT 296.310 324.060 296.630 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 296.340 324.060 296.600 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 296.330 1633.515 296.610 1633.885 ;
        RECT 296.400 324.350 296.540 1633.515 ;
        RECT 296.340 324.030 296.600 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 296.330 1633.560 296.610 1633.840 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 296.305 1633.850 296.635 1633.865 ;
        RECT 300.000 1633.850 304.000 1633.960 ;
        RECT 296.305 1633.550 304.000 1633.850 ;
        RECT 296.305 1633.535 296.635 1633.550 ;
        RECT 300.000 1633.360 304.000 1633.550 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 689.610 3504.960 689.930 3505.020 ;
        RECT 1175.830 3504.960 1176.150 3505.020 ;
        RECT 689.610 3504.820 1176.150 3504.960 ;
        RECT 689.610 3504.760 689.930 3504.820 ;
        RECT 1175.830 3504.760 1176.150 3504.820 ;
        RECT 686.390 3498.500 686.710 3498.560 ;
        RECT 689.610 3498.500 689.930 3498.560 ;
        RECT 686.390 3498.360 689.930 3498.500 ;
        RECT 686.390 3498.300 686.710 3498.360 ;
        RECT 689.610 3498.300 689.930 3498.360 ;
        RECT 284.350 2704.260 284.670 2704.320 ;
        RECT 686.390 2704.260 686.710 2704.320 ;
        RECT 284.350 2704.120 686.710 2704.260 ;
        RECT 284.350 2704.060 284.670 2704.120 ;
        RECT 686.390 2704.060 686.710 2704.120 ;
      LAYER via ;
        RECT 689.640 3504.760 689.900 3505.020 ;
        RECT 1175.860 3504.760 1176.120 3505.020 ;
        RECT 686.420 3498.300 686.680 3498.560 ;
        RECT 689.640 3498.300 689.900 3498.560 ;
        RECT 284.380 2704.060 284.640 2704.320 ;
        RECT 686.420 2704.060 686.680 2704.320 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3505.050 1176.060 3517.600 ;
        RECT 689.640 3504.730 689.900 3505.050 ;
        RECT 1175.860 3504.730 1176.120 3505.050 ;
        RECT 689.700 3498.590 689.840 3504.730 ;
        RECT 686.420 3498.270 686.680 3498.590 ;
        RECT 689.640 3498.270 689.900 3498.590 ;
        RECT 686.480 2704.350 686.620 3498.270 ;
        RECT 284.380 2704.030 284.640 2704.350 ;
        RECT 686.420 2704.030 686.680 2704.350 ;
        RECT 284.440 2184.005 284.580 2704.030 ;
        RECT 284.370 2183.635 284.650 2184.005 ;
      LAYER via2 ;
        RECT 284.370 2183.680 284.650 2183.960 ;
      LAYER met3 ;
        RECT 284.345 2183.970 284.675 2183.985 ;
        RECT 300.000 2183.970 304.000 2184.080 ;
        RECT 284.345 2183.670 304.000 2183.970 ;
        RECT 284.345 2183.655 284.675 2183.670 ;
        RECT 300.000 2183.480 304.000 2183.670 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 850.610 3477.420 850.930 3477.480 ;
        RECT 851.530 3477.420 851.850 3477.480 ;
        RECT 850.610 3477.280 851.850 3477.420 ;
        RECT 850.610 3477.220 850.930 3477.280 ;
        RECT 851.530 3477.220 851.850 3477.280 ;
        RECT 849.230 3429.820 849.550 3429.880 ;
        RECT 850.610 3429.820 850.930 3429.880 ;
        RECT 849.230 3429.680 850.930 3429.820 ;
        RECT 849.230 3429.620 849.550 3429.680 ;
        RECT 850.610 3429.620 850.930 3429.680 ;
        RECT 849.230 3422.340 849.550 3422.400 ;
        RECT 851.070 3422.340 851.390 3422.400 ;
        RECT 849.230 3422.200 851.390 3422.340 ;
        RECT 849.230 3422.140 849.550 3422.200 ;
        RECT 851.070 3422.140 851.390 3422.200 ;
        RECT 849.690 3308.780 850.010 3308.840 ;
        RECT 851.070 3308.780 851.390 3308.840 ;
        RECT 849.690 3308.640 851.390 3308.780 ;
        RECT 849.690 3308.580 850.010 3308.640 ;
        RECT 851.070 3308.580 851.390 3308.640 ;
        RECT 849.690 3284.640 850.010 3284.700 ;
        RECT 850.150 3284.640 850.470 3284.700 ;
        RECT 849.690 3284.500 850.470 3284.640 ;
        RECT 849.690 3284.440 850.010 3284.500 ;
        RECT 850.150 3284.440 850.470 3284.500 ;
        RECT 849.690 3236.360 850.010 3236.420 ;
        RECT 850.150 3236.360 850.470 3236.420 ;
        RECT 849.690 3236.220 850.470 3236.360 ;
        RECT 849.690 3236.160 850.010 3236.220 ;
        RECT 850.150 3236.160 850.470 3236.220 ;
        RECT 849.690 3202.020 850.010 3202.080 ;
        RECT 850.150 3202.020 850.470 3202.080 ;
        RECT 849.690 3201.880 850.470 3202.020 ;
        RECT 849.690 3201.820 850.010 3201.880 ;
        RECT 850.150 3201.820 850.470 3201.880 ;
        RECT 849.230 3153.400 849.550 3153.460 ;
        RECT 850.150 3153.400 850.470 3153.460 ;
        RECT 849.230 3153.260 850.470 3153.400 ;
        RECT 849.230 3153.200 849.550 3153.260 ;
        RECT 850.150 3153.200 850.470 3153.260 ;
        RECT 849.230 3056.840 849.550 3056.900 ;
        RECT 850.150 3056.840 850.470 3056.900 ;
        RECT 849.230 3056.700 850.470 3056.840 ;
        RECT 849.230 3056.640 849.550 3056.700 ;
        RECT 850.150 3056.640 850.470 3056.700 ;
        RECT 849.230 3042.900 849.550 3042.960 ;
        RECT 849.690 3042.900 850.010 3042.960 ;
        RECT 849.230 3042.760 850.010 3042.900 ;
        RECT 849.230 3042.700 849.550 3042.760 ;
        RECT 849.690 3042.700 850.010 3042.760 ;
        RECT 849.230 3008.560 849.550 3008.620 ;
        RECT 850.610 3008.560 850.930 3008.620 ;
        RECT 849.230 3008.420 850.930 3008.560 ;
        RECT 849.230 3008.360 849.550 3008.420 ;
        RECT 850.610 3008.360 850.930 3008.420 ;
        RECT 849.690 2994.620 850.010 2994.680 ;
        RECT 850.610 2994.620 850.930 2994.680 ;
        RECT 849.690 2994.480 850.930 2994.620 ;
        RECT 849.690 2994.420 850.010 2994.480 ;
        RECT 850.610 2994.420 850.930 2994.480 ;
        RECT 849.690 2946.680 850.010 2946.740 ;
        RECT 851.070 2946.680 851.390 2946.740 ;
        RECT 849.690 2946.540 851.390 2946.680 ;
        RECT 849.690 2946.480 850.010 2946.540 ;
        RECT 851.070 2946.480 851.390 2946.540 ;
        RECT 851.070 2912.340 851.390 2912.400 ;
        RECT 850.700 2912.200 851.390 2912.340 ;
        RECT 850.700 2911.720 850.840 2912.200 ;
        RECT 851.070 2912.140 851.390 2912.200 ;
        RECT 850.610 2911.460 850.930 2911.720 ;
        RECT 283.890 2703.920 284.210 2703.980 ;
        RECT 850.150 2703.920 850.470 2703.980 ;
        RECT 283.890 2703.780 850.470 2703.920 ;
        RECT 283.890 2703.720 284.210 2703.780 ;
        RECT 850.150 2703.720 850.470 2703.780 ;
      LAYER via ;
        RECT 850.640 3477.220 850.900 3477.480 ;
        RECT 851.560 3477.220 851.820 3477.480 ;
        RECT 849.260 3429.620 849.520 3429.880 ;
        RECT 850.640 3429.620 850.900 3429.880 ;
        RECT 849.260 3422.140 849.520 3422.400 ;
        RECT 851.100 3422.140 851.360 3422.400 ;
        RECT 849.720 3308.580 849.980 3308.840 ;
        RECT 851.100 3308.580 851.360 3308.840 ;
        RECT 849.720 3284.440 849.980 3284.700 ;
        RECT 850.180 3284.440 850.440 3284.700 ;
        RECT 849.720 3236.160 849.980 3236.420 ;
        RECT 850.180 3236.160 850.440 3236.420 ;
        RECT 849.720 3201.820 849.980 3202.080 ;
        RECT 850.180 3201.820 850.440 3202.080 ;
        RECT 849.260 3153.200 849.520 3153.460 ;
        RECT 850.180 3153.200 850.440 3153.460 ;
        RECT 849.260 3056.640 849.520 3056.900 ;
        RECT 850.180 3056.640 850.440 3056.900 ;
        RECT 849.260 3042.700 849.520 3042.960 ;
        RECT 849.720 3042.700 849.980 3042.960 ;
        RECT 849.260 3008.360 849.520 3008.620 ;
        RECT 850.640 3008.360 850.900 3008.620 ;
        RECT 849.720 2994.420 849.980 2994.680 ;
        RECT 850.640 2994.420 850.900 2994.680 ;
        RECT 849.720 2946.480 849.980 2946.740 ;
        RECT 851.100 2946.480 851.360 2946.740 ;
        RECT 851.100 2912.140 851.360 2912.400 ;
        RECT 850.640 2911.460 850.900 2911.720 ;
        RECT 283.920 2703.720 284.180 2703.980 ;
        RECT 850.180 2703.720 850.440 2703.980 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3477.510 851.760 3517.600 ;
        RECT 850.640 3477.190 850.900 3477.510 ;
        RECT 851.560 3477.190 851.820 3477.510 ;
        RECT 850.700 3429.910 850.840 3477.190 ;
        RECT 849.260 3429.590 849.520 3429.910 ;
        RECT 850.640 3429.590 850.900 3429.910 ;
        RECT 849.320 3422.430 849.460 3429.590 ;
        RECT 849.260 3422.110 849.520 3422.430 ;
        RECT 851.100 3422.110 851.360 3422.430 ;
        RECT 851.160 3308.870 851.300 3422.110 ;
        RECT 849.720 3308.550 849.980 3308.870 ;
        RECT 851.100 3308.550 851.360 3308.870 ;
        RECT 849.780 3284.730 849.920 3308.550 ;
        RECT 849.720 3284.410 849.980 3284.730 ;
        RECT 850.180 3284.410 850.440 3284.730 ;
        RECT 850.240 3236.450 850.380 3284.410 ;
        RECT 849.720 3236.130 849.980 3236.450 ;
        RECT 850.180 3236.130 850.440 3236.450 ;
        RECT 849.780 3202.110 849.920 3236.130 ;
        RECT 849.720 3201.790 849.980 3202.110 ;
        RECT 850.180 3201.790 850.440 3202.110 ;
        RECT 850.240 3153.490 850.380 3201.790 ;
        RECT 849.260 3153.170 849.520 3153.490 ;
        RECT 850.180 3153.170 850.440 3153.490 ;
        RECT 849.320 3152.890 849.460 3153.170 ;
        RECT 849.320 3152.750 849.920 3152.890 ;
        RECT 849.780 3105.290 849.920 3152.750 ;
        RECT 849.780 3105.150 850.380 3105.290 ;
        RECT 850.240 3056.930 850.380 3105.150 ;
        RECT 849.260 3056.610 849.520 3056.930 ;
        RECT 850.180 3056.610 850.440 3056.930 ;
        RECT 849.320 3056.330 849.460 3056.610 ;
        RECT 849.320 3056.190 849.920 3056.330 ;
        RECT 849.780 3042.990 849.920 3056.190 ;
        RECT 849.260 3042.670 849.520 3042.990 ;
        RECT 849.720 3042.670 849.980 3042.990 ;
        RECT 849.320 3008.650 849.460 3042.670 ;
        RECT 849.260 3008.330 849.520 3008.650 ;
        RECT 850.640 3008.330 850.900 3008.650 ;
        RECT 850.700 2994.710 850.840 3008.330 ;
        RECT 849.720 2994.390 849.980 2994.710 ;
        RECT 850.640 2994.390 850.900 2994.710 ;
        RECT 849.780 2946.770 849.920 2994.390 ;
        RECT 849.720 2946.450 849.980 2946.770 ;
        RECT 851.100 2946.450 851.360 2946.770 ;
        RECT 851.160 2912.430 851.300 2946.450 ;
        RECT 851.100 2912.110 851.360 2912.430 ;
        RECT 850.640 2911.430 850.900 2911.750 ;
        RECT 850.700 2863.210 850.840 2911.430 ;
        RECT 849.780 2863.070 850.840 2863.210 ;
        RECT 849.780 2815.610 849.920 2863.070 ;
        RECT 849.320 2815.470 849.920 2815.610 ;
        RECT 849.320 2814.930 849.460 2815.470 ;
        RECT 849.320 2814.790 849.920 2814.930 ;
        RECT 849.780 2767.330 849.920 2814.790 ;
        RECT 849.780 2767.190 850.380 2767.330 ;
        RECT 850.240 2704.010 850.380 2767.190 ;
        RECT 283.920 2703.690 284.180 2704.010 ;
        RECT 850.180 2703.690 850.440 2704.010 ;
        RECT 283.980 2213.245 284.120 2703.690 ;
        RECT 283.910 2212.875 284.190 2213.245 ;
      LAYER via2 ;
        RECT 283.910 2212.920 284.190 2213.200 ;
      LAYER met3 ;
        RECT 283.885 2213.210 284.215 2213.225 ;
        RECT 300.000 2213.210 304.000 2213.320 ;
        RECT 283.885 2212.910 304.000 2213.210 ;
        RECT 283.885 2212.895 284.215 2212.910 ;
        RECT 300.000 2212.720 304.000 2212.910 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 524.930 3491.360 525.250 3491.420 ;
        RECT 527.690 3491.360 528.010 3491.420 ;
        RECT 524.930 3491.220 528.010 3491.360 ;
        RECT 524.930 3491.160 525.250 3491.220 ;
        RECT 527.690 3491.160 528.010 3491.220 ;
        RECT 524.470 3367.600 524.790 3367.660 ;
        RECT 525.390 3367.600 525.710 3367.660 ;
        RECT 524.470 3367.460 525.710 3367.600 ;
        RECT 524.470 3367.400 524.790 3367.460 ;
        RECT 525.390 3367.400 525.710 3367.460 ;
        RECT 288.490 3253.700 288.810 3253.760 ;
        RECT 525.390 3253.700 525.710 3253.760 ;
        RECT 288.490 3253.560 525.710 3253.700 ;
        RECT 288.490 3253.500 288.810 3253.560 ;
        RECT 525.390 3253.500 525.710 3253.560 ;
      LAYER via ;
        RECT 524.960 3491.160 525.220 3491.420 ;
        RECT 527.720 3491.160 527.980 3491.420 ;
        RECT 524.500 3367.400 524.760 3367.660 ;
        RECT 525.420 3367.400 525.680 3367.660 ;
        RECT 288.520 3253.500 288.780 3253.760 ;
        RECT 525.420 3253.500 525.680 3253.760 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3517.370 527.460 3517.600 ;
        RECT 527.320 3517.230 527.920 3517.370 ;
        RECT 527.780 3491.450 527.920 3517.230 ;
        RECT 524.960 3491.130 525.220 3491.450 ;
        RECT 527.720 3491.130 527.980 3491.450 ;
        RECT 525.020 3443.250 525.160 3491.130 ;
        RECT 524.560 3443.110 525.160 3443.250 ;
        RECT 524.560 3415.370 524.700 3443.110 ;
        RECT 524.560 3415.230 525.620 3415.370 ;
        RECT 525.480 3367.690 525.620 3415.230 ;
        RECT 524.500 3367.370 524.760 3367.690 ;
        RECT 525.420 3367.370 525.680 3367.690 ;
        RECT 524.560 3318.810 524.700 3367.370 ;
        RECT 524.560 3318.670 525.620 3318.810 ;
        RECT 525.480 3253.790 525.620 3318.670 ;
        RECT 288.520 3253.470 288.780 3253.790 ;
        RECT 525.420 3253.470 525.680 3253.790 ;
        RECT 288.580 2241.805 288.720 3253.470 ;
        RECT 288.510 2241.435 288.790 2241.805 ;
      LAYER via2 ;
        RECT 288.510 2241.480 288.790 2241.760 ;
      LAYER met3 ;
        RECT 288.485 2241.770 288.815 2241.785 ;
        RECT 300.000 2241.770 304.000 2241.880 ;
        RECT 288.485 2241.470 304.000 2241.770 ;
        RECT 288.485 2241.455 288.815 2241.470 ;
        RECT 300.000 2241.280 304.000 2241.470 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3499.860 202.790 3499.920 ;
        RECT 210.290 3499.860 210.610 3499.920 ;
        RECT 202.470 3499.720 210.610 3499.860 ;
        RECT 202.470 3499.660 202.790 3499.720 ;
        RECT 210.290 3499.660 210.610 3499.720 ;
        RECT 210.290 2276.880 210.610 2276.940 ;
        RECT 282.970 2276.880 283.290 2276.940 ;
        RECT 210.290 2276.740 283.290 2276.880 ;
        RECT 210.290 2276.680 210.610 2276.740 ;
        RECT 282.970 2276.680 283.290 2276.740 ;
      LAYER via ;
        RECT 202.500 3499.660 202.760 3499.920 ;
        RECT 210.320 3499.660 210.580 3499.920 ;
        RECT 210.320 2276.680 210.580 2276.940 ;
        RECT 283.000 2276.680 283.260 2276.940 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3499.950 202.700 3517.600 ;
        RECT 202.500 3499.630 202.760 3499.950 ;
        RECT 210.320 3499.630 210.580 3499.950 ;
        RECT 210.380 2276.970 210.520 3499.630 ;
        RECT 210.320 2276.650 210.580 2276.970 ;
        RECT 283.000 2276.650 283.260 2276.970 ;
        RECT 283.060 2271.045 283.200 2276.650 ;
        RECT 282.990 2270.675 283.270 2271.045 ;
      LAYER via2 ;
        RECT 282.990 2270.720 283.270 2271.000 ;
      LAYER met3 ;
        RECT 282.965 2271.010 283.295 2271.025 ;
        RECT 300.000 2271.010 304.000 2271.120 ;
        RECT 282.965 2270.710 304.000 2271.010 ;
        RECT 282.965 2270.695 283.295 2270.710 ;
        RECT 300.000 2270.520 304.000 2270.710 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2304.420 17.410 2304.480 ;
        RECT 17.090 2304.280 283.660 2304.420 ;
        RECT 17.090 2304.220 17.410 2304.280 ;
        RECT 282.970 2303.740 283.290 2303.800 ;
        RECT 283.520 2303.740 283.660 2304.280 ;
        RECT 282.970 2303.600 283.660 2303.740 ;
        RECT 282.970 2303.540 283.290 2303.600 ;
      LAYER via ;
        RECT 17.120 2304.220 17.380 2304.480 ;
        RECT 283.000 2303.540 283.260 2303.800 ;
      LAYER met2 ;
        RECT 17.110 3411.035 17.390 3411.405 ;
        RECT 17.180 2304.510 17.320 3411.035 ;
        RECT 17.120 2304.190 17.380 2304.510 ;
        RECT 283.000 2303.510 283.260 2303.830 ;
        RECT 283.060 2299.605 283.200 2303.510 ;
        RECT 282.990 2299.235 283.270 2299.605 ;
      LAYER via2 ;
        RECT 17.110 3411.080 17.390 3411.360 ;
        RECT 282.990 2299.280 283.270 2299.560 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.085 3411.370 17.415 3411.385 ;
        RECT -4.800 3411.070 17.415 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.085 3411.055 17.415 3411.070 ;
        RECT 282.965 2299.570 283.295 2299.585 ;
        RECT 300.000 2299.570 304.000 2299.680 ;
        RECT 282.965 2299.270 304.000 2299.570 ;
        RECT 282.965 2299.255 283.295 2299.270 ;
        RECT 300.000 2299.080 304.000 2299.270 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2331.960 17.870 2332.020 ;
        RECT 282.510 2331.960 282.830 2332.020 ;
        RECT 17.550 2331.820 282.830 2331.960 ;
        RECT 17.550 2331.760 17.870 2331.820 ;
        RECT 282.510 2331.760 282.830 2331.820 ;
      LAYER via ;
        RECT 17.580 2331.760 17.840 2332.020 ;
        RECT 282.540 2331.760 282.800 2332.020 ;
      LAYER met2 ;
        RECT 17.570 3124.075 17.850 3124.445 ;
        RECT 17.640 2332.050 17.780 3124.075 ;
        RECT 17.580 2331.730 17.840 2332.050 ;
        RECT 282.540 2331.730 282.800 2332.050 ;
        RECT 282.600 2328.845 282.740 2331.730 ;
        RECT 282.530 2328.475 282.810 2328.845 ;
      LAYER via2 ;
        RECT 17.570 3124.120 17.850 3124.400 ;
        RECT 282.530 2328.520 282.810 2328.800 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.545 3124.410 17.875 3124.425 ;
        RECT -4.800 3124.110 17.875 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.545 3124.095 17.875 3124.110 ;
        RECT 282.505 2328.810 282.835 2328.825 ;
        RECT 300.000 2328.810 304.000 2328.920 ;
        RECT 282.505 2328.510 304.000 2328.810 ;
        RECT 282.505 2328.495 282.835 2328.510 ;
        RECT 300.000 2328.320 304.000 2328.510 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.010 2359.840 18.330 2359.900 ;
        RECT 282.510 2359.840 282.830 2359.900 ;
        RECT 18.010 2359.700 282.830 2359.840 ;
        RECT 18.010 2359.640 18.330 2359.700 ;
        RECT 282.510 2359.640 282.830 2359.700 ;
      LAYER via ;
        RECT 18.040 2359.640 18.300 2359.900 ;
        RECT 282.540 2359.640 282.800 2359.900 ;
      LAYER met2 ;
        RECT 18.030 2836.435 18.310 2836.805 ;
        RECT 18.100 2359.930 18.240 2836.435 ;
        RECT 18.040 2359.610 18.300 2359.930 ;
        RECT 282.540 2359.610 282.800 2359.930 ;
        RECT 282.600 2358.085 282.740 2359.610 ;
        RECT 282.530 2357.715 282.810 2358.085 ;
      LAYER via2 ;
        RECT 18.030 2836.480 18.310 2836.760 ;
        RECT 282.530 2357.760 282.810 2358.040 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 18.005 2836.770 18.335 2836.785 ;
        RECT -4.800 2836.470 18.335 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 18.005 2836.455 18.335 2836.470 ;
        RECT 282.505 2358.050 282.835 2358.065 ;
        RECT 300.000 2358.050 304.000 2358.160 ;
        RECT 282.505 2357.750 304.000 2358.050 ;
        RECT 282.505 2357.735 282.835 2357.750 ;
        RECT 300.000 2357.560 304.000 2357.750 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2387.380 20.630 2387.440 ;
        RECT 282.510 2387.380 282.830 2387.440 ;
        RECT 20.310 2387.240 282.830 2387.380 ;
        RECT 20.310 2387.180 20.630 2387.240 ;
        RECT 282.510 2387.180 282.830 2387.240 ;
      LAYER via ;
        RECT 20.340 2387.180 20.600 2387.440 ;
        RECT 282.540 2387.180 282.800 2387.440 ;
      LAYER met2 ;
        RECT 20.330 2549.475 20.610 2549.845 ;
        RECT 20.400 2387.470 20.540 2549.475 ;
        RECT 20.340 2387.150 20.600 2387.470 ;
        RECT 282.540 2387.150 282.800 2387.470 ;
        RECT 282.600 2386.645 282.740 2387.150 ;
        RECT 282.530 2386.275 282.810 2386.645 ;
      LAYER via2 ;
        RECT 20.330 2549.520 20.610 2549.800 ;
        RECT 282.530 2386.320 282.810 2386.600 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 20.305 2549.810 20.635 2549.825 ;
        RECT -4.800 2549.510 20.635 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 20.305 2549.495 20.635 2549.510 ;
        RECT 282.505 2386.610 282.835 2386.625 ;
        RECT 300.000 2386.610 304.000 2386.720 ;
        RECT 282.505 2386.310 304.000 2386.610 ;
        RECT 282.505 2386.295 282.835 2386.310 ;
        RECT 300.000 2386.120 304.000 2386.310 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 2262.940 17.410 2263.000 ;
        RECT 282.970 2262.940 283.290 2263.000 ;
        RECT 17.090 2262.800 283.290 2262.940 ;
        RECT 17.090 2262.740 17.410 2262.800 ;
        RECT 282.970 2262.740 283.290 2262.800 ;
      LAYER via ;
        RECT 17.120 2262.740 17.380 2263.000 ;
        RECT 283.000 2262.740 283.260 2263.000 ;
      LAYER met2 ;
        RECT 282.990 2415.515 283.270 2415.885 ;
        RECT 283.060 2304.250 283.200 2415.515 ;
        RECT 282.140 2304.110 283.200 2304.250 ;
        RECT 282.140 2298.130 282.280 2304.110 ;
        RECT 282.140 2297.990 283.200 2298.130 ;
        RECT 283.060 2291.330 283.200 2297.990 ;
        RECT 282.600 2291.190 283.200 2291.330 ;
        RECT 282.600 2289.290 282.740 2291.190 ;
        RECT 282.600 2289.150 283.200 2289.290 ;
        RECT 283.060 2284.530 283.200 2289.150 ;
        RECT 282.600 2284.390 283.200 2284.530 ;
        RECT 282.600 2270.250 282.740 2284.390 ;
        RECT 282.600 2270.110 283.200 2270.250 ;
        RECT 283.060 2263.030 283.200 2270.110 ;
        RECT 17.120 2262.710 17.380 2263.030 ;
        RECT 283.000 2262.710 283.260 2263.030 ;
        RECT 17.180 2262.205 17.320 2262.710 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
      LAYER via2 ;
        RECT 282.990 2415.560 283.270 2415.840 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
      LAYER met3 ;
        RECT 282.965 2415.850 283.295 2415.865 ;
        RECT 300.000 2415.850 304.000 2415.960 ;
        RECT 282.965 2415.550 304.000 2415.850 ;
        RECT 282.965 2415.535 283.295 2415.550 ;
        RECT 300.000 2415.360 304.000 2415.550 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 283.430 2408.800 283.750 2408.860 ;
        RECT 283.430 2408.660 284.120 2408.800 ;
        RECT 283.430 2408.600 283.750 2408.660 ;
        RECT 283.430 2405.740 283.750 2405.800 ;
        RECT 283.980 2405.740 284.120 2408.660 ;
        RECT 283.430 2405.600 284.120 2405.740 ;
        RECT 283.430 2405.540 283.750 2405.600 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 283.430 1980.060 283.750 1980.120 ;
        RECT 15.710 1979.920 283.750 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 283.430 1979.860 283.750 1979.920 ;
      LAYER via ;
        RECT 283.460 2408.600 283.720 2408.860 ;
        RECT 283.460 2405.540 283.720 2405.800 ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 283.460 1979.860 283.720 1980.120 ;
      LAYER met2 ;
        RECT 282.990 2444.075 283.270 2444.445 ;
        RECT 283.060 2421.210 283.200 2444.075 ;
        RECT 283.060 2421.070 283.660 2421.210 ;
        RECT 283.520 2408.890 283.660 2421.070 ;
        RECT 283.460 2408.570 283.720 2408.890 ;
        RECT 283.460 2405.510 283.720 2405.830 ;
        RECT 283.520 1980.150 283.660 2405.510 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 283.460 1979.830 283.720 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 282.990 2444.120 283.270 2444.400 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 282.965 2444.410 283.295 2444.425 ;
        RECT 300.000 2444.410 304.000 2444.520 ;
        RECT 282.965 2444.110 304.000 2444.410 ;
        RECT 282.965 2444.095 283.295 2444.110 ;
        RECT 300.000 2443.920 304.000 2444.110 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 295.850 558.860 296.170 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 295.850 558.720 2899.310 558.860 ;
        RECT 295.850 558.660 296.170 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 295.880 558.660 296.140 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 295.870 1662.755 296.150 1663.125 ;
        RECT 295.940 558.950 296.080 1662.755 ;
        RECT 295.880 558.630 296.140 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 295.870 1662.800 296.150 1663.080 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 295.845 1663.090 296.175 1663.105 ;
        RECT 300.000 1663.090 304.000 1663.200 ;
        RECT 295.845 1662.790 304.000 1663.090 ;
        RECT 295.845 1662.775 296.175 1662.790 ;
        RECT 300.000 1662.600 304.000 1662.790 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 287.110 1690.380 287.430 1690.440 ;
        RECT 17.090 1690.240 287.430 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 287.110 1690.180 287.430 1690.240 ;
      LAYER via ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 287.140 1690.180 287.400 1690.440 ;
      LAYER met2 ;
        RECT 287.130 2473.315 287.410 2473.685 ;
        RECT 287.200 1690.470 287.340 2473.315 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 287.140 1690.150 287.400 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 287.130 2473.360 287.410 2473.640 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT 287.105 2473.650 287.435 2473.665 ;
        RECT 300.000 2473.650 304.000 2473.760 ;
        RECT 287.105 2473.350 304.000 2473.650 ;
        RECT 287.105 2473.335 287.435 2473.350 ;
        RECT 300.000 2473.160 304.000 2473.350 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 286.650 1476.520 286.970 1476.580 ;
        RECT 17.090 1476.380 286.970 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 286.650 1476.320 286.970 1476.380 ;
      LAYER via ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 286.680 1476.320 286.940 1476.580 ;
      LAYER met2 ;
        RECT 286.670 2501.875 286.950 2502.245 ;
        RECT 286.740 1476.610 286.880 2501.875 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 286.680 1476.290 286.940 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 286.670 2501.920 286.950 2502.200 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 286.645 2502.210 286.975 2502.225 ;
        RECT 300.000 2502.210 304.000 2502.320 ;
        RECT 286.645 2501.910 304.000 2502.210 ;
        RECT 286.645 2501.895 286.975 2501.910 ;
        RECT 300.000 2501.720 304.000 2501.910 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1262.660 17.410 1262.720 ;
        RECT 286.190 1262.660 286.510 1262.720 ;
        RECT 17.090 1262.520 286.510 1262.660 ;
        RECT 17.090 1262.460 17.410 1262.520 ;
        RECT 286.190 1262.460 286.510 1262.520 ;
      LAYER via ;
        RECT 17.120 1262.460 17.380 1262.720 ;
        RECT 286.220 1262.460 286.480 1262.720 ;
      LAYER met2 ;
        RECT 286.210 2531.115 286.490 2531.485 ;
        RECT 286.280 1262.750 286.420 2531.115 ;
        RECT 17.120 1262.430 17.380 1262.750 ;
        RECT 286.220 1262.430 286.480 1262.750 ;
        RECT 17.180 1256.485 17.320 1262.430 ;
        RECT 17.110 1256.115 17.390 1256.485 ;
      LAYER via2 ;
        RECT 286.210 2531.160 286.490 2531.440 ;
        RECT 17.110 1256.160 17.390 1256.440 ;
      LAYER met3 ;
        RECT 286.185 2531.450 286.515 2531.465 ;
        RECT 300.000 2531.450 304.000 2531.560 ;
        RECT 286.185 2531.150 304.000 2531.450 ;
        RECT 286.185 2531.135 286.515 2531.150 ;
        RECT 300.000 2530.960 304.000 2531.150 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.085 1256.450 17.415 1256.465 ;
        RECT -4.800 1256.150 17.415 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.085 1256.135 17.415 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 25.370 2560.100 25.690 2560.160 ;
        RECT 287.110 2560.100 287.430 2560.160 ;
        RECT 25.370 2559.960 287.430 2560.100 ;
        RECT 25.370 2559.900 25.690 2559.960 ;
        RECT 287.110 2559.900 287.430 2559.960 ;
        RECT 13.870 1040.980 14.190 1041.040 ;
        RECT 25.370 1040.980 25.690 1041.040 ;
        RECT 13.870 1040.840 25.690 1040.980 ;
        RECT 13.870 1040.780 14.190 1040.840 ;
        RECT 25.370 1040.780 25.690 1040.840 ;
      LAYER via ;
        RECT 25.400 2559.900 25.660 2560.160 ;
        RECT 287.140 2559.900 287.400 2560.160 ;
        RECT 13.900 1040.780 14.160 1041.040 ;
        RECT 25.400 1040.780 25.660 1041.040 ;
      LAYER met2 ;
        RECT 287.130 2560.355 287.410 2560.725 ;
        RECT 287.200 2560.190 287.340 2560.355 ;
        RECT 25.400 2559.870 25.660 2560.190 ;
        RECT 287.140 2559.870 287.400 2560.190 ;
        RECT 25.460 1041.070 25.600 2559.870 ;
        RECT 13.900 1040.925 14.160 1041.070 ;
        RECT 13.890 1040.555 14.170 1040.925 ;
        RECT 25.400 1040.750 25.660 1041.070 ;
      LAYER via2 ;
        RECT 287.130 2560.400 287.410 2560.680 ;
        RECT 13.890 1040.600 14.170 1040.880 ;
      LAYER met3 ;
        RECT 287.105 2560.690 287.435 2560.705 ;
        RECT 300.000 2560.690 304.000 2560.800 ;
        RECT 287.105 2560.390 304.000 2560.690 ;
        RECT 287.105 2560.375 287.435 2560.390 ;
        RECT 300.000 2560.200 304.000 2560.390 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 13.865 1040.890 14.195 1040.905 ;
        RECT -4.800 1040.590 14.195 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 13.865 1040.575 14.195 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 2587.640 25.230 2587.700 ;
        RECT 287.110 2587.640 287.430 2587.700 ;
        RECT 24.910 2587.500 287.430 2587.640 ;
        RECT 24.910 2587.440 25.230 2587.500 ;
        RECT 287.110 2587.440 287.430 2587.500 ;
        RECT 13.870 827.460 14.190 827.520 ;
        RECT 24.910 827.460 25.230 827.520 ;
        RECT 13.870 827.320 25.230 827.460 ;
        RECT 13.870 827.260 14.190 827.320 ;
        RECT 24.910 827.260 25.230 827.320 ;
      LAYER via ;
        RECT 24.940 2587.440 25.200 2587.700 ;
        RECT 287.140 2587.440 287.400 2587.700 ;
        RECT 13.900 827.260 14.160 827.520 ;
        RECT 24.940 827.260 25.200 827.520 ;
      LAYER met2 ;
        RECT 287.130 2588.915 287.410 2589.285 ;
        RECT 287.200 2587.730 287.340 2588.915 ;
        RECT 24.940 2587.410 25.200 2587.730 ;
        RECT 287.140 2587.410 287.400 2587.730 ;
        RECT 25.000 827.550 25.140 2587.410 ;
        RECT 13.900 827.230 14.160 827.550 ;
        RECT 24.940 827.230 25.200 827.550 ;
        RECT 13.960 825.365 14.100 827.230 ;
        RECT 13.890 824.995 14.170 825.365 ;
      LAYER via2 ;
        RECT 287.130 2588.960 287.410 2589.240 ;
        RECT 13.890 825.040 14.170 825.320 ;
      LAYER met3 ;
        RECT 287.105 2589.250 287.435 2589.265 ;
        RECT 300.000 2589.250 304.000 2589.360 ;
        RECT 287.105 2588.950 304.000 2589.250 ;
        RECT 287.105 2588.935 287.435 2588.950 ;
        RECT 300.000 2588.760 304.000 2588.950 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 13.865 825.330 14.195 825.345 ;
        RECT -4.800 825.030 14.195 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 13.865 825.015 14.195 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 2615.180 24.770 2615.240 ;
        RECT 287.110 2615.180 287.430 2615.240 ;
        RECT 24.450 2615.040 287.430 2615.180 ;
        RECT 24.450 2614.980 24.770 2615.040 ;
        RECT 287.110 2614.980 287.430 2615.040 ;
        RECT 13.870 611.900 14.190 611.960 ;
        RECT 24.450 611.900 24.770 611.960 ;
        RECT 13.870 611.760 24.770 611.900 ;
        RECT 13.870 611.700 14.190 611.760 ;
        RECT 24.450 611.700 24.770 611.760 ;
      LAYER via ;
        RECT 24.480 2614.980 24.740 2615.240 ;
        RECT 287.140 2614.980 287.400 2615.240 ;
        RECT 13.900 611.700 14.160 611.960 ;
        RECT 24.480 611.700 24.740 611.960 ;
      LAYER met2 ;
        RECT 287.130 2618.155 287.410 2618.525 ;
        RECT 287.200 2615.270 287.340 2618.155 ;
        RECT 24.480 2614.950 24.740 2615.270 ;
        RECT 287.140 2614.950 287.400 2615.270 ;
        RECT 24.540 611.990 24.680 2614.950 ;
        RECT 13.900 611.670 14.160 611.990 ;
        RECT 24.480 611.670 24.740 611.990 ;
        RECT 13.960 610.485 14.100 611.670 ;
        RECT 13.890 610.115 14.170 610.485 ;
      LAYER via2 ;
        RECT 287.130 2618.200 287.410 2618.480 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT 287.105 2618.490 287.435 2618.505 ;
        RECT 300.000 2618.490 304.000 2618.600 ;
        RECT 287.105 2618.190 304.000 2618.490 ;
        RECT 287.105 2618.175 287.435 2618.190 ;
        RECT 300.000 2618.000 304.000 2618.190 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.800 610.150 14.195 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 23.990 2643.060 24.310 2643.120 ;
        RECT 287.110 2643.060 287.430 2643.120 ;
        RECT 23.990 2642.920 287.430 2643.060 ;
        RECT 23.990 2642.860 24.310 2642.920 ;
        RECT 287.110 2642.860 287.430 2642.920 ;
        RECT 13.870 395.320 14.190 395.380 ;
        RECT 23.990 395.320 24.310 395.380 ;
        RECT 13.870 395.180 24.310 395.320 ;
        RECT 13.870 395.120 14.190 395.180 ;
        RECT 23.990 395.120 24.310 395.180 ;
      LAYER via ;
        RECT 24.020 2642.860 24.280 2643.120 ;
        RECT 287.140 2642.860 287.400 2643.120 ;
        RECT 13.900 395.120 14.160 395.380 ;
        RECT 24.020 395.120 24.280 395.380 ;
      LAYER met2 ;
        RECT 287.130 2646.715 287.410 2647.085 ;
        RECT 287.200 2643.150 287.340 2646.715 ;
        RECT 24.020 2642.830 24.280 2643.150 ;
        RECT 287.140 2642.830 287.400 2643.150 ;
        RECT 24.080 395.410 24.220 2642.830 ;
        RECT 13.900 395.090 14.160 395.410 ;
        RECT 24.020 395.090 24.280 395.410 ;
        RECT 13.960 394.925 14.100 395.090 ;
        RECT 13.890 394.555 14.170 394.925 ;
      LAYER via2 ;
        RECT 287.130 2646.760 287.410 2647.040 ;
        RECT 13.890 394.600 14.170 394.880 ;
      LAYER met3 ;
        RECT 287.105 2647.050 287.435 2647.065 ;
        RECT 300.000 2647.050 304.000 2647.160 ;
        RECT 287.105 2646.750 304.000 2647.050 ;
        RECT 287.105 2646.735 287.435 2646.750 ;
        RECT 300.000 2646.560 304.000 2646.750 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 13.865 394.890 14.195 394.905 ;
        RECT -4.800 394.590 14.195 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 13.865 394.575 14.195 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 2670.600 86.410 2670.660 ;
        RECT 287.110 2670.600 287.430 2670.660 ;
        RECT 86.090 2670.460 287.430 2670.600 ;
        RECT 86.090 2670.400 86.410 2670.460 ;
        RECT 287.110 2670.400 287.430 2670.460 ;
        RECT 17.090 179.420 17.410 179.480 ;
        RECT 86.090 179.420 86.410 179.480 ;
        RECT 17.090 179.280 86.410 179.420 ;
        RECT 17.090 179.220 17.410 179.280 ;
        RECT 86.090 179.220 86.410 179.280 ;
      LAYER via ;
        RECT 86.120 2670.400 86.380 2670.660 ;
        RECT 287.140 2670.400 287.400 2670.660 ;
        RECT 17.120 179.220 17.380 179.480 ;
        RECT 86.120 179.220 86.380 179.480 ;
      LAYER met2 ;
        RECT 287.130 2675.955 287.410 2676.325 ;
        RECT 287.200 2670.690 287.340 2675.955 ;
        RECT 86.120 2670.370 86.380 2670.690 ;
        RECT 287.140 2670.370 287.400 2670.690 ;
        RECT 86.180 179.510 86.320 2670.370 ;
        RECT 17.120 179.365 17.380 179.510 ;
        RECT 17.110 178.995 17.390 179.365 ;
        RECT 86.120 179.190 86.380 179.510 ;
      LAYER via2 ;
        RECT 287.130 2676.000 287.410 2676.280 ;
        RECT 17.110 179.040 17.390 179.320 ;
      LAYER met3 ;
        RECT 287.105 2676.290 287.435 2676.305 ;
        RECT 300.000 2676.290 304.000 2676.400 ;
        RECT 287.105 2675.990 304.000 2676.290 ;
        RECT 287.105 2675.975 287.435 2675.990 ;
        RECT 300.000 2675.800 304.000 2675.990 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.085 179.330 17.415 179.345 ;
        RECT -4.800 179.030 17.415 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.085 179.015 17.415 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 295.390 793.460 295.710 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 295.390 793.320 2899.310 793.460 ;
        RECT 295.390 793.260 295.710 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 295.420 793.260 295.680 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 295.410 1691.315 295.690 1691.685 ;
        RECT 295.480 793.550 295.620 1691.315 ;
        RECT 295.420 793.230 295.680 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 295.410 1691.360 295.690 1691.640 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 295.385 1691.650 295.715 1691.665 ;
        RECT 300.000 1691.650 304.000 1691.760 ;
        RECT 295.385 1691.350 304.000 1691.650 ;
        RECT 295.385 1691.335 295.715 1691.350 ;
        RECT 300.000 1691.160 304.000 1691.350 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.770 1028.060 297.090 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 296.770 1027.920 2899.310 1028.060 ;
        RECT 296.770 1027.860 297.090 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 296.800 1027.860 297.060 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 296.790 1720.555 297.070 1720.925 ;
        RECT 296.860 1028.150 297.000 1720.555 ;
        RECT 296.800 1027.830 297.060 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 296.790 1720.600 297.070 1720.880 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 296.765 1720.890 297.095 1720.905 ;
        RECT 300.000 1720.890 304.000 1721.000 ;
        RECT 296.765 1720.590 304.000 1720.890 ;
        RECT 296.765 1720.575 297.095 1720.590 ;
        RECT 300.000 1720.400 304.000 1720.590 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 297.230 1262.660 297.550 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 297.230 1262.520 2899.310 1262.660 ;
        RECT 297.230 1262.460 297.550 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 297.260 1262.460 297.520 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 297.250 1749.115 297.530 1749.485 ;
        RECT 297.320 1262.750 297.460 1749.115 ;
        RECT 297.260 1262.430 297.520 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 297.250 1749.160 297.530 1749.440 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 297.225 1749.450 297.555 1749.465 ;
        RECT 300.000 1749.450 304.000 1749.560 ;
        RECT 297.225 1749.150 304.000 1749.450 ;
        RECT 297.225 1749.135 297.555 1749.150 ;
        RECT 300.000 1748.960 304.000 1749.150 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 283.890 1497.260 284.210 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 283.890 1497.120 2899.310 1497.260 ;
        RECT 283.890 1497.060 284.210 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 283.920 1497.060 284.180 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 283.910 1778.355 284.190 1778.725 ;
        RECT 283.980 1497.350 284.120 1778.355 ;
        RECT 283.920 1497.030 284.180 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 283.910 1778.400 284.190 1778.680 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 283.885 1778.690 284.215 1778.705 ;
        RECT 300.000 1778.690 304.000 1778.800 ;
        RECT 283.885 1778.390 304.000 1778.690 ;
        RECT 283.885 1778.375 284.215 1778.390 ;
        RECT 300.000 1778.200 304.000 1778.390 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.970 1653.320 283.290 1653.380 ;
        RECT 284.350 1653.320 284.670 1653.380 ;
        RECT 282.970 1653.180 284.670 1653.320 ;
        RECT 282.970 1653.120 283.290 1653.180 ;
        RECT 284.350 1653.120 284.670 1653.180 ;
        RECT 282.970 1627.480 283.290 1627.540 ;
        RECT 289.870 1627.480 290.190 1627.540 ;
        RECT 282.970 1627.340 290.190 1627.480 ;
        RECT 282.970 1627.280 283.290 1627.340 ;
        RECT 289.870 1627.280 290.190 1627.340 ;
        RECT 289.870 1603.680 290.190 1603.740 ;
        RECT 2900.830 1603.680 2901.150 1603.740 ;
        RECT 289.870 1603.540 2901.150 1603.680 ;
        RECT 289.870 1603.480 290.190 1603.540 ;
        RECT 2900.830 1603.480 2901.150 1603.540 ;
      LAYER via ;
        RECT 283.000 1653.120 283.260 1653.380 ;
        RECT 284.380 1653.120 284.640 1653.380 ;
        RECT 283.000 1627.280 283.260 1627.540 ;
        RECT 289.900 1627.280 290.160 1627.540 ;
        RECT 289.900 1603.480 290.160 1603.740 ;
        RECT 2900.860 1603.480 2901.120 1603.740 ;
      LAYER met2 ;
        RECT 284.370 1807.595 284.650 1807.965 ;
        RECT 284.440 1653.410 284.580 1807.595 ;
        RECT 2900.850 1730.075 2901.130 1730.445 ;
        RECT 283.000 1653.090 283.260 1653.410 ;
        RECT 284.380 1653.090 284.640 1653.410 ;
        RECT 283.060 1627.570 283.200 1653.090 ;
        RECT 283.000 1627.250 283.260 1627.570 ;
        RECT 289.900 1627.250 290.160 1627.570 ;
        RECT 289.960 1624.930 290.100 1627.250 ;
        RECT 289.500 1624.790 290.100 1624.930 ;
        RECT 289.500 1605.890 289.640 1624.790 ;
        RECT 289.500 1605.750 290.100 1605.890 ;
        RECT 289.960 1603.770 290.100 1605.750 ;
        RECT 2900.920 1603.770 2901.060 1730.075 ;
        RECT 289.900 1603.450 290.160 1603.770 ;
        RECT 2900.860 1603.450 2901.120 1603.770 ;
      LAYER via2 ;
        RECT 284.370 1807.640 284.650 1807.920 ;
        RECT 2900.850 1730.120 2901.130 1730.400 ;
      LAYER met3 ;
        RECT 284.345 1807.930 284.675 1807.945 ;
        RECT 300.000 1807.930 304.000 1808.040 ;
        RECT 284.345 1807.630 304.000 1807.930 ;
        RECT 284.345 1807.615 284.675 1807.630 ;
        RECT 300.000 1807.440 304.000 1807.630 ;
        RECT 2900.825 1730.410 2901.155 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2900.825 1730.110 2924.800 1730.410 ;
        RECT 2900.825 1730.095 2901.155 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 287.570 1603.340 287.890 1603.400 ;
        RECT 2903.590 1603.340 2903.910 1603.400 ;
        RECT 287.570 1603.200 2903.910 1603.340 ;
        RECT 287.570 1603.140 287.890 1603.200 ;
        RECT 2903.590 1603.140 2903.910 1603.200 ;
      LAYER via ;
        RECT 287.600 1603.140 287.860 1603.400 ;
        RECT 2903.620 1603.140 2903.880 1603.400 ;
      LAYER met2 ;
        RECT 2903.610 1964.675 2903.890 1965.045 ;
        RECT 288.050 1836.155 288.330 1836.525 ;
        RECT 288.120 1625.610 288.260 1836.155 ;
        RECT 287.660 1625.470 288.260 1625.610 ;
        RECT 287.660 1603.430 287.800 1625.470 ;
        RECT 2903.680 1603.430 2903.820 1964.675 ;
        RECT 287.600 1603.110 287.860 1603.430 ;
        RECT 2903.620 1603.110 2903.880 1603.430 ;
      LAYER via2 ;
        RECT 2903.610 1964.720 2903.890 1965.000 ;
        RECT 288.050 1836.200 288.330 1836.480 ;
      LAYER met3 ;
        RECT 2903.585 1965.010 2903.915 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2903.585 1964.710 2924.800 1965.010 ;
        RECT 2903.585 1964.695 2903.915 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 288.025 1836.490 288.355 1836.505 ;
        RECT 300.000 1836.490 304.000 1836.600 ;
        RECT 288.025 1836.190 304.000 1836.490 ;
        RECT 288.025 1836.175 288.355 1836.190 ;
        RECT 300.000 1836.000 304.000 1836.190 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 288.490 1625.440 288.810 1625.500 ;
        RECT 298.150 1625.440 298.470 1625.500 ;
        RECT 288.490 1625.300 298.470 1625.440 ;
        RECT 288.490 1625.240 288.810 1625.300 ;
        RECT 298.150 1625.240 298.470 1625.300 ;
        RECT 298.150 1599.940 298.470 1600.000 ;
        RECT 2902.210 1599.940 2902.530 1600.000 ;
        RECT 298.150 1599.800 2902.530 1599.940 ;
        RECT 298.150 1599.740 298.470 1599.800 ;
        RECT 2902.210 1599.740 2902.530 1599.800 ;
      LAYER via ;
        RECT 288.520 1625.240 288.780 1625.500 ;
        RECT 298.180 1625.240 298.440 1625.500 ;
        RECT 298.180 1599.740 298.440 1600.000 ;
        RECT 2902.240 1599.740 2902.500 1600.000 ;
      LAYER met2 ;
        RECT 2902.230 2199.275 2902.510 2199.645 ;
        RECT 288.510 1865.395 288.790 1865.765 ;
        RECT 288.580 1625.530 288.720 1865.395 ;
        RECT 288.520 1625.210 288.780 1625.530 ;
        RECT 298.180 1625.210 298.440 1625.530 ;
        RECT 298.240 1600.030 298.380 1625.210 ;
        RECT 2902.300 1600.030 2902.440 2199.275 ;
        RECT 298.180 1599.710 298.440 1600.030 ;
        RECT 2902.240 1599.710 2902.500 1600.030 ;
      LAYER via2 ;
        RECT 2902.230 2199.320 2902.510 2199.600 ;
        RECT 288.510 1865.440 288.790 1865.720 ;
      LAYER met3 ;
        RECT 2902.205 2199.610 2902.535 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2902.205 2199.310 2924.800 2199.610 ;
        RECT 2902.205 2199.295 2902.535 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 288.485 1865.730 288.815 1865.745 ;
        RECT 300.000 1865.730 304.000 1865.840 ;
        RECT 288.485 1865.430 304.000 1865.730 ;
        RECT 288.485 1865.415 288.815 1865.430 ;
        RECT 300.000 1865.240 304.000 1865.430 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.490 206.960 288.810 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 288.490 206.820 2901.150 206.960 ;
        RECT 288.490 206.760 288.810 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 288.520 206.760 288.780 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 288.510 1614.475 288.790 1614.845 ;
        RECT 288.580 207.050 288.720 1614.475 ;
        RECT 288.520 206.730 288.780 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 288.510 1614.520 288.790 1614.800 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 288.485 1614.810 288.815 1614.825 ;
        RECT 300.000 1614.810 304.000 1614.920 ;
        RECT 288.485 1614.510 304.000 1614.810 ;
        RECT 288.485 1614.495 288.815 1614.510 ;
        RECT 300.000 1614.320 304.000 1614.510 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 287.570 2698.140 287.890 2698.200 ;
        RECT 2904.050 2698.140 2904.370 2698.200 ;
        RECT 287.570 2698.000 2904.370 2698.140 ;
        RECT 287.570 2697.940 287.890 2698.000 ;
        RECT 2904.050 2697.940 2904.370 2698.000 ;
      LAYER via ;
        RECT 287.600 2697.940 287.860 2698.200 ;
        RECT 2904.080 2697.940 2904.340 2698.200 ;
      LAYER met2 ;
        RECT 287.600 2697.910 287.860 2698.230 ;
        RECT 2904.080 2697.910 2904.340 2698.230 ;
        RECT 287.660 1903.845 287.800 2697.910 ;
        RECT 2904.140 2551.885 2904.280 2697.910 ;
        RECT 2904.070 2551.515 2904.350 2551.885 ;
        RECT 287.590 1903.475 287.870 1903.845 ;
      LAYER via2 ;
        RECT 2904.070 2551.560 2904.350 2551.840 ;
        RECT 287.590 1903.520 287.870 1903.800 ;
      LAYER met3 ;
        RECT 2904.045 2551.850 2904.375 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2904.045 2551.550 2924.800 2551.850 ;
        RECT 2904.045 2551.535 2904.375 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 287.565 1903.810 287.895 1903.825 ;
        RECT 300.000 1903.810 304.000 1903.920 ;
        RECT 287.565 1903.510 304.000 1903.810 ;
        RECT 287.565 1903.495 287.895 1903.510 ;
        RECT 300.000 1903.320 304.000 1903.510 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 291.250 2781.100 291.570 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 291.250 2780.960 2901.150 2781.100 ;
        RECT 291.250 2780.900 291.570 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 291.280 2780.900 291.540 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 291.280 2780.870 291.540 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 291.340 1933.085 291.480 2780.870 ;
        RECT 291.270 1932.715 291.550 1933.085 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 291.270 1932.760 291.550 1933.040 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 291.245 1933.050 291.575 1933.065 ;
        RECT 300.000 1933.050 304.000 1933.160 ;
        RECT 291.245 1932.750 304.000 1933.050 ;
        RECT 291.245 1932.735 291.575 1932.750 ;
        RECT 300.000 1932.560 304.000 1932.750 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 290.790 2701.200 291.110 2701.260 ;
        RECT 2902.210 2701.200 2902.530 2701.260 ;
        RECT 290.790 2701.060 2902.530 2701.200 ;
        RECT 290.790 2701.000 291.110 2701.060 ;
        RECT 2902.210 2701.000 2902.530 2701.060 ;
      LAYER via ;
        RECT 290.820 2701.000 291.080 2701.260 ;
        RECT 2902.240 2701.000 2902.500 2701.260 ;
      LAYER met2 ;
        RECT 2902.230 3020.715 2902.510 3021.085 ;
        RECT 2902.300 2701.290 2902.440 3020.715 ;
        RECT 290.820 2700.970 291.080 2701.290 ;
        RECT 2902.240 2700.970 2902.500 2701.290 ;
        RECT 290.880 1962.325 291.020 2700.970 ;
        RECT 290.810 1961.955 291.090 1962.325 ;
      LAYER via2 ;
        RECT 2902.230 3020.760 2902.510 3021.040 ;
        RECT 290.810 1962.000 291.090 1962.280 ;
      LAYER met3 ;
        RECT 2902.205 3021.050 2902.535 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2902.205 3020.750 2924.800 3021.050 ;
        RECT 2902.205 3020.735 2902.535 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 290.785 1962.290 291.115 1962.305 ;
        RECT 300.000 1962.290 304.000 1962.400 ;
        RECT 290.785 1961.990 304.000 1962.290 ;
        RECT 290.785 1961.975 291.115 1961.990 ;
        RECT 300.000 1961.800 304.000 1961.990 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1835.470 3254.040 1835.790 3254.100 ;
        RECT 1852.030 3254.040 1852.350 3254.100 ;
        RECT 1835.470 3253.900 1852.350 3254.040 ;
        RECT 1835.470 3253.840 1835.790 3253.900 ;
        RECT 1852.030 3253.840 1852.350 3253.900 ;
        RECT 1393.870 3253.700 1394.190 3253.760 ;
        RECT 1441.710 3253.700 1442.030 3253.760 ;
        RECT 1393.870 3253.560 1442.030 3253.700 ;
        RECT 1393.870 3253.500 1394.190 3253.560 ;
        RECT 1441.710 3253.500 1442.030 3253.560 ;
        RECT 2863.110 3253.700 2863.430 3253.760 ;
        RECT 2897.610 3253.700 2897.930 3253.760 ;
        RECT 2863.110 3253.560 2897.930 3253.700 ;
        RECT 2863.110 3253.500 2863.430 3253.560 ;
        RECT 2897.610 3253.500 2897.930 3253.560 ;
        RECT 448.110 3253.020 448.430 3253.080 ;
        RECT 482.610 3253.020 482.930 3253.080 ;
        RECT 448.110 3252.880 482.930 3253.020 ;
        RECT 448.110 3252.820 448.430 3252.880 ;
        RECT 482.610 3252.820 482.930 3252.880 ;
        RECT 533.670 3253.020 533.990 3253.080 ;
        RECT 578.750 3253.020 579.070 3253.080 ;
        RECT 533.670 3252.880 579.070 3253.020 ;
        RECT 533.670 3252.820 533.990 3252.880 ;
        RECT 578.750 3252.820 579.070 3252.880 ;
        RECT 1703.910 3253.020 1704.230 3253.080 ;
        RECT 1738.410 3253.020 1738.730 3253.080 ;
        RECT 1703.910 3252.880 1738.730 3253.020 ;
        RECT 1703.910 3252.820 1704.230 3252.880 ;
        RECT 1738.410 3252.820 1738.730 3252.880 ;
        RECT 2801.470 3253.020 2801.790 3253.080 ;
        RECT 2815.730 3253.020 2816.050 3253.080 ;
        RECT 2801.470 3252.880 2816.050 3253.020 ;
        RECT 2801.470 3252.820 2801.790 3252.880 ;
        RECT 2815.730 3252.820 2816.050 3252.880 ;
        RECT 579.670 3252.680 579.990 3252.740 ;
        RECT 603.590 3252.680 603.910 3252.740 ;
        RECT 579.670 3252.540 603.910 3252.680 ;
        RECT 579.670 3252.480 579.990 3252.540 ;
        RECT 603.590 3252.480 603.910 3252.540 ;
        RECT 1449.070 3252.680 1449.390 3252.740 ;
        RECT 1463.330 3252.680 1463.650 3252.740 ;
        RECT 1449.070 3252.540 1463.650 3252.680 ;
        RECT 1449.070 3252.480 1449.390 3252.540 ;
        RECT 1463.330 3252.480 1463.650 3252.540 ;
        RECT 2028.670 3252.680 2028.990 3252.740 ;
        RECT 2066.850 3252.680 2067.170 3252.740 ;
        RECT 2028.670 3252.540 2067.170 3252.680 ;
        RECT 2028.670 3252.480 2028.990 3252.540 ;
        RECT 2066.850 3252.480 2067.170 3252.540 ;
        RECT 2669.910 3252.680 2670.230 3252.740 ;
        RECT 2704.410 3252.680 2704.730 3252.740 ;
        RECT 2669.910 3252.540 2704.730 3252.680 ;
        RECT 2669.910 3252.480 2670.230 3252.540 ;
        RECT 2704.410 3252.480 2704.730 3252.540 ;
        RECT 2283.510 3252.340 2283.830 3252.400 ;
        RECT 2318.010 3252.340 2318.330 3252.400 ;
        RECT 2283.510 3252.200 2318.330 3252.340 ;
        RECT 2283.510 3252.140 2283.830 3252.200 ;
        RECT 2318.010 3252.140 2318.330 3252.200 ;
        RECT 2380.110 3252.340 2380.430 3252.400 ;
        RECT 2414.610 3252.340 2414.930 3252.400 ;
        RECT 2380.110 3252.200 2414.930 3252.340 ;
        RECT 2380.110 3252.140 2380.430 3252.200 ;
        RECT 2414.610 3252.140 2414.930 3252.200 ;
        RECT 2476.710 3252.340 2477.030 3252.400 ;
        RECT 2511.210 3252.340 2511.530 3252.400 ;
        RECT 2476.710 3252.200 2511.530 3252.340 ;
        RECT 2476.710 3252.140 2477.030 3252.200 ;
        RECT 2511.210 3252.140 2511.530 3252.200 ;
        RECT 2573.310 3252.340 2573.630 3252.400 ;
        RECT 2607.810 3252.340 2608.130 3252.400 ;
        RECT 2573.310 3252.200 2608.130 3252.340 ;
        RECT 2573.310 3252.140 2573.630 3252.200 ;
        RECT 2607.810 3252.140 2608.130 3252.200 ;
      LAYER via ;
        RECT 1835.500 3253.840 1835.760 3254.100 ;
        RECT 1852.060 3253.840 1852.320 3254.100 ;
        RECT 1393.900 3253.500 1394.160 3253.760 ;
        RECT 1441.740 3253.500 1442.000 3253.760 ;
        RECT 2863.140 3253.500 2863.400 3253.760 ;
        RECT 2897.640 3253.500 2897.900 3253.760 ;
        RECT 448.140 3252.820 448.400 3253.080 ;
        RECT 482.640 3252.820 482.900 3253.080 ;
        RECT 533.700 3252.820 533.960 3253.080 ;
        RECT 578.780 3252.820 579.040 3253.080 ;
        RECT 1703.940 3252.820 1704.200 3253.080 ;
        RECT 1738.440 3252.820 1738.700 3253.080 ;
        RECT 2801.500 3252.820 2801.760 3253.080 ;
        RECT 2815.760 3252.820 2816.020 3253.080 ;
        RECT 579.700 3252.480 579.960 3252.740 ;
        RECT 603.620 3252.480 603.880 3252.740 ;
        RECT 1449.100 3252.480 1449.360 3252.740 ;
        RECT 1463.360 3252.480 1463.620 3252.740 ;
        RECT 2028.700 3252.480 2028.960 3252.740 ;
        RECT 2066.880 3252.480 2067.140 3252.740 ;
        RECT 2669.940 3252.480 2670.200 3252.740 ;
        RECT 2704.440 3252.480 2704.700 3252.740 ;
        RECT 2283.540 3252.140 2283.800 3252.400 ;
        RECT 2318.040 3252.140 2318.300 3252.400 ;
        RECT 2380.140 3252.140 2380.400 3252.400 ;
        RECT 2414.640 3252.140 2414.900 3252.400 ;
        RECT 2476.740 3252.140 2477.000 3252.400 ;
        RECT 2511.240 3252.140 2511.500 3252.400 ;
        RECT 2573.340 3252.140 2573.600 3252.400 ;
        RECT 2607.840 3252.140 2608.100 3252.400 ;
      LAYER met2 ;
        RECT 1931.630 3256.675 1931.910 3257.045 ;
        RECT 1852.050 3255.315 1852.330 3255.685 ;
        RECT 675.830 3254.635 676.110 3255.005 ;
        RECT 700.210 3254.890 700.490 3255.005 ;
        RECT 1559.950 3254.890 1560.230 3255.005 ;
        RECT 700.210 3254.750 700.880 3254.890 ;
        RECT 700.210 3254.635 700.490 3254.750 ;
        RECT 603.610 3253.955 603.890 3254.325 ;
        RECT 448.130 3253.275 448.410 3253.645 ;
        RECT 533.690 3253.275 533.970 3253.645 ;
        RECT 448.200 3253.110 448.340 3253.275 ;
        RECT 533.760 3253.110 533.900 3253.275 ;
        RECT 448.140 3252.790 448.400 3253.110 ;
        RECT 482.640 3252.965 482.900 3253.110 ;
        RECT 482.630 3252.595 482.910 3252.965 ;
        RECT 533.700 3252.790 533.960 3253.110 ;
        RECT 578.780 3252.965 579.040 3253.110 ;
        RECT 578.770 3252.595 579.050 3252.965 ;
        RECT 579.690 3252.595 579.970 3252.965 ;
        RECT 603.680 3252.770 603.820 3253.955 ;
        RECT 675.900 3252.965 676.040 3254.635 ;
        RECT 700.740 3253.645 700.880 3254.750 ;
        RECT 1559.100 3254.750 1560.230 3254.890 ;
        RECT 1559.100 3254.325 1559.240 3254.750 ;
        RECT 1559.950 3254.635 1560.230 3254.750 ;
        RECT 1545.230 3253.955 1545.510 3254.325 ;
        RECT 1559.030 3253.955 1559.310 3254.325 ;
        RECT 1835.490 3253.955 1835.770 3254.325 ;
        RECT 1852.120 3254.130 1852.260 3255.315 ;
        RECT 1931.700 3255.005 1931.840 3256.675 ;
        RECT 2004.310 3255.315 2004.590 3255.685 ;
        RECT 2916.950 3255.315 2917.230 3255.685 ;
        RECT 1931.630 3254.635 1931.910 3255.005 ;
        RECT 1945.890 3254.890 1946.170 3255.005 ;
        RECT 1945.890 3254.750 1946.560 3254.890 ;
        RECT 1945.890 3254.635 1946.170 3254.750 ;
        RECT 1946.420 3254.325 1946.560 3254.750 ;
        RECT 1393.900 3253.645 1394.160 3253.790 ;
        RECT 700.670 3253.275 700.950 3253.645 ;
        RECT 1393.890 3253.275 1394.170 3253.645 ;
        RECT 1441.740 3253.470 1442.000 3253.790 ;
        RECT 1441.800 3252.965 1441.940 3253.470 ;
        RECT 1463.350 3253.275 1463.630 3253.645 ;
        RECT 579.700 3252.450 579.960 3252.595 ;
        RECT 603.620 3252.450 603.880 3252.770 ;
        RECT 675.830 3252.595 676.110 3252.965 ;
        RECT 1441.730 3252.595 1442.010 3252.965 ;
        RECT 1449.090 3252.595 1449.370 3252.965 ;
        RECT 1463.420 3252.770 1463.560 3253.275 ;
        RECT 1449.100 3252.450 1449.360 3252.595 ;
        RECT 1463.360 3252.450 1463.620 3252.770 ;
        RECT 1545.300 3252.285 1545.440 3253.955 ;
        RECT 1835.500 3253.810 1835.760 3253.955 ;
        RECT 1852.060 3253.810 1852.320 3254.130 ;
        RECT 1946.350 3253.955 1946.630 3254.325 ;
        RECT 1703.930 3253.275 1704.210 3253.645 ;
        RECT 1704.000 3253.110 1704.140 3253.275 ;
        RECT 1607.330 3252.850 1607.610 3252.965 ;
        RECT 1608.250 3252.850 1608.530 3252.965 ;
        RECT 1607.330 3252.710 1608.530 3252.850 ;
        RECT 1703.940 3252.790 1704.200 3253.110 ;
        RECT 1738.440 3252.965 1738.700 3253.110 ;
        RECT 2004.380 3252.965 2004.520 3255.315 ;
        RECT 2917.020 3254.325 2917.160 3255.315 ;
        RECT 2221.430 3253.955 2221.710 3254.325 ;
        RECT 2815.750 3253.955 2816.030 3254.325 ;
        RECT 2916.950 3253.955 2917.230 3254.325 ;
        RECT 2221.500 3252.965 2221.640 3253.955 ;
        RECT 2815.820 3253.110 2815.960 3253.955 ;
        RECT 2863.140 3253.645 2863.400 3253.790 ;
        RECT 2897.640 3253.645 2897.900 3253.790 ;
        RECT 2863.130 3253.275 2863.410 3253.645 ;
        RECT 2897.630 3253.275 2897.910 3253.645 ;
        RECT 2801.500 3252.965 2801.760 3253.110 ;
        RECT 1607.330 3252.595 1607.610 3252.710 ;
        RECT 1608.250 3252.595 1608.530 3252.710 ;
        RECT 1738.430 3252.595 1738.710 3252.965 ;
        RECT 2004.310 3252.595 2004.590 3252.965 ;
        RECT 2028.690 3252.595 2028.970 3252.965 ;
        RECT 2091.250 3252.850 2091.530 3252.965 ;
        RECT 2028.700 3252.450 2028.960 3252.595 ;
        RECT 2066.880 3252.450 2067.140 3252.770 ;
        RECT 2090.400 3252.710 2091.530 3252.850 ;
        RECT 1545.230 3251.915 1545.510 3252.285 ;
        RECT 2066.940 3250.925 2067.080 3252.450 ;
        RECT 2090.400 3251.605 2090.540 3252.710 ;
        RECT 2091.250 3252.595 2091.530 3252.710 ;
        RECT 2221.430 3252.595 2221.710 3252.965 ;
        RECT 2318.030 3252.595 2318.310 3252.965 ;
        RECT 2414.630 3252.595 2414.910 3252.965 ;
        RECT 2511.230 3252.595 2511.510 3252.965 ;
        RECT 2607.830 3252.595 2608.110 3252.965 ;
        RECT 2318.100 3252.430 2318.240 3252.595 ;
        RECT 2414.700 3252.430 2414.840 3252.595 ;
        RECT 2511.300 3252.430 2511.440 3252.595 ;
        RECT 2607.900 3252.430 2608.040 3252.595 ;
        RECT 2669.940 3252.450 2670.200 3252.770 ;
        RECT 2704.430 3252.595 2704.710 3252.965 ;
        RECT 2801.490 3252.595 2801.770 3252.965 ;
        RECT 2815.760 3252.790 2816.020 3253.110 ;
        RECT 2704.440 3252.450 2704.700 3252.595 ;
        RECT 2283.540 3252.285 2283.800 3252.430 ;
        RECT 2283.530 3251.915 2283.810 3252.285 ;
        RECT 2318.040 3252.110 2318.300 3252.430 ;
        RECT 2380.140 3252.285 2380.400 3252.430 ;
        RECT 2380.130 3251.915 2380.410 3252.285 ;
        RECT 2414.640 3252.110 2414.900 3252.430 ;
        RECT 2476.740 3252.285 2477.000 3252.430 ;
        RECT 2476.730 3251.915 2477.010 3252.285 ;
        RECT 2511.240 3252.110 2511.500 3252.430 ;
        RECT 2573.340 3252.285 2573.600 3252.430 ;
        RECT 2573.330 3251.915 2573.610 3252.285 ;
        RECT 2607.840 3252.110 2608.100 3252.430 ;
        RECT 2670.000 3252.285 2670.140 3252.450 ;
        RECT 2669.930 3251.915 2670.210 3252.285 ;
        RECT 2090.330 3251.235 2090.610 3251.605 ;
        RECT 2066.870 3250.555 2067.150 3250.925 ;
      LAYER via2 ;
        RECT 1931.630 3256.720 1931.910 3257.000 ;
        RECT 1852.050 3255.360 1852.330 3255.640 ;
        RECT 675.830 3254.680 676.110 3254.960 ;
        RECT 700.210 3254.680 700.490 3254.960 ;
        RECT 603.610 3254.000 603.890 3254.280 ;
        RECT 448.130 3253.320 448.410 3253.600 ;
        RECT 533.690 3253.320 533.970 3253.600 ;
        RECT 482.630 3252.640 482.910 3252.920 ;
        RECT 578.770 3252.640 579.050 3252.920 ;
        RECT 579.690 3252.640 579.970 3252.920 ;
        RECT 1559.950 3254.680 1560.230 3254.960 ;
        RECT 1545.230 3254.000 1545.510 3254.280 ;
        RECT 1559.030 3254.000 1559.310 3254.280 ;
        RECT 1835.490 3254.000 1835.770 3254.280 ;
        RECT 2004.310 3255.360 2004.590 3255.640 ;
        RECT 2916.950 3255.360 2917.230 3255.640 ;
        RECT 1931.630 3254.680 1931.910 3254.960 ;
        RECT 1945.890 3254.680 1946.170 3254.960 ;
        RECT 700.670 3253.320 700.950 3253.600 ;
        RECT 1393.890 3253.320 1394.170 3253.600 ;
        RECT 1463.350 3253.320 1463.630 3253.600 ;
        RECT 675.830 3252.640 676.110 3252.920 ;
        RECT 1441.730 3252.640 1442.010 3252.920 ;
        RECT 1449.090 3252.640 1449.370 3252.920 ;
        RECT 1946.350 3254.000 1946.630 3254.280 ;
        RECT 1703.930 3253.320 1704.210 3253.600 ;
        RECT 1607.330 3252.640 1607.610 3252.920 ;
        RECT 1608.250 3252.640 1608.530 3252.920 ;
        RECT 2221.430 3254.000 2221.710 3254.280 ;
        RECT 2815.750 3254.000 2816.030 3254.280 ;
        RECT 2916.950 3254.000 2917.230 3254.280 ;
        RECT 2863.130 3253.320 2863.410 3253.600 ;
        RECT 2897.630 3253.320 2897.910 3253.600 ;
        RECT 1738.430 3252.640 1738.710 3252.920 ;
        RECT 2004.310 3252.640 2004.590 3252.920 ;
        RECT 2028.690 3252.640 2028.970 3252.920 ;
        RECT 1545.230 3251.960 1545.510 3252.240 ;
        RECT 2091.250 3252.640 2091.530 3252.920 ;
        RECT 2221.430 3252.640 2221.710 3252.920 ;
        RECT 2318.030 3252.640 2318.310 3252.920 ;
        RECT 2414.630 3252.640 2414.910 3252.920 ;
        RECT 2511.230 3252.640 2511.510 3252.920 ;
        RECT 2607.830 3252.640 2608.110 3252.920 ;
        RECT 2704.430 3252.640 2704.710 3252.920 ;
        RECT 2801.490 3252.640 2801.770 3252.920 ;
        RECT 2283.530 3251.960 2283.810 3252.240 ;
        RECT 2380.130 3251.960 2380.410 3252.240 ;
        RECT 2476.730 3251.960 2477.010 3252.240 ;
        RECT 2573.330 3251.960 2573.610 3252.240 ;
        RECT 2669.930 3251.960 2670.210 3252.240 ;
        RECT 2090.330 3251.280 2090.610 3251.560 ;
        RECT 2066.870 3250.600 2067.150 3250.880 ;
      LAYER met3 ;
        RECT 1883.510 3257.010 1883.890 3257.020 ;
        RECT 1931.605 3257.010 1931.935 3257.025 ;
        RECT 1883.510 3256.710 1931.935 3257.010 ;
        RECT 1883.510 3256.700 1883.890 3256.710 ;
        RECT 1931.605 3256.695 1931.935 3256.710 ;
        RECT 1852.025 3255.650 1852.355 3255.665 ;
        RECT 1883.510 3255.650 1883.890 3255.660 ;
        RECT 1852.025 3255.350 1883.890 3255.650 ;
        RECT 1852.025 3255.335 1852.355 3255.350 ;
        RECT 1883.510 3255.340 1883.890 3255.350 ;
        RECT 1980.110 3255.650 1980.490 3255.660 ;
        RECT 2004.285 3255.650 2004.615 3255.665 ;
        RECT 1980.110 3255.350 2004.615 3255.650 ;
        RECT 1980.110 3255.340 1980.490 3255.350 ;
        RECT 2004.285 3255.335 2004.615 3255.350 ;
        RECT 2916.925 3255.650 2917.255 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2916.925 3255.350 2924.800 3255.650 ;
        RECT 2916.925 3255.335 2917.255 3255.350 ;
        RECT 675.805 3254.970 676.135 3254.985 ;
        RECT 700.185 3254.970 700.515 3254.985 ;
        RECT 675.805 3254.670 700.515 3254.970 ;
        RECT 675.805 3254.655 676.135 3254.670 ;
        RECT 700.185 3254.655 700.515 3254.670 ;
        RECT 1559.925 3254.970 1560.255 3254.985 ;
        RECT 1593.710 3254.970 1594.090 3254.980 ;
        RECT 1559.925 3254.670 1594.090 3254.970 ;
        RECT 1559.925 3254.655 1560.255 3254.670 ;
        RECT 1593.710 3254.660 1594.090 3254.670 ;
        RECT 1931.605 3254.970 1931.935 3254.985 ;
        RECT 1945.865 3254.970 1946.195 3254.985 ;
        RECT 1931.605 3254.670 1946.195 3254.970 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 1931.605 3254.655 1931.935 3254.670 ;
        RECT 1945.865 3254.655 1946.195 3254.670 ;
        RECT 290.990 3254.290 291.370 3254.300 ;
        RECT 603.585 3254.290 603.915 3254.305 ;
        RECT 627.710 3254.290 628.090 3254.300 ;
        RECT 1545.205 3254.290 1545.535 3254.305 ;
        RECT 1559.005 3254.290 1559.335 3254.305 ;
        RECT 1835.465 3254.290 1835.795 3254.305 ;
        RECT 290.990 3253.990 352.050 3254.290 ;
        RECT 290.990 3253.980 291.370 3253.990 ;
        RECT 351.750 3252.930 352.050 3253.990 ;
        RECT 603.585 3253.990 628.090 3254.290 ;
        RECT 603.585 3253.975 603.915 3253.990 ;
        RECT 627.710 3253.980 628.090 3253.990 ;
        RECT 734.470 3253.990 835.050 3254.290 ;
        RECT 448.105 3253.610 448.435 3253.625 ;
        RECT 533.665 3253.610 533.995 3253.625 ;
        RECT 400.510 3253.310 448.435 3253.610 ;
        RECT 400.510 3252.930 400.810 3253.310 ;
        RECT 448.105 3253.295 448.435 3253.310 ;
        RECT 497.110 3253.310 533.995 3253.610 ;
        RECT 351.750 3252.630 400.810 3252.930 ;
        RECT 482.605 3252.930 482.935 3252.945 ;
        RECT 497.110 3252.930 497.410 3253.310 ;
        RECT 533.665 3253.295 533.995 3253.310 ;
        RECT 700.645 3253.610 700.975 3253.625 ;
        RECT 734.470 3253.610 734.770 3253.990 ;
        RECT 700.645 3253.310 734.770 3253.610 ;
        RECT 700.645 3253.295 700.975 3253.310 ;
        RECT 482.605 3252.630 497.410 3252.930 ;
        RECT 578.745 3252.930 579.075 3252.945 ;
        RECT 579.665 3252.930 579.995 3252.945 ;
        RECT 578.745 3252.630 579.995 3252.930 ;
        RECT 482.605 3252.615 482.935 3252.630 ;
        RECT 578.745 3252.615 579.075 3252.630 ;
        RECT 579.665 3252.615 579.995 3252.630 ;
        RECT 627.710 3252.930 628.090 3252.940 ;
        RECT 675.805 3252.930 676.135 3252.945 ;
        RECT 627.710 3252.630 676.135 3252.930 ;
        RECT 834.750 3252.930 835.050 3253.990 ;
        RECT 1545.205 3253.990 1559.335 3254.290 ;
        RECT 1545.205 3253.975 1545.535 3253.990 ;
        RECT 1559.005 3253.975 1559.335 3253.990 ;
        RECT 1800.750 3253.990 1835.795 3254.290 ;
        RECT 1393.865 3253.610 1394.195 3253.625 ;
        RECT 883.510 3253.310 930.730 3253.610 ;
        RECT 883.510 3252.930 883.810 3253.310 ;
        RECT 834.750 3252.630 883.810 3252.930 ;
        RECT 930.430 3252.930 930.730 3253.310 ;
        RECT 980.110 3253.310 1018.130 3253.610 ;
        RECT 980.110 3252.930 980.410 3253.310 ;
        RECT 930.430 3252.630 980.410 3252.930 ;
        RECT 1017.830 3252.930 1018.130 3253.310 ;
        RECT 1076.710 3253.310 1107.370 3253.610 ;
        RECT 1076.710 3252.930 1077.010 3253.310 ;
        RECT 1017.830 3252.630 1077.010 3252.930 ;
        RECT 1107.070 3252.930 1107.370 3253.310 ;
        RECT 1173.310 3253.310 1211.330 3253.610 ;
        RECT 1173.310 3252.930 1173.610 3253.310 ;
        RECT 1107.070 3252.630 1173.610 3252.930 ;
        RECT 1211.030 3252.930 1211.330 3253.310 ;
        RECT 1269.910 3253.310 1318.165 3253.610 ;
        RECT 1269.910 3252.930 1270.210 3253.310 ;
        RECT 1211.030 3252.630 1270.210 3252.930 ;
        RECT 1317.865 3252.930 1318.165 3253.310 ;
        RECT 1366.510 3253.310 1394.195 3253.610 ;
        RECT 1366.510 3252.930 1366.810 3253.310 ;
        RECT 1393.865 3253.295 1394.195 3253.310 ;
        RECT 1463.325 3253.610 1463.655 3253.625 ;
        RECT 1497.110 3253.610 1497.490 3253.620 ;
        RECT 1703.905 3253.610 1704.235 3253.625 ;
        RECT 1463.325 3253.310 1497.490 3253.610 ;
        RECT 1463.325 3253.295 1463.655 3253.310 ;
        RECT 1497.110 3253.300 1497.490 3253.310 ;
        RECT 1656.310 3253.310 1704.235 3253.610 ;
        RECT 1317.865 3252.630 1366.810 3252.930 ;
        RECT 1441.705 3252.930 1442.035 3252.945 ;
        RECT 1449.065 3252.930 1449.395 3252.945 ;
        RECT 1441.705 3252.630 1449.395 3252.930 ;
        RECT 627.710 3252.620 628.090 3252.630 ;
        RECT 675.805 3252.615 676.135 3252.630 ;
        RECT 1441.705 3252.615 1442.035 3252.630 ;
        RECT 1449.065 3252.615 1449.395 3252.630 ;
        RECT 1593.710 3252.930 1594.090 3252.940 ;
        RECT 1607.305 3252.930 1607.635 3252.945 ;
        RECT 1593.710 3252.630 1607.635 3252.930 ;
        RECT 1593.710 3252.620 1594.090 3252.630 ;
        RECT 1607.305 3252.615 1607.635 3252.630 ;
        RECT 1608.225 3252.930 1608.555 3252.945 ;
        RECT 1656.310 3252.930 1656.610 3253.310 ;
        RECT 1703.905 3253.295 1704.235 3253.310 ;
        RECT 1608.225 3252.630 1656.610 3252.930 ;
        RECT 1738.405 3252.930 1738.735 3252.945 ;
        RECT 1800.750 3252.930 1801.050 3253.990 ;
        RECT 1835.465 3253.975 1835.795 3253.990 ;
        RECT 1946.325 3254.290 1946.655 3254.305 ;
        RECT 1980.110 3254.290 1980.490 3254.300 ;
        RECT 1946.325 3253.990 1980.490 3254.290 ;
        RECT 1946.325 3253.975 1946.655 3253.990 ;
        RECT 1980.110 3253.980 1980.490 3253.990 ;
        RECT 2173.310 3254.290 2173.690 3254.300 ;
        RECT 2221.405 3254.290 2221.735 3254.305 ;
        RECT 2173.310 3253.990 2221.735 3254.290 ;
        RECT 2173.310 3253.980 2173.690 3253.990 ;
        RECT 2221.405 3253.975 2221.735 3253.990 ;
        RECT 2815.725 3254.290 2816.055 3254.305 ;
        RECT 2898.270 3254.290 2898.650 3254.300 ;
        RECT 2916.925 3254.290 2917.255 3254.305 ;
        RECT 2815.725 3253.990 2849.850 3254.290 ;
        RECT 2815.725 3253.975 2816.055 3253.990 ;
        RECT 2849.550 3253.610 2849.850 3253.990 ;
        RECT 2898.270 3253.990 2917.255 3254.290 ;
        RECT 2898.270 3253.980 2898.650 3253.990 ;
        RECT 2916.925 3253.975 2917.255 3253.990 ;
        RECT 2863.105 3253.610 2863.435 3253.625 ;
        RECT 2849.550 3253.310 2863.435 3253.610 ;
        RECT 2863.105 3253.295 2863.435 3253.310 ;
        RECT 2897.605 3253.610 2897.935 3253.625 ;
        RECT 2897.605 3253.310 2898.610 3253.610 ;
        RECT 2897.605 3253.295 2897.935 3253.310 ;
        RECT 1738.405 3252.630 1801.050 3252.930 ;
        RECT 2004.285 3252.930 2004.615 3252.945 ;
        RECT 2028.665 3252.930 2028.995 3252.945 ;
        RECT 2004.285 3252.630 2028.995 3252.930 ;
        RECT 1608.225 3252.615 1608.555 3252.630 ;
        RECT 1738.405 3252.615 1738.735 3252.630 ;
        RECT 2004.285 3252.615 2004.615 3252.630 ;
        RECT 2028.665 3252.615 2028.995 3252.630 ;
        RECT 2091.225 3252.930 2091.555 3252.945 ;
        RECT 2221.405 3252.930 2221.735 3252.945 ;
        RECT 2318.005 3252.930 2318.335 3252.945 ;
        RECT 2414.605 3252.930 2414.935 3252.945 ;
        RECT 2511.205 3252.930 2511.535 3252.945 ;
        RECT 2607.805 3252.930 2608.135 3252.945 ;
        RECT 2704.405 3252.930 2704.735 3252.945 ;
        RECT 2801.465 3252.930 2801.795 3252.945 ;
        RECT 2898.310 3252.940 2898.610 3253.310 ;
        RECT 2091.225 3252.630 2139.610 3252.930 ;
        RECT 2091.225 3252.615 2091.555 3252.630 ;
        RECT 1497.110 3252.250 1497.490 3252.260 ;
        RECT 1545.205 3252.250 1545.535 3252.265 ;
        RECT 1497.110 3251.950 1545.535 3252.250 ;
        RECT 2139.310 3252.250 2139.610 3252.630 ;
        RECT 2221.405 3252.630 2236.210 3252.930 ;
        RECT 2221.405 3252.615 2221.735 3252.630 ;
        RECT 2173.310 3252.250 2173.690 3252.260 ;
        RECT 2139.310 3251.950 2173.690 3252.250 ;
        RECT 2235.910 3252.250 2236.210 3252.630 ;
        RECT 2318.005 3252.630 2332.810 3252.930 ;
        RECT 2318.005 3252.615 2318.335 3252.630 ;
        RECT 2283.505 3252.250 2283.835 3252.265 ;
        RECT 2235.910 3251.950 2283.835 3252.250 ;
        RECT 2332.510 3252.250 2332.810 3252.630 ;
        RECT 2414.605 3252.630 2429.410 3252.930 ;
        RECT 2414.605 3252.615 2414.935 3252.630 ;
        RECT 2380.105 3252.250 2380.435 3252.265 ;
        RECT 2332.510 3251.950 2380.435 3252.250 ;
        RECT 2429.110 3252.250 2429.410 3252.630 ;
        RECT 2511.205 3252.630 2526.010 3252.930 ;
        RECT 2511.205 3252.615 2511.535 3252.630 ;
        RECT 2476.705 3252.250 2477.035 3252.265 ;
        RECT 2429.110 3251.950 2477.035 3252.250 ;
        RECT 2525.710 3252.250 2526.010 3252.630 ;
        RECT 2607.805 3252.630 2622.610 3252.930 ;
        RECT 2607.805 3252.615 2608.135 3252.630 ;
        RECT 2573.305 3252.250 2573.635 3252.265 ;
        RECT 2525.710 3251.950 2573.635 3252.250 ;
        RECT 2622.310 3252.250 2622.610 3252.630 ;
        RECT 2704.405 3252.630 2719.210 3252.930 ;
        RECT 2704.405 3252.615 2704.735 3252.630 ;
        RECT 2669.905 3252.250 2670.235 3252.265 ;
        RECT 2622.310 3251.950 2670.235 3252.250 ;
        RECT 2718.910 3252.250 2719.210 3252.630 ;
        RECT 2800.790 3252.630 2801.795 3252.930 ;
        RECT 2718.910 3251.950 2753.250 3252.250 ;
        RECT 1497.110 3251.940 1497.490 3251.950 ;
        RECT 1545.205 3251.935 1545.535 3251.950 ;
        RECT 2173.310 3251.940 2173.690 3251.950 ;
        RECT 2283.505 3251.935 2283.835 3251.950 ;
        RECT 2380.105 3251.935 2380.435 3251.950 ;
        RECT 2476.705 3251.935 2477.035 3251.950 ;
        RECT 2573.305 3251.935 2573.635 3251.950 ;
        RECT 2669.905 3251.935 2670.235 3251.950 ;
        RECT 2090.305 3251.570 2090.635 3251.585 ;
        RECT 2076.750 3251.270 2090.635 3251.570 ;
        RECT 2066.845 3250.890 2067.175 3250.905 ;
        RECT 2076.750 3250.890 2077.050 3251.270 ;
        RECT 2090.305 3251.255 2090.635 3251.270 ;
        RECT 2066.845 3250.590 2077.050 3250.890 ;
        RECT 2752.950 3250.890 2753.250 3251.950 ;
        RECT 2800.790 3250.890 2801.090 3252.630 ;
        RECT 2801.465 3252.615 2801.795 3252.630 ;
        RECT 2898.270 3252.620 2898.650 3252.940 ;
        RECT 2752.950 3250.590 2801.090 3250.890 ;
        RECT 2066.845 3250.575 2067.175 3250.590 ;
        RECT 290.990 1990.850 291.370 1990.860 ;
        RECT 300.000 1990.850 304.000 1990.960 ;
        RECT 290.990 1990.550 304.000 1990.850 ;
        RECT 290.990 1990.540 291.370 1990.550 ;
        RECT 300.000 1990.360 304.000 1990.550 ;
      LAYER via3 ;
        RECT 1883.540 3256.700 1883.860 3257.020 ;
        RECT 1883.540 3255.340 1883.860 3255.660 ;
        RECT 1980.140 3255.340 1980.460 3255.660 ;
        RECT 1593.740 3254.660 1594.060 3254.980 ;
        RECT 291.020 3253.980 291.340 3254.300 ;
        RECT 627.740 3253.980 628.060 3254.300 ;
        RECT 627.740 3252.620 628.060 3252.940 ;
        RECT 1497.140 3253.300 1497.460 3253.620 ;
        RECT 1593.740 3252.620 1594.060 3252.940 ;
        RECT 1980.140 3253.980 1980.460 3254.300 ;
        RECT 2173.340 3253.980 2173.660 3254.300 ;
        RECT 2898.300 3253.980 2898.620 3254.300 ;
        RECT 1497.140 3251.940 1497.460 3252.260 ;
        RECT 2173.340 3251.940 2173.660 3252.260 ;
        RECT 2898.300 3252.620 2898.620 3252.940 ;
        RECT 291.020 1990.540 291.340 1990.860 ;
      LAYER met4 ;
        RECT 1883.535 3256.695 1883.865 3257.025 ;
        RECT 1883.550 3255.665 1883.850 3256.695 ;
        RECT 1883.535 3255.335 1883.865 3255.665 ;
        RECT 1980.135 3255.335 1980.465 3255.665 ;
        RECT 1593.735 3254.655 1594.065 3254.985 ;
        RECT 291.015 3253.975 291.345 3254.305 ;
        RECT 627.735 3253.975 628.065 3254.305 ;
        RECT 291.030 1990.865 291.330 3253.975 ;
        RECT 627.750 3252.945 628.050 3253.975 ;
        RECT 1497.135 3253.295 1497.465 3253.625 ;
        RECT 627.735 3252.615 628.065 3252.945 ;
        RECT 1497.150 3252.265 1497.450 3253.295 ;
        RECT 1593.750 3252.945 1594.050 3254.655 ;
        RECT 1980.150 3254.305 1980.450 3255.335 ;
        RECT 1980.135 3253.975 1980.465 3254.305 ;
        RECT 2173.335 3253.975 2173.665 3254.305 ;
        RECT 2898.295 3253.975 2898.625 3254.305 ;
        RECT 1593.735 3252.615 1594.065 3252.945 ;
        RECT 2173.350 3252.265 2173.650 3253.975 ;
        RECT 2898.310 3252.945 2898.610 3253.975 ;
        RECT 2898.295 3252.615 2898.625 3252.945 ;
        RECT 1497.135 3251.935 1497.465 3252.265 ;
        RECT 2173.335 3251.935 2173.665 3252.265 ;
        RECT 291.015 1990.535 291.345 1990.865 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2801.470 3486.600 2801.790 3486.660 ;
        RECT 2825.850 3486.600 2826.170 3486.660 ;
        RECT 2801.470 3486.460 2826.170 3486.600 ;
        RECT 2801.470 3486.400 2801.790 3486.460 ;
        RECT 2825.850 3486.400 2826.170 3486.460 ;
        RECT 2704.870 3485.920 2705.190 3485.980 ;
        RECT 2743.050 3485.920 2743.370 3485.980 ;
        RECT 2704.870 3485.780 2743.370 3485.920 ;
        RECT 2704.870 3485.720 2705.190 3485.780 ;
        RECT 2743.050 3485.720 2743.370 3485.780 ;
        RECT 351.510 3485.580 351.830 3485.640 ;
        RECT 386.010 3485.580 386.330 3485.640 ;
        RECT 351.510 3485.440 386.330 3485.580 ;
        RECT 351.510 3485.380 351.830 3485.440 ;
        RECT 386.010 3485.380 386.330 3485.440 ;
        RECT 448.110 3485.580 448.430 3485.640 ;
        RECT 482.610 3485.580 482.930 3485.640 ;
        RECT 448.110 3485.440 482.930 3485.580 ;
        RECT 448.110 3485.380 448.430 3485.440 ;
        RECT 482.610 3485.380 482.930 3485.440 ;
        RECT 544.710 3485.580 545.030 3485.640 ;
        RECT 579.210 3485.580 579.530 3485.640 ;
        RECT 544.710 3485.440 579.530 3485.580 ;
        RECT 544.710 3485.380 545.030 3485.440 ;
        RECT 579.210 3485.380 579.530 3485.440 ;
        RECT 641.310 3485.580 641.630 3485.640 ;
        RECT 675.810 3485.580 676.130 3485.640 ;
        RECT 641.310 3485.440 676.130 3485.580 ;
        RECT 641.310 3485.380 641.630 3485.440 ;
        RECT 675.810 3485.380 676.130 3485.440 ;
        RECT 737.910 3485.580 738.230 3485.640 ;
        RECT 772.410 3485.580 772.730 3485.640 ;
        RECT 737.910 3485.440 772.730 3485.580 ;
        RECT 737.910 3485.380 738.230 3485.440 ;
        RECT 772.410 3485.380 772.730 3485.440 ;
        RECT 834.510 3485.580 834.830 3485.640 ;
        RECT 869.010 3485.580 869.330 3485.640 ;
        RECT 834.510 3485.440 869.330 3485.580 ;
        RECT 834.510 3485.380 834.830 3485.440 ;
        RECT 869.010 3485.380 869.330 3485.440 ;
        RECT 931.110 3485.580 931.430 3485.640 ;
        RECT 965.610 3485.580 965.930 3485.640 ;
        RECT 931.110 3485.440 965.930 3485.580 ;
        RECT 931.110 3485.380 931.430 3485.440 ;
        RECT 965.610 3485.380 965.930 3485.440 ;
        RECT 1027.710 3485.580 1028.030 3485.640 ;
        RECT 1062.210 3485.580 1062.530 3485.640 ;
        RECT 1027.710 3485.440 1062.530 3485.580 ;
        RECT 1027.710 3485.380 1028.030 3485.440 ;
        RECT 1062.210 3485.380 1062.530 3485.440 ;
        RECT 1124.310 3485.580 1124.630 3485.640 ;
        RECT 1158.810 3485.580 1159.130 3485.640 ;
        RECT 1124.310 3485.440 1159.130 3485.580 ;
        RECT 1124.310 3485.380 1124.630 3485.440 ;
        RECT 1158.810 3485.380 1159.130 3485.440 ;
        RECT 1220.910 3485.580 1221.230 3485.640 ;
        RECT 1255.410 3485.580 1255.730 3485.640 ;
        RECT 1220.910 3485.440 1255.730 3485.580 ;
        RECT 1220.910 3485.380 1221.230 3485.440 ;
        RECT 1255.410 3485.380 1255.730 3485.440 ;
        RECT 1317.510 3485.580 1317.830 3485.640 ;
        RECT 1352.010 3485.580 1352.330 3485.640 ;
        RECT 1317.510 3485.440 1352.330 3485.580 ;
        RECT 1317.510 3485.380 1317.830 3485.440 ;
        RECT 1352.010 3485.380 1352.330 3485.440 ;
        RECT 1414.110 3485.580 1414.430 3485.640 ;
        RECT 1448.610 3485.580 1448.930 3485.640 ;
        RECT 1414.110 3485.440 1448.930 3485.580 ;
        RECT 1414.110 3485.380 1414.430 3485.440 ;
        RECT 1448.610 3485.380 1448.930 3485.440 ;
        RECT 1510.710 3485.580 1511.030 3485.640 ;
        RECT 1545.210 3485.580 1545.530 3485.640 ;
        RECT 1510.710 3485.440 1545.530 3485.580 ;
        RECT 1510.710 3485.380 1511.030 3485.440 ;
        RECT 1545.210 3485.380 1545.530 3485.440 ;
        RECT 1607.310 3485.580 1607.630 3485.640 ;
        RECT 1641.810 3485.580 1642.130 3485.640 ;
        RECT 1607.310 3485.440 1642.130 3485.580 ;
        RECT 1607.310 3485.380 1607.630 3485.440 ;
        RECT 1641.810 3485.380 1642.130 3485.440 ;
      LAYER via ;
        RECT 2801.500 3486.400 2801.760 3486.660 ;
        RECT 2825.880 3486.400 2826.140 3486.660 ;
        RECT 2704.900 3485.720 2705.160 3485.980 ;
        RECT 2743.080 3485.720 2743.340 3485.980 ;
        RECT 351.540 3485.380 351.800 3485.640 ;
        RECT 386.040 3485.380 386.300 3485.640 ;
        RECT 448.140 3485.380 448.400 3485.640 ;
        RECT 482.640 3485.380 482.900 3485.640 ;
        RECT 544.740 3485.380 545.000 3485.640 ;
        RECT 579.240 3485.380 579.500 3485.640 ;
        RECT 641.340 3485.380 641.600 3485.640 ;
        RECT 675.840 3485.380 676.100 3485.640 ;
        RECT 737.940 3485.380 738.200 3485.640 ;
        RECT 772.440 3485.380 772.700 3485.640 ;
        RECT 834.540 3485.380 834.800 3485.640 ;
        RECT 869.040 3485.380 869.300 3485.640 ;
        RECT 931.140 3485.380 931.400 3485.640 ;
        RECT 965.640 3485.380 965.900 3485.640 ;
        RECT 1027.740 3485.380 1028.000 3485.640 ;
        RECT 1062.240 3485.380 1062.500 3485.640 ;
        RECT 1124.340 3485.380 1124.600 3485.640 ;
        RECT 1158.840 3485.380 1159.100 3485.640 ;
        RECT 1220.940 3485.380 1221.200 3485.640 ;
        RECT 1255.440 3485.380 1255.700 3485.640 ;
        RECT 1317.540 3485.380 1317.800 3485.640 ;
        RECT 1352.040 3485.380 1352.300 3485.640 ;
        RECT 1414.140 3485.380 1414.400 3485.640 ;
        RECT 1448.640 3485.380 1448.900 3485.640 ;
        RECT 1510.740 3485.380 1511.000 3485.640 ;
        RECT 1545.240 3485.380 1545.500 3485.640 ;
        RECT 1607.340 3485.380 1607.600 3485.640 ;
        RECT 1641.840 3485.380 1642.100 3485.640 ;
      LAYER met2 ;
        RECT 2766.530 3486.770 2766.810 3486.885 ;
        RECT 2767.450 3486.770 2767.730 3486.885 ;
        RECT 2766.530 3486.630 2767.730 3486.770 ;
        RECT 2766.530 3486.515 2766.810 3486.630 ;
        RECT 2767.450 3486.515 2767.730 3486.630 ;
        RECT 2801.490 3486.515 2801.770 3486.885 ;
        RECT 2801.500 3486.370 2801.760 3486.515 ;
        RECT 2825.880 3486.370 2826.140 3486.690 ;
        RECT 2825.940 3486.205 2826.080 3486.370 ;
        RECT 386.030 3485.835 386.310 3486.205 ;
        RECT 482.630 3485.835 482.910 3486.205 ;
        RECT 579.230 3485.835 579.510 3486.205 ;
        RECT 675.830 3485.835 676.110 3486.205 ;
        RECT 772.430 3485.835 772.710 3486.205 ;
        RECT 869.030 3485.835 869.310 3486.205 ;
        RECT 965.630 3485.835 965.910 3486.205 ;
        RECT 1062.230 3485.835 1062.510 3486.205 ;
        RECT 1158.830 3485.835 1159.110 3486.205 ;
        RECT 1255.430 3485.835 1255.710 3486.205 ;
        RECT 1352.030 3485.835 1352.310 3486.205 ;
        RECT 1448.630 3485.835 1448.910 3486.205 ;
        RECT 1545.230 3485.835 1545.510 3486.205 ;
        RECT 1641.830 3485.835 1642.110 3486.205 ;
        RECT 2704.890 3485.835 2705.170 3486.205 ;
        RECT 386.100 3485.670 386.240 3485.835 ;
        RECT 482.700 3485.670 482.840 3485.835 ;
        RECT 579.300 3485.670 579.440 3485.835 ;
        RECT 675.900 3485.670 676.040 3485.835 ;
        RECT 772.500 3485.670 772.640 3485.835 ;
        RECT 869.100 3485.670 869.240 3485.835 ;
        RECT 965.700 3485.670 965.840 3485.835 ;
        RECT 1062.300 3485.670 1062.440 3485.835 ;
        RECT 1158.900 3485.670 1159.040 3485.835 ;
        RECT 1255.500 3485.670 1255.640 3485.835 ;
        RECT 1352.100 3485.670 1352.240 3485.835 ;
        RECT 1448.700 3485.670 1448.840 3485.835 ;
        RECT 1545.300 3485.670 1545.440 3485.835 ;
        RECT 1641.900 3485.670 1642.040 3485.835 ;
        RECT 2704.900 3485.690 2705.160 3485.835 ;
        RECT 2743.080 3485.690 2743.340 3486.010 ;
        RECT 2825.870 3485.835 2826.150 3486.205 ;
        RECT 2863.590 3486.090 2863.870 3486.205 ;
        RECT 2863.200 3485.950 2863.870 3486.090 ;
        RECT 351.540 3485.525 351.800 3485.670 ;
        RECT 351.530 3485.155 351.810 3485.525 ;
        RECT 386.040 3485.350 386.300 3485.670 ;
        RECT 448.140 3485.525 448.400 3485.670 ;
        RECT 448.130 3485.155 448.410 3485.525 ;
        RECT 482.640 3485.350 482.900 3485.670 ;
        RECT 544.740 3485.525 545.000 3485.670 ;
        RECT 544.730 3485.155 545.010 3485.525 ;
        RECT 579.240 3485.350 579.500 3485.670 ;
        RECT 641.340 3485.525 641.600 3485.670 ;
        RECT 641.330 3485.155 641.610 3485.525 ;
        RECT 675.840 3485.350 676.100 3485.670 ;
        RECT 737.940 3485.525 738.200 3485.670 ;
        RECT 737.930 3485.155 738.210 3485.525 ;
        RECT 772.440 3485.350 772.700 3485.670 ;
        RECT 834.540 3485.525 834.800 3485.670 ;
        RECT 834.530 3485.155 834.810 3485.525 ;
        RECT 869.040 3485.350 869.300 3485.670 ;
        RECT 931.140 3485.525 931.400 3485.670 ;
        RECT 931.130 3485.155 931.410 3485.525 ;
        RECT 965.640 3485.350 965.900 3485.670 ;
        RECT 1027.740 3485.525 1028.000 3485.670 ;
        RECT 1027.730 3485.155 1028.010 3485.525 ;
        RECT 1062.240 3485.350 1062.500 3485.670 ;
        RECT 1124.340 3485.525 1124.600 3485.670 ;
        RECT 1124.330 3485.155 1124.610 3485.525 ;
        RECT 1158.840 3485.350 1159.100 3485.670 ;
        RECT 1220.940 3485.525 1221.200 3485.670 ;
        RECT 1220.930 3485.155 1221.210 3485.525 ;
        RECT 1255.440 3485.350 1255.700 3485.670 ;
        RECT 1317.540 3485.525 1317.800 3485.670 ;
        RECT 1317.530 3485.155 1317.810 3485.525 ;
        RECT 1352.040 3485.350 1352.300 3485.670 ;
        RECT 1414.140 3485.525 1414.400 3485.670 ;
        RECT 1414.130 3485.155 1414.410 3485.525 ;
        RECT 1448.640 3485.350 1448.900 3485.670 ;
        RECT 1510.740 3485.525 1511.000 3485.670 ;
        RECT 1510.730 3485.155 1511.010 3485.525 ;
        RECT 1545.240 3485.350 1545.500 3485.670 ;
        RECT 1607.340 3485.525 1607.600 3485.670 ;
        RECT 1607.330 3485.155 1607.610 3485.525 ;
        RECT 1641.840 3485.350 1642.100 3485.670 ;
        RECT 2743.140 3484.845 2743.280 3485.690 ;
        RECT 2863.200 3485.525 2863.340 3485.950 ;
        RECT 2863.590 3485.835 2863.870 3485.950 ;
        RECT 2863.130 3485.155 2863.410 3485.525 ;
        RECT 2743.070 3484.475 2743.350 3484.845 ;
      LAYER via2 ;
        RECT 2766.530 3486.560 2766.810 3486.840 ;
        RECT 2767.450 3486.560 2767.730 3486.840 ;
        RECT 2801.490 3486.560 2801.770 3486.840 ;
        RECT 386.030 3485.880 386.310 3486.160 ;
        RECT 482.630 3485.880 482.910 3486.160 ;
        RECT 579.230 3485.880 579.510 3486.160 ;
        RECT 675.830 3485.880 676.110 3486.160 ;
        RECT 772.430 3485.880 772.710 3486.160 ;
        RECT 869.030 3485.880 869.310 3486.160 ;
        RECT 965.630 3485.880 965.910 3486.160 ;
        RECT 1062.230 3485.880 1062.510 3486.160 ;
        RECT 1158.830 3485.880 1159.110 3486.160 ;
        RECT 1255.430 3485.880 1255.710 3486.160 ;
        RECT 1352.030 3485.880 1352.310 3486.160 ;
        RECT 1448.630 3485.880 1448.910 3486.160 ;
        RECT 1545.230 3485.880 1545.510 3486.160 ;
        RECT 1641.830 3485.880 1642.110 3486.160 ;
        RECT 2704.890 3485.880 2705.170 3486.160 ;
        RECT 2825.870 3485.880 2826.150 3486.160 ;
        RECT 351.530 3485.200 351.810 3485.480 ;
        RECT 448.130 3485.200 448.410 3485.480 ;
        RECT 544.730 3485.200 545.010 3485.480 ;
        RECT 641.330 3485.200 641.610 3485.480 ;
        RECT 737.930 3485.200 738.210 3485.480 ;
        RECT 834.530 3485.200 834.810 3485.480 ;
        RECT 931.130 3485.200 931.410 3485.480 ;
        RECT 1027.730 3485.200 1028.010 3485.480 ;
        RECT 1124.330 3485.200 1124.610 3485.480 ;
        RECT 1220.930 3485.200 1221.210 3485.480 ;
        RECT 1317.530 3485.200 1317.810 3485.480 ;
        RECT 1414.130 3485.200 1414.410 3485.480 ;
        RECT 1510.730 3485.200 1511.010 3485.480 ;
        RECT 1607.330 3485.200 1607.610 3485.480 ;
        RECT 2863.590 3485.880 2863.870 3486.160 ;
        RECT 2863.130 3485.200 2863.410 3485.480 ;
        RECT 2743.070 3484.520 2743.350 3484.800 ;
      LAYER met3 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2916.710 3489.950 2924.800 3490.250 ;
        RECT 2752.910 3486.850 2753.290 3486.860 ;
        RECT 2766.505 3486.850 2766.835 3486.865 ;
        RECT 2752.910 3486.550 2766.835 3486.850 ;
        RECT 2752.910 3486.540 2753.290 3486.550 ;
        RECT 2766.505 3486.535 2766.835 3486.550 ;
        RECT 2767.425 3486.850 2767.755 3486.865 ;
        RECT 2801.465 3486.850 2801.795 3486.865 ;
        RECT 2767.425 3486.550 2801.795 3486.850 ;
        RECT 2767.425 3486.535 2767.755 3486.550 ;
        RECT 2801.465 3486.535 2801.795 3486.550 ;
        RECT 295.590 3486.170 295.970 3486.180 ;
        RECT 386.005 3486.170 386.335 3486.185 ;
        RECT 482.605 3486.170 482.935 3486.185 ;
        RECT 579.205 3486.170 579.535 3486.185 ;
        RECT 675.805 3486.170 676.135 3486.185 ;
        RECT 772.405 3486.170 772.735 3486.185 ;
        RECT 869.005 3486.170 869.335 3486.185 ;
        RECT 965.605 3486.170 965.935 3486.185 ;
        RECT 1062.205 3486.170 1062.535 3486.185 ;
        RECT 1158.805 3486.170 1159.135 3486.185 ;
        RECT 1255.405 3486.170 1255.735 3486.185 ;
        RECT 1352.005 3486.170 1352.335 3486.185 ;
        RECT 1448.605 3486.170 1448.935 3486.185 ;
        RECT 1545.205 3486.170 1545.535 3486.185 ;
        RECT 1641.805 3486.170 1642.135 3486.185 ;
        RECT 2704.865 3486.170 2705.195 3486.185 ;
        RECT 295.590 3485.870 304.210 3486.170 ;
        RECT 295.590 3485.860 295.970 3485.870 ;
        RECT 303.910 3485.490 304.210 3485.870 ;
        RECT 386.005 3485.870 400.810 3486.170 ;
        RECT 386.005 3485.855 386.335 3485.870 ;
        RECT 351.505 3485.490 351.835 3485.505 ;
        RECT 303.910 3485.190 351.835 3485.490 ;
        RECT 400.510 3485.490 400.810 3485.870 ;
        RECT 482.605 3485.870 497.410 3486.170 ;
        RECT 482.605 3485.855 482.935 3485.870 ;
        RECT 448.105 3485.490 448.435 3485.505 ;
        RECT 400.510 3485.190 448.435 3485.490 ;
        RECT 497.110 3485.490 497.410 3485.870 ;
        RECT 579.205 3485.870 594.010 3486.170 ;
        RECT 579.205 3485.855 579.535 3485.870 ;
        RECT 544.705 3485.490 545.035 3485.505 ;
        RECT 497.110 3485.190 545.035 3485.490 ;
        RECT 593.710 3485.490 594.010 3485.870 ;
        RECT 675.805 3485.870 690.610 3486.170 ;
        RECT 675.805 3485.855 676.135 3485.870 ;
        RECT 641.305 3485.490 641.635 3485.505 ;
        RECT 593.710 3485.190 641.635 3485.490 ;
        RECT 690.310 3485.490 690.610 3485.870 ;
        RECT 772.405 3485.870 787.210 3486.170 ;
        RECT 772.405 3485.855 772.735 3485.870 ;
        RECT 737.905 3485.490 738.235 3485.505 ;
        RECT 690.310 3485.190 738.235 3485.490 ;
        RECT 786.910 3485.490 787.210 3485.870 ;
        RECT 869.005 3485.870 883.810 3486.170 ;
        RECT 869.005 3485.855 869.335 3485.870 ;
        RECT 834.505 3485.490 834.835 3485.505 ;
        RECT 786.910 3485.190 834.835 3485.490 ;
        RECT 883.510 3485.490 883.810 3485.870 ;
        RECT 965.605 3485.870 980.410 3486.170 ;
        RECT 965.605 3485.855 965.935 3485.870 ;
        RECT 931.105 3485.490 931.435 3485.505 ;
        RECT 883.510 3485.190 931.435 3485.490 ;
        RECT 980.110 3485.490 980.410 3485.870 ;
        RECT 1062.205 3485.870 1077.010 3486.170 ;
        RECT 1062.205 3485.855 1062.535 3485.870 ;
        RECT 1027.705 3485.490 1028.035 3485.505 ;
        RECT 980.110 3485.190 1028.035 3485.490 ;
        RECT 1076.710 3485.490 1077.010 3485.870 ;
        RECT 1158.805 3485.870 1173.610 3486.170 ;
        RECT 1158.805 3485.855 1159.135 3485.870 ;
        RECT 1124.305 3485.490 1124.635 3485.505 ;
        RECT 1076.710 3485.190 1124.635 3485.490 ;
        RECT 1173.310 3485.490 1173.610 3485.870 ;
        RECT 1255.405 3485.870 1270.210 3486.170 ;
        RECT 1255.405 3485.855 1255.735 3485.870 ;
        RECT 1220.905 3485.490 1221.235 3485.505 ;
        RECT 1173.310 3485.190 1221.235 3485.490 ;
        RECT 1269.910 3485.490 1270.210 3485.870 ;
        RECT 1352.005 3485.870 1366.810 3486.170 ;
        RECT 1352.005 3485.855 1352.335 3485.870 ;
        RECT 1317.505 3485.490 1317.835 3485.505 ;
        RECT 1269.910 3485.190 1317.835 3485.490 ;
        RECT 1366.510 3485.490 1366.810 3485.870 ;
        RECT 1448.605 3485.870 1463.410 3486.170 ;
        RECT 1448.605 3485.855 1448.935 3485.870 ;
        RECT 1414.105 3485.490 1414.435 3485.505 ;
        RECT 1366.510 3485.190 1414.435 3485.490 ;
        RECT 1463.110 3485.490 1463.410 3485.870 ;
        RECT 1545.205 3485.870 1560.010 3486.170 ;
        RECT 1545.205 3485.855 1545.535 3485.870 ;
        RECT 1510.705 3485.490 1511.035 3485.505 ;
        RECT 1463.110 3485.190 1511.035 3485.490 ;
        RECT 1559.710 3485.490 1560.010 3485.870 ;
        RECT 1641.805 3485.870 1704.450 3486.170 ;
        RECT 1641.805 3485.855 1642.135 3485.870 ;
        RECT 1607.305 3485.490 1607.635 3485.505 ;
        RECT 1559.710 3485.190 1607.635 3485.490 ;
        RECT 1704.150 3485.490 1704.450 3485.870 ;
        RECT 1869.750 3485.870 1917.890 3486.170 ;
        RECT 1704.150 3485.190 1752.290 3485.490 ;
        RECT 351.505 3485.175 351.835 3485.190 ;
        RECT 448.105 3485.175 448.435 3485.190 ;
        RECT 544.705 3485.175 545.035 3485.190 ;
        RECT 641.305 3485.175 641.635 3485.190 ;
        RECT 737.905 3485.175 738.235 3485.190 ;
        RECT 834.505 3485.175 834.835 3485.190 ;
        RECT 931.105 3485.175 931.435 3485.190 ;
        RECT 1027.705 3485.175 1028.035 3485.190 ;
        RECT 1124.305 3485.175 1124.635 3485.190 ;
        RECT 1220.905 3485.175 1221.235 3485.190 ;
        RECT 1317.505 3485.175 1317.835 3485.190 ;
        RECT 1414.105 3485.175 1414.435 3485.190 ;
        RECT 1510.705 3485.175 1511.035 3485.190 ;
        RECT 1607.305 3485.175 1607.635 3485.190 ;
        RECT 1751.990 3484.810 1752.290 3485.190 ;
        RECT 1869.750 3484.810 1870.050 3485.870 ;
        RECT 1751.990 3484.510 1870.050 3484.810 ;
        RECT 1917.590 3484.810 1917.890 3485.870 ;
        RECT 1918.510 3485.870 1966.650 3486.170 ;
        RECT 1918.510 3484.810 1918.810 3485.870 ;
        RECT 1966.350 3485.490 1966.650 3485.870 ;
        RECT 2015.110 3485.870 2063.250 3486.170 ;
        RECT 1966.350 3485.190 2014.490 3485.490 ;
        RECT 1917.590 3484.510 1918.810 3484.810 ;
        RECT 2014.190 3484.810 2014.490 3485.190 ;
        RECT 2015.110 3484.810 2015.410 3485.870 ;
        RECT 2062.950 3485.490 2063.250 3485.870 ;
        RECT 2111.710 3485.870 2159.850 3486.170 ;
        RECT 2062.950 3485.190 2111.090 3485.490 ;
        RECT 2014.190 3484.510 2015.410 3484.810 ;
        RECT 2110.790 3484.810 2111.090 3485.190 ;
        RECT 2111.710 3484.810 2112.010 3485.870 ;
        RECT 2159.550 3485.490 2159.850 3485.870 ;
        RECT 2208.310 3485.870 2256.450 3486.170 ;
        RECT 2159.550 3485.190 2207.690 3485.490 ;
        RECT 2110.790 3484.510 2112.010 3484.810 ;
        RECT 2207.390 3484.810 2207.690 3485.190 ;
        RECT 2208.310 3484.810 2208.610 3485.870 ;
        RECT 2256.150 3485.490 2256.450 3485.870 ;
        RECT 2304.910 3485.870 2353.050 3486.170 ;
        RECT 2256.150 3485.190 2304.290 3485.490 ;
        RECT 2207.390 3484.510 2208.610 3484.810 ;
        RECT 2303.990 3484.810 2304.290 3485.190 ;
        RECT 2304.910 3484.810 2305.210 3485.870 ;
        RECT 2352.750 3485.490 2353.050 3485.870 ;
        RECT 2401.510 3485.870 2449.650 3486.170 ;
        RECT 2352.750 3485.190 2400.890 3485.490 ;
        RECT 2303.990 3484.510 2305.210 3484.810 ;
        RECT 2400.590 3484.810 2400.890 3485.190 ;
        RECT 2401.510 3484.810 2401.810 3485.870 ;
        RECT 2449.350 3485.490 2449.650 3485.870 ;
        RECT 2498.110 3485.870 2546.250 3486.170 ;
        RECT 2449.350 3485.190 2497.490 3485.490 ;
        RECT 2400.590 3484.510 2401.810 3484.810 ;
        RECT 2497.190 3484.810 2497.490 3485.190 ;
        RECT 2498.110 3484.810 2498.410 3485.870 ;
        RECT 2545.950 3485.490 2546.250 3485.870 ;
        RECT 2594.710 3485.870 2642.850 3486.170 ;
        RECT 2545.950 3485.190 2594.090 3485.490 ;
        RECT 2497.190 3484.510 2498.410 3484.810 ;
        RECT 2593.790 3484.810 2594.090 3485.190 ;
        RECT 2594.710 3484.810 2595.010 3485.870 ;
        RECT 2642.550 3485.490 2642.850 3485.870 ;
        RECT 2691.310 3485.870 2705.195 3486.170 ;
        RECT 2642.550 3485.190 2690.690 3485.490 ;
        RECT 2593.790 3484.510 2595.010 3484.810 ;
        RECT 2690.390 3484.810 2690.690 3485.190 ;
        RECT 2691.310 3484.810 2691.610 3485.870 ;
        RECT 2704.865 3485.855 2705.195 3485.870 ;
        RECT 2825.845 3486.170 2826.175 3486.185 ;
        RECT 2863.565 3486.170 2863.895 3486.185 ;
        RECT 2825.845 3485.870 2849.850 3486.170 ;
        RECT 2825.845 3485.855 2826.175 3485.870 ;
        RECT 2849.550 3485.490 2849.850 3485.870 ;
        RECT 2863.565 3485.870 2884.810 3486.170 ;
        RECT 2863.565 3485.855 2863.895 3485.870 ;
        RECT 2863.105 3485.490 2863.435 3485.505 ;
        RECT 2849.550 3485.190 2863.435 3485.490 ;
        RECT 2884.510 3485.490 2884.810 3485.870 ;
        RECT 2916.710 3485.490 2917.010 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2884.510 3485.190 2917.010 3485.490 ;
        RECT 2863.105 3485.175 2863.435 3485.190 ;
        RECT 2690.390 3484.510 2691.610 3484.810 ;
        RECT 2743.045 3484.810 2743.375 3484.825 ;
        RECT 2752.910 3484.810 2753.290 3484.820 ;
        RECT 2743.045 3484.510 2753.290 3484.810 ;
        RECT 2743.045 3484.495 2743.375 3484.510 ;
        RECT 2752.910 3484.500 2753.290 3484.510 ;
        RECT 295.590 2020.090 295.970 2020.100 ;
        RECT 300.000 2020.090 304.000 2020.200 ;
        RECT 295.590 2019.790 304.000 2020.090 ;
        RECT 295.590 2019.780 295.970 2019.790 ;
        RECT 300.000 2019.600 304.000 2019.790 ;
      LAYER via3 ;
        RECT 2752.940 3486.540 2753.260 3486.860 ;
        RECT 295.620 3485.860 295.940 3486.180 ;
        RECT 2752.940 3484.500 2753.260 3484.820 ;
        RECT 295.620 2019.780 295.940 2020.100 ;
      LAYER met4 ;
        RECT 2752.935 3486.535 2753.265 3486.865 ;
        RECT 295.615 3485.855 295.945 3486.185 ;
        RECT 295.630 2020.105 295.930 3485.855 ;
        RECT 2752.950 3484.825 2753.250 3486.535 ;
        RECT 2752.935 3484.495 2753.265 3484.825 ;
        RECT 295.615 2019.775 295.945 2020.105 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 296.770 3501.560 297.090 3501.620 ;
        RECT 2635.870 3501.560 2636.190 3501.620 ;
        RECT 296.770 3501.420 2636.190 3501.560 ;
        RECT 296.770 3501.360 297.090 3501.420 ;
        RECT 2635.870 3501.360 2636.190 3501.420 ;
      LAYER via ;
        RECT 296.800 3501.360 297.060 3501.620 ;
        RECT 2635.900 3501.360 2636.160 3501.620 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3501.650 2636.100 3517.600 ;
        RECT 296.800 3501.330 297.060 3501.650 ;
        RECT 2635.900 3501.330 2636.160 3501.650 ;
        RECT 296.860 2048.685 297.000 3501.330 ;
        RECT 296.790 2048.315 297.070 2048.685 ;
      LAYER via2 ;
        RECT 296.790 2048.360 297.070 2048.640 ;
      LAYER met3 ;
        RECT 296.765 2048.650 297.095 2048.665 ;
        RECT 300.000 2048.650 304.000 2048.760 ;
        RECT 296.765 2048.350 304.000 2048.650 ;
        RECT 296.765 2048.335 297.095 2048.350 ;
        RECT 300.000 2048.160 304.000 2048.350 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.870 2702.900 290.190 2702.960 ;
        RECT 2311.570 2702.900 2311.890 2702.960 ;
        RECT 289.870 2702.760 2311.890 2702.900 ;
        RECT 289.870 2702.700 290.190 2702.760 ;
        RECT 2311.570 2702.700 2311.890 2702.760 ;
      LAYER via ;
        RECT 289.900 2702.700 290.160 2702.960 ;
        RECT 2311.600 2702.700 2311.860 2702.960 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 2702.990 2311.800 3517.600 ;
        RECT 289.900 2702.670 290.160 2702.990 ;
        RECT 2311.600 2702.670 2311.860 2702.990 ;
        RECT 289.960 2077.925 290.100 2702.670 ;
        RECT 289.890 2077.555 290.170 2077.925 ;
      LAYER via2 ;
        RECT 289.890 2077.600 290.170 2077.880 ;
      LAYER met3 ;
        RECT 289.865 2077.890 290.195 2077.905 ;
        RECT 300.000 2077.890 304.000 2078.000 ;
        RECT 289.865 2077.590 304.000 2077.890 ;
        RECT 289.865 2077.575 290.195 2077.590 ;
        RECT 300.000 2077.400 304.000 2077.590 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.850 3502.580 296.170 3502.640 ;
        RECT 1987.270 3502.580 1987.590 3502.640 ;
        RECT 295.850 3502.440 1987.590 3502.580 ;
        RECT 295.850 3502.380 296.170 3502.440 ;
        RECT 1987.270 3502.380 1987.590 3502.440 ;
      LAYER via ;
        RECT 295.880 3502.380 296.140 3502.640 ;
        RECT 1987.300 3502.380 1987.560 3502.640 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3502.670 1987.500 3517.600 ;
        RECT 295.880 3502.350 296.140 3502.670 ;
        RECT 1987.300 3502.350 1987.560 3502.670 ;
        RECT 295.940 2107.165 296.080 3502.350 ;
        RECT 295.870 2106.795 296.150 2107.165 ;
      LAYER via2 ;
        RECT 295.870 2106.840 296.150 2107.120 ;
      LAYER met3 ;
        RECT 295.845 2107.130 296.175 2107.145 ;
        RECT 300.000 2107.130 304.000 2107.240 ;
        RECT 295.845 2106.830 304.000 2107.130 ;
        RECT 295.845 2106.815 296.175 2106.830 ;
        RECT 300.000 2106.640 304.000 2106.830 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.930 3503.260 295.250 3503.320 ;
        RECT 1662.510 3503.260 1662.830 3503.320 ;
        RECT 294.930 3503.120 1662.830 3503.260 ;
        RECT 294.930 3503.060 295.250 3503.120 ;
        RECT 1662.510 3503.060 1662.830 3503.120 ;
      LAYER via ;
        RECT 294.960 3503.060 295.220 3503.320 ;
        RECT 1662.540 3503.060 1662.800 3503.320 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.350 1662.740 3517.600 ;
        RECT 294.960 3503.030 295.220 3503.350 ;
        RECT 1662.540 3503.030 1662.800 3503.350 ;
        RECT 295.020 2135.725 295.160 3503.030 ;
        RECT 294.950 2135.355 295.230 2135.725 ;
      LAYER via2 ;
        RECT 294.950 2135.400 295.230 2135.680 ;
      LAYER met3 ;
        RECT 294.925 2135.690 295.255 2135.705 ;
        RECT 300.000 2135.690 304.000 2135.800 ;
        RECT 294.925 2135.390 304.000 2135.690 ;
        RECT 294.925 2135.375 295.255 2135.390 ;
        RECT 300.000 2135.200 304.000 2135.390 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.470 3503.940 294.790 3504.000 ;
        RECT 1338.210 3503.940 1338.530 3504.000 ;
        RECT 294.470 3503.800 1338.530 3503.940 ;
        RECT 294.470 3503.740 294.790 3503.800 ;
        RECT 1338.210 3503.740 1338.530 3503.800 ;
      LAYER via ;
        RECT 294.500 3503.740 294.760 3504.000 ;
        RECT 1338.240 3503.740 1338.500 3504.000 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3504.030 1338.440 3517.600 ;
        RECT 294.500 3503.710 294.760 3504.030 ;
        RECT 1338.240 3503.710 1338.500 3504.030 ;
        RECT 294.560 2164.965 294.700 3503.710 ;
        RECT 294.490 2164.595 294.770 2164.965 ;
      LAYER via2 ;
        RECT 294.490 2164.640 294.770 2164.920 ;
      LAYER met3 ;
        RECT 294.465 2164.930 294.795 2164.945 ;
        RECT 300.000 2164.930 304.000 2165.040 ;
        RECT 294.465 2164.630 304.000 2164.930 ;
        RECT 294.465 2164.615 294.795 2164.630 ;
        RECT 300.000 2164.440 304.000 2164.630 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.270 441.560 285.590 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 285.270 441.420 2901.150 441.560 ;
        RECT 285.270 441.360 285.590 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 285.300 441.360 285.560 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 285.290 1643.035 285.570 1643.405 ;
        RECT 285.360 441.650 285.500 1643.035 ;
        RECT 285.300 441.330 285.560 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 285.290 1643.080 285.570 1643.360 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 285.265 1643.370 285.595 1643.385 ;
        RECT 300.000 1643.370 304.000 1643.480 ;
        RECT 285.265 1643.070 304.000 1643.370 ;
        RECT 285.265 1643.055 285.595 1643.070 ;
        RECT 300.000 1642.880 304.000 1643.070 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.550 3504.620 293.870 3504.680 ;
        RECT 1013.910 3504.620 1014.230 3504.680 ;
        RECT 293.550 3504.480 1014.230 3504.620 ;
        RECT 293.550 3504.420 293.870 3504.480 ;
        RECT 1013.910 3504.420 1014.230 3504.480 ;
      LAYER via ;
        RECT 293.580 3504.420 293.840 3504.680 ;
        RECT 1013.940 3504.420 1014.200 3504.680 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3504.710 1014.140 3517.600 ;
        RECT 293.580 3504.390 293.840 3504.710 ;
        RECT 1013.940 3504.390 1014.200 3504.710 ;
        RECT 293.640 2193.525 293.780 3504.390 ;
        RECT 293.570 2193.155 293.850 2193.525 ;
      LAYER via2 ;
        RECT 293.570 2193.200 293.850 2193.480 ;
      LAYER met3 ;
        RECT 293.545 2193.490 293.875 2193.505 ;
        RECT 300.000 2193.490 304.000 2193.600 ;
        RECT 293.545 2193.190 304.000 2193.490 ;
        RECT 293.545 2193.175 293.875 2193.190 ;
        RECT 300.000 2193.000 304.000 2193.190 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 293.090 3504.960 293.410 3505.020 ;
        RECT 689.150 3504.960 689.470 3505.020 ;
        RECT 293.090 3504.820 689.470 3504.960 ;
        RECT 293.090 3504.760 293.410 3504.820 ;
        RECT 689.150 3504.760 689.470 3504.820 ;
      LAYER via ;
        RECT 293.120 3504.760 293.380 3505.020 ;
        RECT 689.180 3504.760 689.440 3505.020 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3505.050 689.380 3517.600 ;
        RECT 293.120 3504.730 293.380 3505.050 ;
        RECT 689.180 3504.730 689.440 3505.050 ;
        RECT 293.180 2222.765 293.320 3504.730 ;
        RECT 293.110 2222.395 293.390 2222.765 ;
      LAYER via2 ;
        RECT 293.110 2222.440 293.390 2222.720 ;
      LAYER met3 ;
        RECT 293.085 2222.730 293.415 2222.745 ;
        RECT 300.000 2222.730 304.000 2222.840 ;
        RECT 293.085 2222.430 304.000 2222.730 ;
        RECT 293.085 2222.415 293.415 2222.430 ;
        RECT 300.000 2222.240 304.000 2222.430 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.170 3500.540 292.490 3500.600 ;
        RECT 364.850 3500.540 365.170 3500.600 ;
        RECT 292.170 3500.400 365.170 3500.540 ;
        RECT 292.170 3500.340 292.490 3500.400 ;
        RECT 364.850 3500.340 365.170 3500.400 ;
      LAYER via ;
        RECT 292.200 3500.340 292.460 3500.600 ;
        RECT 364.880 3500.340 365.140 3500.600 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3500.630 365.080 3517.600 ;
        RECT 292.200 3500.310 292.460 3500.630 ;
        RECT 364.880 3500.310 365.140 3500.630 ;
        RECT 292.260 2251.325 292.400 3500.310 ;
        RECT 292.190 2250.955 292.470 2251.325 ;
      LAYER via2 ;
        RECT 292.190 2251.000 292.470 2251.280 ;
      LAYER met3 ;
        RECT 292.165 2251.290 292.495 2251.305 ;
        RECT 300.000 2251.290 304.000 2251.400 ;
        RECT 292.165 2250.990 304.000 2251.290 ;
        RECT 292.165 2250.975 292.495 2250.990 ;
        RECT 300.000 2250.800 304.000 2250.990 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3498.500 40.870 3498.560 ;
        RECT 51.590 3498.500 51.910 3498.560 ;
        RECT 40.550 3498.360 51.910 3498.500 ;
        RECT 40.550 3498.300 40.870 3498.360 ;
        RECT 51.590 3498.300 51.910 3498.360 ;
        RECT 51.590 2283.680 51.910 2283.740 ;
        RECT 282.970 2283.680 283.290 2283.740 ;
        RECT 51.590 2283.540 283.290 2283.680 ;
        RECT 51.590 2283.480 51.910 2283.540 ;
        RECT 282.970 2283.480 283.290 2283.540 ;
      LAYER via ;
        RECT 40.580 3498.300 40.840 3498.560 ;
        RECT 51.620 3498.300 51.880 3498.560 ;
        RECT 51.620 2283.480 51.880 2283.740 ;
        RECT 283.000 2283.480 283.260 2283.740 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3498.590 40.780 3517.600 ;
        RECT 40.580 3498.270 40.840 3498.590 ;
        RECT 51.620 3498.270 51.880 3498.590 ;
        RECT 51.680 2283.770 51.820 3498.270 ;
        RECT 51.620 2283.450 51.880 2283.770 ;
        RECT 283.000 2283.450 283.260 2283.770 ;
        RECT 283.060 2280.565 283.200 2283.450 ;
        RECT 282.990 2280.195 283.270 2280.565 ;
      LAYER via2 ;
        RECT 282.990 2280.240 283.270 2280.520 ;
      LAYER met3 ;
        RECT 282.965 2280.530 283.295 2280.545 ;
        RECT 300.000 2280.530 304.000 2280.640 ;
        RECT 282.965 2280.230 304.000 2280.530 ;
        RECT 282.965 2280.215 283.295 2280.230 ;
        RECT 300.000 2280.040 304.000 2280.230 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 65.390 3263.900 65.710 3263.960 ;
        RECT 15.250 3263.760 65.710 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 65.390 3263.700 65.710 3263.760 ;
        RECT 65.390 2311.560 65.710 2311.620 ;
        RECT 282.510 2311.560 282.830 2311.620 ;
        RECT 65.390 2311.420 282.830 2311.560 ;
        RECT 65.390 2311.360 65.710 2311.420 ;
        RECT 282.510 2311.360 282.830 2311.420 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 65.420 3263.700 65.680 3263.960 ;
        RECT 65.420 2311.360 65.680 2311.620 ;
        RECT 282.540 2311.360 282.800 2311.620 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 65.420 3263.670 65.680 3263.990 ;
        RECT 65.480 2311.650 65.620 3263.670 ;
        RECT 65.420 2311.330 65.680 2311.650 ;
        RECT 282.540 2311.330 282.800 2311.650 ;
        RECT 282.600 2309.805 282.740 2311.330 ;
        RECT 282.530 2309.435 282.810 2309.805 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 282.530 2309.480 282.810 2309.760 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 282.505 2309.770 282.835 2309.785 ;
        RECT 300.000 2309.770 304.000 2309.880 ;
        RECT 282.505 2309.470 304.000 2309.770 ;
        RECT 282.505 2309.455 282.835 2309.470 ;
        RECT 300.000 2309.280 304.000 2309.470 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2974.220 16.950 2974.280 ;
        RECT 72.290 2974.220 72.610 2974.280 ;
        RECT 16.630 2974.080 72.610 2974.220 ;
        RECT 16.630 2974.020 16.950 2974.080 ;
        RECT 72.290 2974.020 72.610 2974.080 ;
        RECT 72.290 2339.100 72.610 2339.160 ;
        RECT 282.510 2339.100 282.830 2339.160 ;
        RECT 72.290 2338.960 282.830 2339.100 ;
        RECT 72.290 2338.900 72.610 2338.960 ;
        RECT 282.510 2338.900 282.830 2338.960 ;
      LAYER via ;
        RECT 16.660 2974.020 16.920 2974.280 ;
        RECT 72.320 2974.020 72.580 2974.280 ;
        RECT 72.320 2338.900 72.580 2339.160 ;
        RECT 282.540 2338.900 282.800 2339.160 ;
      LAYER met2 ;
        RECT 16.650 2979.915 16.930 2980.285 ;
        RECT 16.720 2974.310 16.860 2979.915 ;
        RECT 16.660 2973.990 16.920 2974.310 ;
        RECT 72.320 2973.990 72.580 2974.310 ;
        RECT 72.380 2339.190 72.520 2973.990 ;
        RECT 72.320 2338.870 72.580 2339.190 ;
        RECT 282.540 2338.870 282.800 2339.190 ;
        RECT 282.600 2338.365 282.740 2338.870 ;
        RECT 282.530 2337.995 282.810 2338.365 ;
      LAYER via2 ;
        RECT 16.650 2979.960 16.930 2980.240 ;
        RECT 282.530 2338.040 282.810 2338.320 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.625 2980.250 16.955 2980.265 ;
        RECT -4.800 2979.950 16.955 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.625 2979.935 16.955 2979.950 ;
        RECT 282.505 2338.330 282.835 2338.345 ;
        RECT 300.000 2338.330 304.000 2338.440 ;
        RECT 282.505 2338.030 304.000 2338.330 ;
        RECT 282.505 2338.015 282.835 2338.030 ;
        RECT 300.000 2337.840 304.000 2338.030 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 2373.440 19.250 2373.500 ;
        RECT 282.510 2373.440 282.830 2373.500 ;
        RECT 18.930 2373.300 282.830 2373.440 ;
        RECT 18.930 2373.240 19.250 2373.300 ;
        RECT 282.510 2373.240 282.830 2373.300 ;
      LAYER via ;
        RECT 18.960 2373.240 19.220 2373.500 ;
        RECT 282.540 2373.240 282.800 2373.500 ;
      LAYER met2 ;
        RECT 18.950 2692.955 19.230 2693.325 ;
        RECT 19.020 2373.530 19.160 2692.955 ;
        RECT 18.960 2373.210 19.220 2373.530 ;
        RECT 282.540 2373.210 282.800 2373.530 ;
        RECT 282.600 2367.605 282.740 2373.210 ;
        RECT 282.530 2367.235 282.810 2367.605 ;
      LAYER via2 ;
        RECT 18.950 2693.000 19.230 2693.280 ;
        RECT 282.530 2367.280 282.810 2367.560 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 18.925 2693.290 19.255 2693.305 ;
        RECT -4.800 2692.990 19.255 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 18.925 2692.975 19.255 2692.990 ;
        RECT 282.505 2367.570 282.835 2367.585 ;
        RECT 300.000 2367.570 304.000 2367.680 ;
        RECT 282.505 2367.270 304.000 2367.570 ;
        RECT 282.505 2367.255 282.835 2367.270 ;
        RECT 300.000 2367.080 304.000 2367.270 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 2400.980 14.650 2401.040 ;
        RECT 282.510 2400.980 282.830 2401.040 ;
        RECT 14.330 2400.840 282.830 2400.980 ;
        RECT 14.330 2400.780 14.650 2400.840 ;
        RECT 282.510 2400.780 282.830 2400.840 ;
      LAYER via ;
        RECT 14.360 2400.780 14.620 2401.040 ;
        RECT 282.540 2400.780 282.800 2401.040 ;
      LAYER met2 ;
        RECT 14.350 2405.315 14.630 2405.685 ;
        RECT 14.420 2401.070 14.560 2405.315 ;
        RECT 14.360 2400.750 14.620 2401.070 ;
        RECT 282.540 2400.750 282.800 2401.070 ;
        RECT 282.600 2396.165 282.740 2400.750 ;
        RECT 282.530 2395.795 282.810 2396.165 ;
      LAYER via2 ;
        RECT 14.350 2405.360 14.630 2405.640 ;
        RECT 282.530 2395.840 282.810 2396.120 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 14.325 2405.650 14.655 2405.665 ;
        RECT -4.800 2405.350 14.655 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 14.325 2405.335 14.655 2405.350 ;
        RECT 282.505 2396.130 282.835 2396.145 ;
        RECT 300.000 2396.130 304.000 2396.240 ;
        RECT 282.505 2395.830 304.000 2396.130 ;
        RECT 282.505 2395.815 282.835 2395.830 ;
        RECT 300.000 2395.640 304.000 2395.830 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.390 2422.060 19.710 2422.120 ;
        RECT 283.430 2422.060 283.750 2422.120 ;
        RECT 19.390 2421.920 283.750 2422.060 ;
        RECT 19.390 2421.860 19.710 2421.920 ;
        RECT 283.430 2421.860 283.750 2421.920 ;
      LAYER via ;
        RECT 19.420 2421.860 19.680 2422.120 ;
        RECT 283.460 2421.860 283.720 2422.120 ;
      LAYER met2 ;
        RECT 283.450 2425.035 283.730 2425.405 ;
        RECT 283.520 2422.150 283.660 2425.035 ;
        RECT 19.420 2421.830 19.680 2422.150 ;
        RECT 283.460 2421.830 283.720 2422.150 ;
        RECT 19.480 2118.725 19.620 2421.830 ;
        RECT 19.410 2118.355 19.690 2118.725 ;
      LAYER via2 ;
        RECT 283.450 2425.080 283.730 2425.360 ;
        RECT 19.410 2118.400 19.690 2118.680 ;
      LAYER met3 ;
        RECT 283.425 2425.370 283.755 2425.385 ;
        RECT 300.000 2425.370 304.000 2425.480 ;
        RECT 283.425 2425.070 304.000 2425.370 ;
        RECT 283.425 2425.055 283.755 2425.070 ;
        RECT 300.000 2424.880 304.000 2425.070 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 19.385 2118.690 19.715 2118.705 ;
        RECT -4.800 2118.390 19.715 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 19.385 2118.375 19.715 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.190 2449.600 79.510 2449.660 ;
        RECT 283.430 2449.600 283.750 2449.660 ;
        RECT 79.190 2449.460 283.750 2449.600 ;
        RECT 79.190 2449.400 79.510 2449.460 ;
        RECT 283.430 2449.400 283.750 2449.460 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 79.190 1835.220 79.510 1835.280 ;
        RECT 15.710 1835.080 79.510 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 79.190 1835.020 79.510 1835.080 ;
      LAYER via ;
        RECT 79.220 2449.400 79.480 2449.660 ;
        RECT 283.460 2449.400 283.720 2449.660 ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 79.220 1835.020 79.480 1835.280 ;
      LAYER met2 ;
        RECT 283.450 2453.595 283.730 2453.965 ;
        RECT 283.520 2449.690 283.660 2453.595 ;
        RECT 79.220 2449.370 79.480 2449.690 ;
        RECT 283.460 2449.370 283.720 2449.690 ;
        RECT 79.280 1835.310 79.420 2449.370 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 79.220 1834.990 79.480 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 283.450 2453.640 283.730 2453.920 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 283.425 2453.930 283.755 2453.945 ;
        RECT 300.000 2453.930 304.000 2454.040 ;
        RECT 283.425 2453.630 304.000 2453.930 ;
        RECT 283.425 2453.615 283.755 2453.630 ;
        RECT 300.000 2453.440 304.000 2453.630 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 287.110 676.160 287.430 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 287.110 676.020 2901.150 676.160 ;
        RECT 287.110 675.960 287.430 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 287.140 675.960 287.400 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 287.130 1672.275 287.410 1672.645 ;
        RECT 287.200 676.250 287.340 1672.275 ;
        RECT 287.140 675.930 287.400 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 287.130 1672.320 287.410 1672.600 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 287.105 1672.610 287.435 1672.625 ;
        RECT 300.000 1672.610 304.000 1672.720 ;
        RECT 287.105 1672.310 304.000 1672.610 ;
        RECT 287.105 1672.295 287.435 1672.310 ;
        RECT 300.000 1672.120 304.000 1672.310 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 100.350 2477.480 100.670 2477.540 ;
        RECT 287.110 2477.480 287.430 2477.540 ;
        RECT 100.350 2477.340 287.430 2477.480 ;
        RECT 100.350 2477.280 100.670 2477.340 ;
        RECT 287.110 2477.280 287.430 2477.340 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 100.350 1545.540 100.670 1545.600 ;
        RECT 16.630 1545.400 100.670 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 100.350 1545.340 100.670 1545.400 ;
      LAYER via ;
        RECT 100.380 2477.280 100.640 2477.540 ;
        RECT 287.140 2477.280 287.400 2477.540 ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 100.380 1545.340 100.640 1545.600 ;
      LAYER met2 ;
        RECT 287.130 2482.835 287.410 2483.205 ;
        RECT 287.200 2477.570 287.340 2482.835 ;
        RECT 100.380 2477.250 100.640 2477.570 ;
        RECT 287.140 2477.250 287.400 2477.570 ;
        RECT 100.440 1545.630 100.580 2477.250 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 100.380 1545.310 100.640 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 287.130 2482.880 287.410 2483.160 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 287.105 2483.170 287.435 2483.185 ;
        RECT 300.000 2483.170 304.000 2483.280 ;
        RECT 287.105 2482.870 304.000 2483.170 ;
        RECT 287.105 2482.855 287.435 2482.870 ;
        RECT 300.000 2482.680 304.000 2482.870 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 141.750 2511.820 142.070 2511.880 ;
        RECT 287.110 2511.820 287.430 2511.880 ;
        RECT 141.750 2511.680 287.430 2511.820 ;
        RECT 141.750 2511.620 142.070 2511.680 ;
        RECT 287.110 2511.620 287.430 2511.680 ;
        RECT 14.330 1331.680 14.650 1331.740 ;
        RECT 141.750 1331.680 142.070 1331.740 ;
        RECT 14.330 1331.540 142.070 1331.680 ;
        RECT 14.330 1331.480 14.650 1331.540 ;
        RECT 141.750 1331.480 142.070 1331.540 ;
      LAYER via ;
        RECT 141.780 2511.620 142.040 2511.880 ;
        RECT 287.140 2511.620 287.400 2511.880 ;
        RECT 14.360 1331.480 14.620 1331.740 ;
        RECT 141.780 1331.480 142.040 1331.740 ;
      LAYER met2 ;
        RECT 287.130 2512.075 287.410 2512.445 ;
        RECT 287.200 2511.910 287.340 2512.075 ;
        RECT 141.780 2511.590 142.040 2511.910 ;
        RECT 287.140 2511.590 287.400 2511.910 ;
        RECT 141.840 1331.770 141.980 2511.590 ;
        RECT 14.360 1331.450 14.620 1331.770 ;
        RECT 141.780 1331.450 142.040 1331.770 ;
        RECT 14.420 1328.565 14.560 1331.450 ;
        RECT 14.350 1328.195 14.630 1328.565 ;
      LAYER via2 ;
        RECT 287.130 2512.120 287.410 2512.400 ;
        RECT 14.350 1328.240 14.630 1328.520 ;
      LAYER met3 ;
        RECT 287.105 2512.410 287.435 2512.425 ;
        RECT 300.000 2512.410 304.000 2512.520 ;
        RECT 287.105 2512.110 304.000 2512.410 ;
        RECT 287.105 2512.095 287.435 2512.110 ;
        RECT 300.000 2511.920 304.000 2512.110 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 14.325 1328.530 14.655 1328.545 ;
        RECT -4.800 1328.230 14.655 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 14.325 1328.215 14.655 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 169.350 2539.360 169.670 2539.420 ;
        RECT 287.110 2539.360 287.430 2539.420 ;
        RECT 169.350 2539.220 287.430 2539.360 ;
        RECT 169.350 2539.160 169.670 2539.220 ;
        RECT 287.110 2539.160 287.430 2539.220 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 169.350 1117.820 169.670 1117.880 ;
        RECT 15.710 1117.680 169.670 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 169.350 1117.620 169.670 1117.680 ;
      LAYER via ;
        RECT 169.380 2539.160 169.640 2539.420 ;
        RECT 287.140 2539.160 287.400 2539.420 ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 169.380 1117.620 169.640 1117.880 ;
      LAYER met2 ;
        RECT 287.130 2540.635 287.410 2541.005 ;
        RECT 287.200 2539.450 287.340 2540.635 ;
        RECT 169.380 2539.130 169.640 2539.450 ;
        RECT 287.140 2539.130 287.400 2539.450 ;
        RECT 169.440 1117.910 169.580 2539.130 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 169.380 1117.590 169.640 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 287.130 2540.680 287.410 2540.960 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 287.105 2540.970 287.435 2540.985 ;
        RECT 300.000 2540.970 304.000 2541.080 ;
        RECT 287.105 2540.670 304.000 2540.970 ;
        RECT 287.105 2540.655 287.435 2540.670 ;
        RECT 300.000 2540.480 304.000 2540.670 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 2566.900 176.110 2566.960 ;
        RECT 287.110 2566.900 287.430 2566.960 ;
        RECT 175.790 2566.760 287.430 2566.900 ;
        RECT 175.790 2566.700 176.110 2566.760 ;
        RECT 287.110 2566.700 287.430 2566.760 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 175.790 903.960 176.110 904.020 ;
        RECT 16.170 903.820 176.110 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 175.790 903.760 176.110 903.820 ;
      LAYER via ;
        RECT 175.820 2566.700 176.080 2566.960 ;
        RECT 287.140 2566.700 287.400 2566.960 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 175.820 903.760 176.080 904.020 ;
      LAYER met2 ;
        RECT 287.130 2569.875 287.410 2570.245 ;
        RECT 287.200 2566.990 287.340 2569.875 ;
        RECT 175.820 2566.670 176.080 2566.990 ;
        RECT 287.140 2566.670 287.400 2566.990 ;
        RECT 175.880 904.050 176.020 2566.670 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 175.820 903.730 176.080 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 287.130 2569.920 287.410 2570.200 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT 287.105 2570.210 287.435 2570.225 ;
        RECT 300.000 2570.210 304.000 2570.320 ;
        RECT 287.105 2569.910 304.000 2570.210 ;
        RECT 287.105 2569.895 287.435 2569.910 ;
        RECT 300.000 2569.720 304.000 2569.910 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 217.190 2594.780 217.510 2594.840 ;
        RECT 287.110 2594.780 287.430 2594.840 ;
        RECT 217.190 2594.640 287.430 2594.780 ;
        RECT 217.190 2594.580 217.510 2594.640 ;
        RECT 287.110 2594.580 287.430 2594.640 ;
        RECT 16.170 682.960 16.490 683.020 ;
        RECT 217.190 682.960 217.510 683.020 ;
        RECT 16.170 682.820 217.510 682.960 ;
        RECT 16.170 682.760 16.490 682.820 ;
        RECT 217.190 682.760 217.510 682.820 ;
      LAYER via ;
        RECT 217.220 2594.580 217.480 2594.840 ;
        RECT 287.140 2594.580 287.400 2594.840 ;
        RECT 16.200 682.760 16.460 683.020 ;
        RECT 217.220 682.760 217.480 683.020 ;
      LAYER met2 ;
        RECT 287.130 2598.435 287.410 2598.805 ;
        RECT 287.200 2594.870 287.340 2598.435 ;
        RECT 217.220 2594.550 217.480 2594.870 ;
        RECT 287.140 2594.550 287.400 2594.870 ;
        RECT 217.280 683.050 217.420 2594.550 ;
        RECT 16.200 682.730 16.460 683.050 ;
        RECT 217.220 682.730 217.480 683.050 ;
        RECT 16.260 681.885 16.400 682.730 ;
        RECT 16.190 681.515 16.470 681.885 ;
      LAYER via2 ;
        RECT 287.130 2598.480 287.410 2598.760 ;
        RECT 16.190 681.560 16.470 681.840 ;
      LAYER met3 ;
        RECT 287.105 2598.770 287.435 2598.785 ;
        RECT 300.000 2598.770 304.000 2598.880 ;
        RECT 287.105 2598.470 304.000 2598.770 ;
        RECT 287.105 2598.455 287.435 2598.470 ;
        RECT 300.000 2598.280 304.000 2598.470 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 16.165 681.850 16.495 681.865 ;
        RECT -4.800 681.550 16.495 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 16.165 681.535 16.495 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 230.990 2622.320 231.310 2622.380 ;
        RECT 287.110 2622.320 287.430 2622.380 ;
        RECT 230.990 2622.180 287.430 2622.320 ;
        RECT 230.990 2622.120 231.310 2622.180 ;
        RECT 287.110 2622.120 287.430 2622.180 ;
        RECT 17.090 469.100 17.410 469.160 ;
        RECT 230.990 469.100 231.310 469.160 ;
        RECT 17.090 468.960 231.310 469.100 ;
        RECT 17.090 468.900 17.410 468.960 ;
        RECT 230.990 468.900 231.310 468.960 ;
      LAYER via ;
        RECT 231.020 2622.120 231.280 2622.380 ;
        RECT 287.140 2622.120 287.400 2622.380 ;
        RECT 17.120 468.900 17.380 469.160 ;
        RECT 231.020 468.900 231.280 469.160 ;
      LAYER met2 ;
        RECT 287.130 2627.675 287.410 2628.045 ;
        RECT 287.200 2622.410 287.340 2627.675 ;
        RECT 231.020 2622.090 231.280 2622.410 ;
        RECT 287.140 2622.090 287.400 2622.410 ;
        RECT 231.080 469.190 231.220 2622.090 ;
        RECT 17.120 468.870 17.380 469.190 ;
        RECT 231.020 468.870 231.280 469.190 ;
        RECT 17.180 466.325 17.320 468.870 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 287.130 2627.720 287.410 2628.000 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT 287.105 2628.010 287.435 2628.025 ;
        RECT 300.000 2628.010 304.000 2628.120 ;
        RECT 287.105 2627.710 304.000 2628.010 ;
        RECT 287.105 2627.695 287.435 2627.710 ;
        RECT 300.000 2627.520 304.000 2627.710 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 244.790 2657.000 245.110 2657.060 ;
        RECT 287.110 2657.000 287.430 2657.060 ;
        RECT 244.790 2656.860 287.430 2657.000 ;
        RECT 244.790 2656.800 245.110 2656.860 ;
        RECT 287.110 2656.800 287.430 2656.860 ;
        RECT 17.090 255.240 17.410 255.300 ;
        RECT 244.790 255.240 245.110 255.300 ;
        RECT 17.090 255.100 245.110 255.240 ;
        RECT 17.090 255.040 17.410 255.100 ;
        RECT 244.790 255.040 245.110 255.100 ;
      LAYER via ;
        RECT 244.820 2656.800 245.080 2657.060 ;
        RECT 287.140 2656.800 287.400 2657.060 ;
        RECT 17.120 255.040 17.380 255.300 ;
        RECT 244.820 255.040 245.080 255.300 ;
      LAYER met2 ;
        RECT 244.820 2656.770 245.080 2657.090 ;
        RECT 287.130 2656.915 287.410 2657.285 ;
        RECT 287.140 2656.770 287.400 2656.915 ;
        RECT 244.880 255.330 245.020 2656.770 ;
        RECT 17.120 255.010 17.380 255.330 ;
        RECT 244.820 255.010 245.080 255.330 ;
        RECT 17.180 250.765 17.320 255.010 ;
        RECT 17.110 250.395 17.390 250.765 ;
      LAYER via2 ;
        RECT 287.130 2656.960 287.410 2657.240 ;
        RECT 17.110 250.440 17.390 250.720 ;
      LAYER met3 ;
        RECT 287.105 2657.250 287.435 2657.265 ;
        RECT 300.000 2657.250 304.000 2657.360 ;
        RECT 287.105 2656.950 304.000 2657.250 ;
        RECT 287.105 2656.935 287.435 2656.950 ;
        RECT 300.000 2656.760 304.000 2656.950 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 17.085 250.730 17.415 250.745 ;
        RECT -4.800 250.430 17.415 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 17.085 250.415 17.415 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 99.890 2684.200 100.210 2684.260 ;
        RECT 287.110 2684.200 287.430 2684.260 ;
        RECT 99.890 2684.060 287.430 2684.200 ;
        RECT 99.890 2684.000 100.210 2684.060 ;
        RECT 287.110 2684.000 287.430 2684.060 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 99.890 41.380 100.210 41.440 ;
        RECT 17.090 41.240 100.210 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 99.890 41.180 100.210 41.240 ;
      LAYER via ;
        RECT 99.920 2684.000 100.180 2684.260 ;
        RECT 287.140 2684.000 287.400 2684.260 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 99.920 41.180 100.180 41.440 ;
      LAYER met2 ;
        RECT 287.130 2685.475 287.410 2685.845 ;
        RECT 287.200 2684.290 287.340 2685.475 ;
        RECT 99.920 2683.970 100.180 2684.290 ;
        RECT 287.140 2683.970 287.400 2684.290 ;
        RECT 99.980 41.470 100.120 2683.970 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 99.920 41.150 100.180 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 287.130 2685.520 287.410 2685.800 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 287.105 2685.810 287.435 2685.825 ;
        RECT 300.000 2685.810 304.000 2685.920 ;
        RECT 287.105 2685.510 304.000 2685.810 ;
        RECT 287.105 2685.495 287.435 2685.510 ;
        RECT 300.000 2685.320 304.000 2685.510 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 346.910 905.320 347.230 905.380 ;
        RECT 386.010 905.320 386.330 905.380 ;
        RECT 346.910 905.180 386.330 905.320 ;
        RECT 346.910 905.120 347.230 905.180 ;
        RECT 386.010 905.120 386.330 905.180 ;
      LAYER via ;
        RECT 346.940 905.120 347.200 905.380 ;
        RECT 386.040 905.120 386.300 905.380 ;
      LAYER met2 ;
        RECT 555.310 907.275 555.590 907.645 ;
        RECT 346.940 905.090 347.200 905.410 ;
        RECT 386.030 905.235 386.310 905.605 ;
        RECT 386.040 905.090 386.300 905.235 ;
        RECT 347.000 904.925 347.140 905.090 ;
        RECT 346.930 904.555 347.210 904.925 ;
        RECT 555.380 904.245 555.520 907.275 ;
        RECT 641.330 904.810 641.610 904.925 ;
        RECT 642.250 904.810 642.530 904.925 ;
        RECT 641.330 904.670 642.530 904.810 ;
        RECT 641.330 904.555 641.610 904.670 ;
        RECT 642.250 904.555 642.530 904.670 ;
        RECT 555.310 903.875 555.590 904.245 ;
      LAYER via2 ;
        RECT 555.310 907.320 555.590 907.600 ;
        RECT 386.030 905.280 386.310 905.560 ;
        RECT 346.930 904.600 347.210 904.880 ;
        RECT 641.330 904.600 641.610 904.880 ;
        RECT 642.250 904.600 642.530 904.880 ;
        RECT 555.310 903.920 555.590 904.200 ;
      LAYER met3 ;
        RECT 287.310 1701.170 287.690 1701.180 ;
        RECT 300.000 1701.170 304.000 1701.280 ;
        RECT 287.310 1700.870 304.000 1701.170 ;
        RECT 287.310 1700.860 287.690 1700.870 ;
        RECT 300.000 1700.680 304.000 1700.870 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2916.710 909.350 2924.800 909.650 ;
        RECT 531.110 907.610 531.490 907.620 ;
        RECT 555.285 907.610 555.615 907.625 ;
        RECT 531.110 907.310 555.615 907.610 ;
        RECT 531.110 907.300 531.490 907.310 ;
        RECT 555.285 907.295 555.615 907.310 ;
        RECT 531.110 906.250 531.490 906.260 ;
        RECT 497.110 905.950 531.490 906.250 ;
        RECT 287.310 905.570 287.690 905.580 ;
        RECT 386.005 905.570 386.335 905.585 ;
        RECT 287.310 905.270 304.210 905.570 ;
        RECT 287.310 905.260 287.690 905.270 ;
        RECT 303.910 904.890 304.210 905.270 ;
        RECT 386.005 905.270 410.930 905.570 ;
        RECT 386.005 905.255 386.335 905.270 ;
        RECT 346.905 904.890 347.235 904.905 ;
        RECT 303.910 904.590 347.235 904.890 ;
        RECT 346.905 904.575 347.235 904.590 ;
        RECT 410.630 904.210 410.930 905.270 ;
        RECT 482.350 904.890 482.730 904.900 ;
        RECT 497.110 904.890 497.410 905.950 ;
        RECT 531.110 905.940 531.490 905.950 ;
        RECT 834.750 905.270 882.890 905.570 ;
        RECT 641.305 904.890 641.635 904.905 ;
        RECT 482.350 904.590 497.410 904.890 ;
        RECT 593.710 904.590 641.635 904.890 ;
        RECT 482.350 904.580 482.730 904.590 ;
        RECT 482.350 904.210 482.730 904.220 ;
        RECT 410.630 903.910 482.730 904.210 ;
        RECT 482.350 903.900 482.730 903.910 ;
        RECT 555.285 904.210 555.615 904.225 ;
        RECT 593.710 904.210 594.010 904.590 ;
        RECT 641.305 904.575 641.635 904.590 ;
        RECT 642.225 904.890 642.555 904.905 ;
        RECT 642.225 904.590 689.690 904.890 ;
        RECT 642.225 904.575 642.555 904.590 ;
        RECT 555.285 903.910 594.010 904.210 ;
        RECT 689.390 904.210 689.690 904.590 ;
        RECT 834.750 904.210 835.050 905.270 ;
        RECT 689.390 903.910 835.050 904.210 ;
        RECT 882.590 904.210 882.890 905.270 ;
        RECT 931.350 905.270 979.490 905.570 ;
        RECT 931.350 904.210 931.650 905.270 ;
        RECT 882.590 903.910 931.650 904.210 ;
        RECT 979.190 904.210 979.490 905.270 ;
        RECT 1027.950 905.270 1076.090 905.570 ;
        RECT 1027.950 904.210 1028.250 905.270 ;
        RECT 979.190 903.910 1028.250 904.210 ;
        RECT 1075.790 904.210 1076.090 905.270 ;
        RECT 1124.550 905.270 1172.690 905.570 ;
        RECT 1124.550 904.210 1124.850 905.270 ;
        RECT 1075.790 903.910 1124.850 904.210 ;
        RECT 1172.390 904.210 1172.690 905.270 ;
        RECT 1221.150 905.270 1269.290 905.570 ;
        RECT 1221.150 904.210 1221.450 905.270 ;
        RECT 1172.390 903.910 1221.450 904.210 ;
        RECT 1268.990 904.210 1269.290 905.270 ;
        RECT 1317.750 905.270 1365.890 905.570 ;
        RECT 1317.750 904.210 1318.050 905.270 ;
        RECT 1268.990 903.910 1318.050 904.210 ;
        RECT 1365.590 904.210 1365.890 905.270 ;
        RECT 1386.750 905.270 1483.650 905.570 ;
        RECT 1386.750 904.210 1387.050 905.270 ;
        RECT 1483.350 904.890 1483.650 905.270 ;
        RECT 1532.110 905.270 1580.250 905.570 ;
        RECT 1483.350 904.590 1531.490 904.890 ;
        RECT 1365.590 903.910 1387.050 904.210 ;
        RECT 1531.190 904.210 1531.490 904.590 ;
        RECT 1532.110 904.210 1532.410 905.270 ;
        RECT 1579.950 904.890 1580.250 905.270 ;
        RECT 1628.710 905.270 1676.850 905.570 ;
        RECT 1579.950 904.590 1628.090 904.890 ;
        RECT 1531.190 903.910 1532.410 904.210 ;
        RECT 1627.790 904.210 1628.090 904.590 ;
        RECT 1628.710 904.210 1629.010 905.270 ;
        RECT 1676.550 904.890 1676.850 905.270 ;
        RECT 1725.310 905.270 1773.450 905.570 ;
        RECT 1676.550 904.590 1724.690 904.890 ;
        RECT 1627.790 903.910 1629.010 904.210 ;
        RECT 1724.390 904.210 1724.690 904.590 ;
        RECT 1725.310 904.210 1725.610 905.270 ;
        RECT 1773.150 904.890 1773.450 905.270 ;
        RECT 1821.910 905.270 1870.050 905.570 ;
        RECT 1773.150 904.590 1821.290 904.890 ;
        RECT 1724.390 903.910 1725.610 904.210 ;
        RECT 1820.990 904.210 1821.290 904.590 ;
        RECT 1821.910 904.210 1822.210 905.270 ;
        RECT 1869.750 904.890 1870.050 905.270 ;
        RECT 1918.510 905.270 1966.650 905.570 ;
        RECT 1869.750 904.590 1917.890 904.890 ;
        RECT 1820.990 903.910 1822.210 904.210 ;
        RECT 1917.590 904.210 1917.890 904.590 ;
        RECT 1918.510 904.210 1918.810 905.270 ;
        RECT 1966.350 904.890 1966.650 905.270 ;
        RECT 2015.110 905.270 2063.250 905.570 ;
        RECT 1966.350 904.590 2014.490 904.890 ;
        RECT 1917.590 903.910 1918.810 904.210 ;
        RECT 2014.190 904.210 2014.490 904.590 ;
        RECT 2015.110 904.210 2015.410 905.270 ;
        RECT 2062.950 904.890 2063.250 905.270 ;
        RECT 2111.710 905.270 2159.850 905.570 ;
        RECT 2062.950 904.590 2111.090 904.890 ;
        RECT 2014.190 903.910 2015.410 904.210 ;
        RECT 2110.790 904.210 2111.090 904.590 ;
        RECT 2111.710 904.210 2112.010 905.270 ;
        RECT 2159.550 904.890 2159.850 905.270 ;
        RECT 2208.310 905.270 2256.450 905.570 ;
        RECT 2159.550 904.590 2207.690 904.890 ;
        RECT 2110.790 903.910 2112.010 904.210 ;
        RECT 2207.390 904.210 2207.690 904.590 ;
        RECT 2208.310 904.210 2208.610 905.270 ;
        RECT 2256.150 904.890 2256.450 905.270 ;
        RECT 2304.910 905.270 2353.050 905.570 ;
        RECT 2256.150 904.590 2304.290 904.890 ;
        RECT 2207.390 903.910 2208.610 904.210 ;
        RECT 2303.990 904.210 2304.290 904.590 ;
        RECT 2304.910 904.210 2305.210 905.270 ;
        RECT 2352.750 904.890 2353.050 905.270 ;
        RECT 2401.510 905.270 2449.650 905.570 ;
        RECT 2352.750 904.590 2400.890 904.890 ;
        RECT 2303.990 903.910 2305.210 904.210 ;
        RECT 2400.590 904.210 2400.890 904.590 ;
        RECT 2401.510 904.210 2401.810 905.270 ;
        RECT 2449.350 904.890 2449.650 905.270 ;
        RECT 2498.110 905.270 2546.250 905.570 ;
        RECT 2449.350 904.590 2497.490 904.890 ;
        RECT 2400.590 903.910 2401.810 904.210 ;
        RECT 2497.190 904.210 2497.490 904.590 ;
        RECT 2498.110 904.210 2498.410 905.270 ;
        RECT 2545.950 904.890 2546.250 905.270 ;
        RECT 2594.710 905.270 2642.850 905.570 ;
        RECT 2545.950 904.590 2594.090 904.890 ;
        RECT 2497.190 903.910 2498.410 904.210 ;
        RECT 2593.790 904.210 2594.090 904.590 ;
        RECT 2594.710 904.210 2595.010 905.270 ;
        RECT 2642.550 904.890 2642.850 905.270 ;
        RECT 2691.310 905.270 2739.450 905.570 ;
        RECT 2642.550 904.590 2690.690 904.890 ;
        RECT 2593.790 903.910 2595.010 904.210 ;
        RECT 2690.390 904.210 2690.690 904.590 ;
        RECT 2691.310 904.210 2691.610 905.270 ;
        RECT 2739.150 904.890 2739.450 905.270 ;
        RECT 2787.910 905.270 2836.050 905.570 ;
        RECT 2739.150 904.590 2787.290 904.890 ;
        RECT 2690.390 903.910 2691.610 904.210 ;
        RECT 2786.990 904.210 2787.290 904.590 ;
        RECT 2787.910 904.210 2788.210 905.270 ;
        RECT 2835.750 904.890 2836.050 905.270 ;
        RECT 2916.710 904.890 2917.010 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
        RECT 2835.750 904.590 2883.890 904.890 ;
        RECT 2786.990 903.910 2788.210 904.210 ;
        RECT 2883.590 904.210 2883.890 904.590 ;
        RECT 2884.510 904.590 2917.010 904.890 ;
        RECT 2884.510 904.210 2884.810 904.590 ;
        RECT 2883.590 903.910 2884.810 904.210 ;
        RECT 555.285 903.895 555.615 903.910 ;
      LAYER via3 ;
        RECT 287.340 1700.860 287.660 1701.180 ;
        RECT 531.140 907.300 531.460 907.620 ;
        RECT 287.340 905.260 287.660 905.580 ;
        RECT 482.380 904.580 482.700 904.900 ;
        RECT 531.140 905.940 531.460 906.260 ;
        RECT 482.380 903.900 482.700 904.220 ;
      LAYER met4 ;
        RECT 287.335 1700.855 287.665 1701.185 ;
        RECT 287.350 905.585 287.650 1700.855 ;
        RECT 531.135 907.295 531.465 907.625 ;
        RECT 531.150 906.265 531.450 907.295 ;
        RECT 531.135 905.935 531.465 906.265 ;
        RECT 287.335 905.255 287.665 905.585 ;
        RECT 482.375 904.575 482.705 904.905 ;
        RECT 482.390 904.225 482.690 904.575 ;
        RECT 482.375 903.895 482.705 904.225 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 331.270 1139.920 331.590 1139.980 ;
        RECT 379.110 1139.920 379.430 1139.980 ;
        RECT 331.270 1139.780 379.430 1139.920 ;
        RECT 331.270 1139.720 331.590 1139.780 ;
        RECT 379.110 1139.720 379.430 1139.780 ;
        RECT 737.910 1139.580 738.230 1139.640 ;
        RECT 772.410 1139.580 772.730 1139.640 ;
        RECT 737.910 1139.440 772.730 1139.580 ;
        RECT 737.910 1139.380 738.230 1139.440 ;
        RECT 772.410 1139.380 772.730 1139.440 ;
        RECT 579.670 1138.900 579.990 1138.960 ;
        RECT 593.930 1138.900 594.250 1138.960 ;
        RECT 579.670 1138.760 594.250 1138.900 ;
        RECT 579.670 1138.700 579.990 1138.760 ;
        RECT 593.930 1138.700 594.250 1138.760 ;
      LAYER via ;
        RECT 331.300 1139.720 331.560 1139.980 ;
        RECT 379.140 1139.720 379.400 1139.980 ;
        RECT 737.940 1139.380 738.200 1139.640 ;
        RECT 772.440 1139.380 772.700 1139.640 ;
        RECT 579.700 1138.700 579.960 1138.960 ;
        RECT 593.960 1138.700 594.220 1138.960 ;
      LAYER met2 ;
        RECT 555.310 1141.875 555.590 1142.245 ;
        RECT 331.300 1139.690 331.560 1140.010 ;
        RECT 379.130 1139.835 379.410 1140.205 ;
        RECT 379.140 1139.690 379.400 1139.835 ;
        RECT 331.360 1139.525 331.500 1139.690 ;
        RECT 331.290 1139.155 331.570 1139.525 ;
        RECT 555.380 1138.845 555.520 1141.875 ;
        RECT 675.830 1141.195 676.110 1141.565 ;
        RECT 593.950 1139.835 594.230 1140.205 ;
        RECT 594.020 1138.990 594.160 1139.835 ;
        RECT 675.900 1139.525 676.040 1141.195 ;
        RECT 700.210 1140.515 700.490 1140.885 ;
        RECT 675.830 1139.155 676.110 1139.525 ;
        RECT 579.700 1138.845 579.960 1138.990 ;
        RECT 555.310 1138.475 555.590 1138.845 ;
        RECT 579.690 1138.475 579.970 1138.845 ;
        RECT 593.960 1138.670 594.220 1138.990 ;
        RECT 700.280 1138.845 700.420 1140.515 ;
        RECT 772.430 1139.835 772.710 1140.205 ;
        RECT 772.500 1139.670 772.640 1139.835 ;
        RECT 737.940 1139.525 738.200 1139.670 ;
        RECT 737.930 1139.155 738.210 1139.525 ;
        RECT 772.440 1139.350 772.700 1139.670 ;
        RECT 700.210 1138.475 700.490 1138.845 ;
      LAYER via2 ;
        RECT 555.310 1141.920 555.590 1142.200 ;
        RECT 379.130 1139.880 379.410 1140.160 ;
        RECT 331.290 1139.200 331.570 1139.480 ;
        RECT 675.830 1141.240 676.110 1141.520 ;
        RECT 593.950 1139.880 594.230 1140.160 ;
        RECT 700.210 1140.560 700.490 1140.840 ;
        RECT 675.830 1139.200 676.110 1139.480 ;
        RECT 555.310 1138.520 555.590 1138.800 ;
        RECT 579.690 1138.520 579.970 1138.800 ;
        RECT 772.430 1139.880 772.710 1140.160 ;
        RECT 737.930 1139.200 738.210 1139.480 ;
        RECT 700.210 1138.520 700.490 1138.800 ;
      LAYER met3 ;
        RECT 285.470 1730.410 285.850 1730.420 ;
        RECT 300.000 1730.410 304.000 1730.520 ;
        RECT 285.470 1730.110 304.000 1730.410 ;
        RECT 285.470 1730.100 285.850 1730.110 ;
        RECT 300.000 1729.920 304.000 1730.110 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2916.710 1143.950 2924.800 1144.250 ;
        RECT 531.110 1142.210 531.490 1142.220 ;
        RECT 555.285 1142.210 555.615 1142.225 ;
        RECT 531.110 1141.910 555.615 1142.210 ;
        RECT 531.110 1141.900 531.490 1141.910 ;
        RECT 555.285 1141.895 555.615 1141.910 ;
        RECT 627.710 1141.530 628.090 1141.540 ;
        RECT 675.805 1141.530 676.135 1141.545 ;
        RECT 627.710 1141.230 676.135 1141.530 ;
        RECT 627.710 1141.220 628.090 1141.230 ;
        RECT 675.805 1141.215 676.135 1141.230 ;
        RECT 531.110 1140.850 531.490 1140.860 ;
        RECT 700.185 1140.850 700.515 1140.865 ;
        RECT 497.110 1140.550 531.490 1140.850 ;
        RECT 285.470 1140.170 285.850 1140.180 ;
        RECT 379.105 1140.170 379.435 1140.185 ;
        RECT 285.470 1139.870 304.210 1140.170 ;
        RECT 285.470 1139.860 285.850 1139.870 ;
        RECT 303.910 1139.490 304.210 1139.870 ;
        RECT 379.105 1139.870 410.930 1140.170 ;
        RECT 379.105 1139.855 379.435 1139.870 ;
        RECT 331.265 1139.490 331.595 1139.505 ;
        RECT 303.910 1139.190 331.595 1139.490 ;
        RECT 331.265 1139.175 331.595 1139.190 ;
        RECT 410.630 1138.810 410.930 1139.870 ;
        RECT 482.350 1139.490 482.730 1139.500 ;
        RECT 497.110 1139.490 497.410 1140.550 ;
        RECT 531.110 1140.540 531.490 1140.550 ;
        RECT 676.510 1140.550 700.515 1140.850 ;
        RECT 593.925 1140.170 594.255 1140.185 ;
        RECT 627.710 1140.170 628.090 1140.180 ;
        RECT 593.925 1139.870 628.090 1140.170 ;
        RECT 593.925 1139.855 594.255 1139.870 ;
        RECT 627.710 1139.860 628.090 1139.870 ;
        RECT 482.350 1139.190 497.410 1139.490 ;
        RECT 675.805 1139.490 676.135 1139.505 ;
        RECT 676.510 1139.490 676.810 1140.550 ;
        RECT 700.185 1140.535 700.515 1140.550 ;
        RECT 772.405 1140.170 772.735 1140.185 ;
        RECT 772.405 1139.870 807.450 1140.170 ;
        RECT 772.405 1139.855 772.735 1139.870 ;
        RECT 737.905 1139.490 738.235 1139.505 ;
        RECT 675.805 1139.190 676.810 1139.490 ;
        RECT 724.350 1139.190 738.235 1139.490 ;
        RECT 807.150 1139.490 807.450 1139.870 ;
        RECT 855.910 1139.870 904.050 1140.170 ;
        RECT 807.150 1139.190 855.290 1139.490 ;
        RECT 482.350 1139.180 482.730 1139.190 ;
        RECT 675.805 1139.175 676.135 1139.190 ;
        RECT 434.510 1138.810 434.890 1138.820 ;
        RECT 410.630 1138.510 434.890 1138.810 ;
        RECT 434.510 1138.500 434.890 1138.510 ;
        RECT 555.285 1138.810 555.615 1138.825 ;
        RECT 579.665 1138.810 579.995 1138.825 ;
        RECT 555.285 1138.510 579.995 1138.810 ;
        RECT 555.285 1138.495 555.615 1138.510 ;
        RECT 579.665 1138.495 579.995 1138.510 ;
        RECT 700.185 1138.810 700.515 1138.825 ;
        RECT 724.350 1138.810 724.650 1139.190 ;
        RECT 737.905 1139.175 738.235 1139.190 ;
        RECT 700.185 1138.510 724.650 1138.810 ;
        RECT 854.990 1138.810 855.290 1139.190 ;
        RECT 855.910 1138.810 856.210 1139.870 ;
        RECT 903.750 1139.490 904.050 1139.870 ;
        RECT 952.510 1139.870 1000.650 1140.170 ;
        RECT 903.750 1139.190 951.890 1139.490 ;
        RECT 854.990 1138.510 856.210 1138.810 ;
        RECT 951.590 1138.810 951.890 1139.190 ;
        RECT 952.510 1138.810 952.810 1139.870 ;
        RECT 1000.350 1139.490 1000.650 1139.870 ;
        RECT 1049.110 1139.870 1097.250 1140.170 ;
        RECT 1000.350 1139.190 1048.490 1139.490 ;
        RECT 951.590 1138.510 952.810 1138.810 ;
        RECT 1048.190 1138.810 1048.490 1139.190 ;
        RECT 1049.110 1138.810 1049.410 1139.870 ;
        RECT 1096.950 1139.490 1097.250 1139.870 ;
        RECT 1145.710 1139.870 1193.850 1140.170 ;
        RECT 1096.950 1139.190 1145.090 1139.490 ;
        RECT 1048.190 1138.510 1049.410 1138.810 ;
        RECT 1144.790 1138.810 1145.090 1139.190 ;
        RECT 1145.710 1138.810 1146.010 1139.870 ;
        RECT 1193.550 1139.490 1193.850 1139.870 ;
        RECT 1242.310 1139.870 1290.450 1140.170 ;
        RECT 1193.550 1139.190 1241.690 1139.490 ;
        RECT 1144.790 1138.510 1146.010 1138.810 ;
        RECT 1241.390 1138.810 1241.690 1139.190 ;
        RECT 1242.310 1138.810 1242.610 1139.870 ;
        RECT 1290.150 1139.490 1290.450 1139.870 ;
        RECT 1338.910 1139.870 1387.050 1140.170 ;
        RECT 1290.150 1139.190 1338.290 1139.490 ;
        RECT 1241.390 1138.510 1242.610 1138.810 ;
        RECT 1337.990 1138.810 1338.290 1139.190 ;
        RECT 1338.910 1138.810 1339.210 1139.870 ;
        RECT 1386.750 1139.490 1387.050 1139.870 ;
        RECT 1435.510 1139.870 1483.650 1140.170 ;
        RECT 1386.750 1139.190 1434.890 1139.490 ;
        RECT 1337.990 1138.510 1339.210 1138.810 ;
        RECT 1434.590 1138.810 1434.890 1139.190 ;
        RECT 1435.510 1138.810 1435.810 1139.870 ;
        RECT 1483.350 1139.490 1483.650 1139.870 ;
        RECT 1532.110 1139.870 1580.250 1140.170 ;
        RECT 1483.350 1139.190 1531.490 1139.490 ;
        RECT 1434.590 1138.510 1435.810 1138.810 ;
        RECT 1531.190 1138.810 1531.490 1139.190 ;
        RECT 1532.110 1138.810 1532.410 1139.870 ;
        RECT 1579.950 1139.490 1580.250 1139.870 ;
        RECT 1628.710 1139.870 1676.850 1140.170 ;
        RECT 1579.950 1139.190 1628.090 1139.490 ;
        RECT 1531.190 1138.510 1532.410 1138.810 ;
        RECT 1627.790 1138.810 1628.090 1139.190 ;
        RECT 1628.710 1138.810 1629.010 1139.870 ;
        RECT 1676.550 1139.490 1676.850 1139.870 ;
        RECT 1725.310 1139.870 1773.450 1140.170 ;
        RECT 1676.550 1139.190 1724.690 1139.490 ;
        RECT 1627.790 1138.510 1629.010 1138.810 ;
        RECT 1724.390 1138.810 1724.690 1139.190 ;
        RECT 1725.310 1138.810 1725.610 1139.870 ;
        RECT 1773.150 1139.490 1773.450 1139.870 ;
        RECT 1821.910 1139.870 1870.050 1140.170 ;
        RECT 1773.150 1139.190 1821.290 1139.490 ;
        RECT 1724.390 1138.510 1725.610 1138.810 ;
        RECT 1820.990 1138.810 1821.290 1139.190 ;
        RECT 1821.910 1138.810 1822.210 1139.870 ;
        RECT 1869.750 1139.490 1870.050 1139.870 ;
        RECT 1918.510 1139.870 1966.650 1140.170 ;
        RECT 1869.750 1139.190 1917.890 1139.490 ;
        RECT 1820.990 1138.510 1822.210 1138.810 ;
        RECT 1917.590 1138.810 1917.890 1139.190 ;
        RECT 1918.510 1138.810 1918.810 1139.870 ;
        RECT 1966.350 1139.490 1966.650 1139.870 ;
        RECT 2015.110 1139.870 2063.250 1140.170 ;
        RECT 1966.350 1139.190 2014.490 1139.490 ;
        RECT 1917.590 1138.510 1918.810 1138.810 ;
        RECT 2014.190 1138.810 2014.490 1139.190 ;
        RECT 2015.110 1138.810 2015.410 1139.870 ;
        RECT 2062.950 1139.490 2063.250 1139.870 ;
        RECT 2111.710 1139.870 2159.850 1140.170 ;
        RECT 2062.950 1139.190 2111.090 1139.490 ;
        RECT 2014.190 1138.510 2015.410 1138.810 ;
        RECT 2110.790 1138.810 2111.090 1139.190 ;
        RECT 2111.710 1138.810 2112.010 1139.870 ;
        RECT 2159.550 1139.490 2159.850 1139.870 ;
        RECT 2208.310 1139.870 2256.450 1140.170 ;
        RECT 2159.550 1139.190 2207.690 1139.490 ;
        RECT 2110.790 1138.510 2112.010 1138.810 ;
        RECT 2207.390 1138.810 2207.690 1139.190 ;
        RECT 2208.310 1138.810 2208.610 1139.870 ;
        RECT 2256.150 1139.490 2256.450 1139.870 ;
        RECT 2304.910 1139.870 2353.050 1140.170 ;
        RECT 2256.150 1139.190 2304.290 1139.490 ;
        RECT 2207.390 1138.510 2208.610 1138.810 ;
        RECT 2303.990 1138.810 2304.290 1139.190 ;
        RECT 2304.910 1138.810 2305.210 1139.870 ;
        RECT 2352.750 1139.490 2353.050 1139.870 ;
        RECT 2401.510 1139.870 2449.650 1140.170 ;
        RECT 2352.750 1139.190 2400.890 1139.490 ;
        RECT 2303.990 1138.510 2305.210 1138.810 ;
        RECT 2400.590 1138.810 2400.890 1139.190 ;
        RECT 2401.510 1138.810 2401.810 1139.870 ;
        RECT 2449.350 1139.490 2449.650 1139.870 ;
        RECT 2498.110 1139.870 2546.250 1140.170 ;
        RECT 2449.350 1139.190 2497.490 1139.490 ;
        RECT 2400.590 1138.510 2401.810 1138.810 ;
        RECT 2497.190 1138.810 2497.490 1139.190 ;
        RECT 2498.110 1138.810 2498.410 1139.870 ;
        RECT 2545.950 1139.490 2546.250 1139.870 ;
        RECT 2594.710 1139.870 2642.850 1140.170 ;
        RECT 2545.950 1139.190 2594.090 1139.490 ;
        RECT 2497.190 1138.510 2498.410 1138.810 ;
        RECT 2593.790 1138.810 2594.090 1139.190 ;
        RECT 2594.710 1138.810 2595.010 1139.870 ;
        RECT 2642.550 1139.490 2642.850 1139.870 ;
        RECT 2691.310 1139.870 2739.450 1140.170 ;
        RECT 2642.550 1139.190 2690.690 1139.490 ;
        RECT 2593.790 1138.510 2595.010 1138.810 ;
        RECT 2690.390 1138.810 2690.690 1139.190 ;
        RECT 2691.310 1138.810 2691.610 1139.870 ;
        RECT 2739.150 1139.490 2739.450 1139.870 ;
        RECT 2787.910 1139.870 2836.050 1140.170 ;
        RECT 2739.150 1139.190 2787.290 1139.490 ;
        RECT 2690.390 1138.510 2691.610 1138.810 ;
        RECT 2786.990 1138.810 2787.290 1139.190 ;
        RECT 2787.910 1138.810 2788.210 1139.870 ;
        RECT 2835.750 1139.490 2836.050 1139.870 ;
        RECT 2916.710 1139.490 2917.010 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 2835.750 1139.190 2883.890 1139.490 ;
        RECT 2786.990 1138.510 2788.210 1138.810 ;
        RECT 2883.590 1138.810 2883.890 1139.190 ;
        RECT 2884.510 1139.190 2917.010 1139.490 ;
        RECT 2884.510 1138.810 2884.810 1139.190 ;
        RECT 2883.590 1138.510 2884.810 1138.810 ;
        RECT 700.185 1138.495 700.515 1138.510 ;
        RECT 434.510 1137.450 434.890 1137.460 ;
        RECT 482.350 1137.450 482.730 1137.460 ;
        RECT 434.510 1137.150 482.730 1137.450 ;
        RECT 434.510 1137.140 434.890 1137.150 ;
        RECT 482.350 1137.140 482.730 1137.150 ;
      LAYER via3 ;
        RECT 285.500 1730.100 285.820 1730.420 ;
        RECT 531.140 1141.900 531.460 1142.220 ;
        RECT 627.740 1141.220 628.060 1141.540 ;
        RECT 285.500 1139.860 285.820 1140.180 ;
        RECT 482.380 1139.180 482.700 1139.500 ;
        RECT 531.140 1140.540 531.460 1140.860 ;
        RECT 627.740 1139.860 628.060 1140.180 ;
        RECT 434.540 1138.500 434.860 1138.820 ;
        RECT 434.540 1137.140 434.860 1137.460 ;
        RECT 482.380 1137.140 482.700 1137.460 ;
      LAYER met4 ;
        RECT 285.495 1730.095 285.825 1730.425 ;
        RECT 285.510 1140.185 285.810 1730.095 ;
        RECT 531.135 1141.895 531.465 1142.225 ;
        RECT 531.150 1140.865 531.450 1141.895 ;
        RECT 627.735 1141.215 628.065 1141.545 ;
        RECT 531.135 1140.535 531.465 1140.865 ;
        RECT 627.750 1140.185 628.050 1141.215 ;
        RECT 285.495 1139.855 285.825 1140.185 ;
        RECT 627.735 1139.855 628.065 1140.185 ;
        RECT 482.375 1139.175 482.705 1139.505 ;
        RECT 434.535 1138.495 434.865 1138.825 ;
        RECT 434.550 1137.465 434.850 1138.495 ;
        RECT 482.390 1137.465 482.690 1139.175 ;
        RECT 434.535 1137.135 434.865 1137.465 ;
        RECT 482.375 1137.135 482.705 1137.465 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.730 1379.960 286.050 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 285.730 1379.820 2901.150 1379.960 ;
        RECT 285.730 1379.760 286.050 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 285.760 1379.760 286.020 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 285.750 1759.315 286.030 1759.685 ;
        RECT 285.820 1380.050 285.960 1759.315 ;
        RECT 285.760 1379.730 286.020 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 285.750 1759.360 286.030 1759.640 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 285.725 1759.650 286.055 1759.665 ;
        RECT 300.000 1759.650 304.000 1759.760 ;
        RECT 285.725 1759.350 304.000 1759.650 ;
        RECT 285.725 1759.335 286.055 1759.350 ;
        RECT 300.000 1759.160 304.000 1759.350 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 282.970 1654.000 283.290 1654.060 ;
        RECT 282.970 1653.860 285.500 1654.000 ;
        RECT 282.970 1653.800 283.290 1653.860 ;
        RECT 285.360 1652.360 285.500 1653.860 ;
        RECT 285.270 1652.100 285.590 1652.360 ;
        RECT 285.270 1646.180 285.590 1646.240 ;
        RECT 288.950 1646.180 289.270 1646.240 ;
        RECT 285.270 1646.040 289.270 1646.180 ;
        RECT 285.270 1645.980 285.590 1646.040 ;
        RECT 288.950 1645.980 289.270 1646.040 ;
        RECT 288.030 1603.000 288.350 1603.060 ;
        RECT 1400.310 1603.000 1400.630 1603.060 ;
        RECT 288.030 1602.860 1400.630 1603.000 ;
        RECT 288.030 1602.800 288.350 1602.860 ;
        RECT 1400.310 1602.800 1400.630 1602.860 ;
      LAYER via ;
        RECT 283.000 1653.800 283.260 1654.060 ;
        RECT 285.300 1652.100 285.560 1652.360 ;
        RECT 285.300 1645.980 285.560 1646.240 ;
        RECT 288.980 1645.980 289.240 1646.240 ;
        RECT 288.060 1602.800 288.320 1603.060 ;
        RECT 1400.340 1602.800 1400.600 1603.060 ;
      LAYER met2 ;
        RECT 282.990 1787.875 283.270 1788.245 ;
        RECT 283.060 1654.090 283.200 1787.875 ;
        RECT 283.000 1653.770 283.260 1654.090 ;
        RECT 285.300 1652.070 285.560 1652.390 ;
        RECT 285.360 1646.270 285.500 1652.070 ;
        RECT 285.300 1645.950 285.560 1646.270 ;
        RECT 288.980 1645.950 289.240 1646.270 ;
        RECT 289.040 1624.930 289.180 1645.950 ;
        RECT 288.120 1624.790 289.180 1624.930 ;
        RECT 288.120 1603.090 288.260 1624.790 ;
        RECT 2899.930 1613.115 2900.210 1613.485 ;
        RECT 2900.000 1603.285 2900.140 1613.115 ;
        RECT 288.060 1602.770 288.320 1603.090 ;
        RECT 1400.330 1602.915 1400.610 1603.285 ;
        RECT 1698.870 1602.915 1699.150 1603.285 ;
        RECT 1749.930 1602.915 1750.210 1603.285 ;
        RECT 2899.930 1602.915 2900.210 1603.285 ;
        RECT 1400.340 1602.770 1400.600 1602.915 ;
        RECT 1698.940 1601.925 1699.080 1602.915 ;
        RECT 1750.000 1601.925 1750.140 1602.915 ;
        RECT 1698.870 1601.555 1699.150 1601.925 ;
        RECT 1749.930 1601.555 1750.210 1601.925 ;
      LAYER via2 ;
        RECT 282.990 1787.920 283.270 1788.200 ;
        RECT 2899.930 1613.160 2900.210 1613.440 ;
        RECT 1400.330 1602.960 1400.610 1603.240 ;
        RECT 1698.870 1602.960 1699.150 1603.240 ;
        RECT 1749.930 1602.960 1750.210 1603.240 ;
        RECT 2899.930 1602.960 2900.210 1603.240 ;
        RECT 1698.870 1601.600 1699.150 1601.880 ;
        RECT 1749.930 1601.600 1750.210 1601.880 ;
      LAYER met3 ;
        RECT 282.965 1788.210 283.295 1788.225 ;
        RECT 300.000 1788.210 304.000 1788.320 ;
        RECT 282.965 1787.910 304.000 1788.210 ;
        RECT 282.965 1787.895 283.295 1787.910 ;
        RECT 300.000 1787.720 304.000 1787.910 ;
        RECT 2899.905 1613.450 2900.235 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2899.905 1613.150 2924.800 1613.450 ;
        RECT 2899.905 1613.135 2900.235 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 1400.305 1603.250 1400.635 1603.265 ;
        RECT 1698.845 1603.250 1699.175 1603.265 ;
        RECT 1400.305 1602.950 1699.175 1603.250 ;
        RECT 1400.305 1602.935 1400.635 1602.950 ;
        RECT 1698.845 1602.935 1699.175 1602.950 ;
        RECT 1749.905 1603.250 1750.235 1603.265 ;
        RECT 2899.905 1603.250 2900.235 1603.265 ;
        RECT 1749.905 1602.950 2900.235 1603.250 ;
        RECT 1749.905 1602.935 1750.235 1602.950 ;
        RECT 2899.905 1602.935 2900.235 1602.950 ;
        RECT 1698.845 1601.890 1699.175 1601.905 ;
        RECT 1749.905 1601.890 1750.235 1601.905 ;
        RECT 1698.845 1601.590 1750.235 1601.890 ;
        RECT 1698.845 1601.575 1699.175 1601.590 ;
        RECT 1749.905 1601.575 1750.235 1601.590 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.350 1626.120 284.670 1626.180 ;
        RECT 287.570 1626.120 287.890 1626.180 ;
        RECT 284.350 1625.980 287.890 1626.120 ;
        RECT 284.350 1625.920 284.670 1625.980 ;
        RECT 287.570 1625.920 287.890 1625.980 ;
        RECT 284.350 1600.620 284.670 1600.680 ;
        RECT 2904.050 1600.620 2904.370 1600.680 ;
        RECT 284.350 1600.480 2904.370 1600.620 ;
        RECT 284.350 1600.420 284.670 1600.480 ;
        RECT 2904.050 1600.420 2904.370 1600.480 ;
      LAYER via ;
        RECT 284.380 1625.920 284.640 1626.180 ;
        RECT 287.600 1625.920 287.860 1626.180 ;
        RECT 284.380 1600.420 284.640 1600.680 ;
        RECT 2904.080 1600.420 2904.340 1600.680 ;
      LAYER met2 ;
        RECT 2904.070 1847.715 2904.350 1848.085 ;
        RECT 287.590 1817.115 287.870 1817.485 ;
        RECT 287.660 1626.210 287.800 1817.115 ;
        RECT 284.380 1625.890 284.640 1626.210 ;
        RECT 287.600 1625.890 287.860 1626.210 ;
        RECT 284.440 1600.710 284.580 1625.890 ;
        RECT 2904.140 1600.710 2904.280 1847.715 ;
        RECT 284.380 1600.390 284.640 1600.710 ;
        RECT 2904.080 1600.390 2904.340 1600.710 ;
      LAYER via2 ;
        RECT 2904.070 1847.760 2904.350 1848.040 ;
        RECT 287.590 1817.160 287.870 1817.440 ;
      LAYER met3 ;
        RECT 2904.045 1848.050 2904.375 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2904.045 1847.750 2924.800 1848.050 ;
        RECT 2904.045 1847.735 2904.375 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 287.565 1817.450 287.895 1817.465 ;
        RECT 300.000 1817.450 304.000 1817.560 ;
        RECT 287.565 1817.150 304.000 1817.450 ;
        RECT 287.565 1817.135 287.895 1817.150 ;
        RECT 300.000 1816.960 304.000 1817.150 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1625.780 289.730 1625.840 ;
        RECT 297.690 1625.780 298.010 1625.840 ;
        RECT 289.410 1625.640 298.010 1625.780 ;
        RECT 289.410 1625.580 289.730 1625.640 ;
        RECT 297.690 1625.580 298.010 1625.640 ;
        RECT 297.690 1602.660 298.010 1602.720 ;
        RECT 1399.850 1602.660 1400.170 1602.720 ;
        RECT 297.690 1602.520 1400.170 1602.660 ;
        RECT 297.690 1602.460 298.010 1602.520 ;
        RECT 1399.850 1602.460 1400.170 1602.520 ;
      LAYER via ;
        RECT 289.440 1625.580 289.700 1625.840 ;
        RECT 297.720 1625.580 297.980 1625.840 ;
        RECT 297.720 1602.460 297.980 1602.720 ;
        RECT 1399.880 1602.460 1400.140 1602.720 ;
      LAYER met2 ;
        RECT 2902.690 2082.315 2902.970 2082.685 ;
        RECT 289.430 1845.675 289.710 1846.045 ;
        RECT 289.500 1625.870 289.640 1845.675 ;
        RECT 289.440 1625.550 289.700 1625.870 ;
        RECT 297.720 1625.550 297.980 1625.870 ;
        RECT 297.780 1602.750 297.920 1625.550 ;
        RECT 2902.760 1604.645 2902.900 2082.315 ;
        RECT 1399.870 1604.275 1400.150 1604.645 ;
        RECT 2902.690 1604.275 2902.970 1604.645 ;
        RECT 1399.940 1602.750 1400.080 1604.275 ;
        RECT 297.720 1602.430 297.980 1602.750 ;
        RECT 1399.880 1602.430 1400.140 1602.750 ;
      LAYER via2 ;
        RECT 2902.690 2082.360 2902.970 2082.640 ;
        RECT 289.430 1845.720 289.710 1846.000 ;
        RECT 1399.870 1604.320 1400.150 1604.600 ;
        RECT 2902.690 1604.320 2902.970 1604.600 ;
      LAYER met3 ;
        RECT 2902.665 2082.650 2902.995 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2902.665 2082.350 2924.800 2082.650 ;
        RECT 2902.665 2082.335 2902.995 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 289.405 1846.010 289.735 1846.025 ;
        RECT 300.000 1846.010 304.000 1846.120 ;
        RECT 289.405 1845.710 304.000 1846.010 ;
        RECT 289.405 1845.695 289.735 1845.710 ;
        RECT 300.000 1845.520 304.000 1845.710 ;
        RECT 1399.845 1604.610 1400.175 1604.625 ;
        RECT 2902.665 1604.610 2902.995 1604.625 ;
        RECT 1399.845 1604.310 1699.850 1604.610 ;
        RECT 1399.845 1604.295 1400.175 1604.310 ;
        RECT 1699.550 1603.250 1699.850 1604.310 ;
        RECT 1748.310 1604.310 2902.995 1604.610 ;
        RECT 1748.310 1603.250 1748.610 1604.310 ;
        RECT 2902.665 1604.295 2902.995 1604.310 ;
        RECT 1699.550 1602.950 1748.610 1603.250 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 298.610 1602.320 298.930 1602.380 ;
        RECT 1400.310 1602.320 1400.630 1602.380 ;
        RECT 298.610 1602.180 1400.630 1602.320 ;
        RECT 298.610 1602.120 298.930 1602.180 ;
        RECT 1400.310 1602.120 1400.630 1602.180 ;
      LAYER via ;
        RECT 298.640 1602.120 298.900 1602.380 ;
        RECT 1400.340 1602.120 1400.600 1602.380 ;
      LAYER met2 ;
        RECT 2901.310 2316.915 2901.590 2317.285 ;
        RECT 298.630 1653.235 298.910 1653.605 ;
        RECT 298.700 1602.410 298.840 1653.235 ;
        RECT 2901.380 1602.605 2901.520 2316.915 ;
        RECT 298.640 1602.090 298.900 1602.410 ;
        RECT 1400.330 1602.235 1400.610 1602.605 ;
        RECT 2901.310 1602.235 2901.590 1602.605 ;
        RECT 1400.340 1602.090 1400.600 1602.235 ;
      LAYER via2 ;
        RECT 2901.310 2316.960 2901.590 2317.240 ;
        RECT 298.630 1653.280 298.910 1653.560 ;
        RECT 1400.330 1602.280 1400.610 1602.560 ;
        RECT 2901.310 1602.280 2901.590 1602.560 ;
      LAYER met3 ;
        RECT 2901.285 2317.250 2901.615 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2901.285 2316.950 2924.800 2317.250 ;
        RECT 2901.285 2316.935 2901.615 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 289.150 1875.250 289.530 1875.260 ;
        RECT 300.000 1875.250 304.000 1875.360 ;
        RECT 289.150 1874.950 304.000 1875.250 ;
        RECT 289.150 1874.940 289.530 1874.950 ;
        RECT 300.000 1874.760 304.000 1874.950 ;
        RECT 289.150 1653.570 289.530 1653.580 ;
        RECT 298.605 1653.570 298.935 1653.585 ;
        RECT 289.150 1653.270 298.935 1653.570 ;
        RECT 289.150 1653.260 289.530 1653.270 ;
        RECT 298.605 1653.255 298.935 1653.270 ;
        RECT 1400.305 1602.570 1400.635 1602.585 ;
        RECT 2901.285 1602.570 2901.615 1602.585 ;
        RECT 1400.305 1602.270 2901.615 1602.570 ;
        RECT 1400.305 1602.255 1400.635 1602.270 ;
        RECT 2901.285 1602.255 2901.615 1602.270 ;
      LAYER via3 ;
        RECT 289.180 1874.940 289.500 1875.260 ;
        RECT 289.180 1653.260 289.500 1653.580 ;
      LAYER met4 ;
        RECT 289.175 1874.935 289.505 1875.265 ;
        RECT 289.190 1653.585 289.490 1874.935 ;
        RECT 289.175 1653.255 289.505 1653.585 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 151.540 289.270 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 288.950 151.400 2901.150 151.540 ;
        RECT 288.950 151.340 289.270 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 288.980 151.340 289.240 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 288.970 1623.995 289.250 1624.365 ;
        RECT 289.040 151.630 289.180 1623.995 ;
        RECT 288.980 151.310 289.240 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 288.970 1624.040 289.250 1624.320 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 288.945 1624.330 289.275 1624.345 ;
        RECT 300.000 1624.330 304.000 1624.440 ;
        RECT 288.945 1624.030 304.000 1624.330 ;
        RECT 288.945 1624.015 289.275 1624.030 ;
        RECT 300.000 1623.840 304.000 1624.030 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 285.730 2696.100 286.050 2696.160 ;
        RECT 2901.290 2696.100 2901.610 2696.160 ;
        RECT 285.730 2695.960 2901.610 2696.100 ;
        RECT 285.730 2695.900 286.050 2695.960 ;
        RECT 2901.290 2695.900 2901.610 2695.960 ;
      LAYER via ;
        RECT 285.760 2695.900 286.020 2696.160 ;
        RECT 2901.320 2695.900 2901.580 2696.160 ;
      LAYER met2 ;
        RECT 285.760 2695.870 286.020 2696.190 ;
        RECT 2901.320 2695.870 2901.580 2696.190 ;
        RECT 285.820 1914.045 285.960 2695.870 ;
        RECT 2901.380 2493.405 2901.520 2695.870 ;
        RECT 2901.310 2493.035 2901.590 2493.405 ;
        RECT 285.750 1913.675 286.030 1914.045 ;
      LAYER via2 ;
        RECT 2901.310 2493.080 2901.590 2493.360 ;
        RECT 285.750 1913.720 286.030 1914.000 ;
      LAYER met3 ;
        RECT 2901.285 2493.370 2901.615 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2901.285 2493.070 2924.800 2493.370 ;
        RECT 2901.285 2493.055 2901.615 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 285.725 1914.010 286.055 1914.025 ;
        RECT 300.000 1914.010 304.000 1914.120 ;
        RECT 285.725 1913.710 304.000 1914.010 ;
        RECT 285.725 1913.695 286.055 1913.710 ;
        RECT 300.000 1913.520 304.000 1913.710 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2801.470 2727.720 2801.790 2727.780 ;
        RECT 2815.730 2727.720 2816.050 2727.780 ;
        RECT 2801.470 2727.580 2816.050 2727.720 ;
        RECT 2801.470 2727.520 2801.790 2727.580 ;
        RECT 2815.730 2727.520 2816.050 2727.580 ;
        RECT 1510.710 2727.380 1511.030 2727.440 ;
        RECT 1545.210 2727.380 1545.530 2727.440 ;
        RECT 1510.710 2727.240 1545.530 2727.380 ;
        RECT 1510.710 2727.180 1511.030 2727.240 ;
        RECT 1545.210 2727.180 1545.530 2727.240 ;
        RECT 2863.110 2727.380 2863.430 2727.440 ;
        RECT 2897.610 2727.380 2897.930 2727.440 ;
        RECT 2863.110 2727.240 2897.930 2727.380 ;
        RECT 2863.110 2727.180 2863.430 2727.240 ;
        RECT 2897.610 2727.180 2897.930 2727.240 ;
        RECT 579.670 2727.040 579.990 2727.100 ;
        RECT 627.050 2727.040 627.370 2727.100 ;
        RECT 579.670 2726.900 627.370 2727.040 ;
        RECT 579.670 2726.840 579.990 2726.900 ;
        RECT 627.050 2726.840 627.370 2726.900 ;
        RECT 676.270 2727.040 676.590 2727.100 ;
        RECT 724.110 2727.040 724.430 2727.100 ;
        RECT 676.270 2726.900 724.430 2727.040 ;
        RECT 676.270 2726.840 676.590 2726.900 ;
        RECT 724.110 2726.840 724.430 2726.900 ;
        RECT 979.410 2727.040 979.730 2727.100 ;
        RECT 1007.010 2727.040 1007.330 2727.100 ;
        RECT 979.410 2726.900 1007.330 2727.040 ;
        RECT 979.410 2726.840 979.730 2726.900 ;
        RECT 1007.010 2726.840 1007.330 2726.900 ;
        RECT 1062.670 2727.040 1062.990 2727.100 ;
        RECT 1110.050 2727.040 1110.370 2727.100 ;
        RECT 1062.670 2726.900 1110.370 2727.040 ;
        RECT 1062.670 2726.840 1062.990 2726.900 ;
        RECT 1110.050 2726.840 1110.370 2726.900 ;
        RECT 1159.270 2727.040 1159.590 2727.100 ;
        RECT 1207.110 2727.040 1207.430 2727.100 ;
        RECT 1159.270 2726.900 1207.430 2727.040 ;
        RECT 1159.270 2726.840 1159.590 2726.900 ;
        RECT 1207.110 2726.840 1207.430 2726.900 ;
        RECT 1255.870 2727.040 1256.190 2727.100 ;
        RECT 1303.710 2727.040 1304.030 2727.100 ;
        RECT 1255.870 2726.900 1304.030 2727.040 ;
        RECT 1255.870 2726.840 1256.190 2726.900 ;
        RECT 1303.710 2726.840 1304.030 2726.900 ;
        RECT 2415.070 2727.040 2415.390 2727.100 ;
        RECT 2429.330 2727.040 2429.650 2727.100 ;
        RECT 2415.070 2726.900 2429.650 2727.040 ;
        RECT 2415.070 2726.840 2415.390 2726.900 ;
        RECT 2429.330 2726.840 2429.650 2726.900 ;
        RECT 2704.870 2727.040 2705.190 2727.100 ;
        RECT 2743.050 2727.040 2743.370 2727.100 ;
        RECT 2704.870 2726.900 2743.370 2727.040 ;
        RECT 2704.870 2726.840 2705.190 2726.900 ;
        RECT 2743.050 2726.840 2743.370 2726.900 ;
        RECT 427.870 2726.700 428.190 2726.760 ;
        RECT 475.250 2726.700 475.570 2726.760 ;
        RECT 427.870 2726.560 475.570 2726.700 ;
        RECT 427.870 2726.500 428.190 2726.560 ;
        RECT 475.250 2726.500 475.570 2726.560 ;
        RECT 834.510 2726.700 834.830 2726.760 ;
        RECT 886.490 2726.700 886.810 2726.760 ;
        RECT 834.510 2726.560 886.810 2726.700 ;
        RECT 834.510 2726.500 834.830 2726.560 ;
        RECT 886.490 2726.500 886.810 2726.560 ;
        RECT 1607.310 2726.700 1607.630 2726.760 ;
        RECT 1641.810 2726.700 1642.130 2726.760 ;
        RECT 1607.310 2726.560 1642.130 2726.700 ;
        RECT 1607.310 2726.500 1607.630 2726.560 ;
        RECT 1641.810 2726.500 1642.130 2726.560 ;
        RECT 483.070 2726.360 483.390 2726.420 ;
        RECT 524.010 2726.360 524.330 2726.420 ;
        RECT 483.070 2726.220 524.330 2726.360 ;
        RECT 483.070 2726.160 483.390 2726.220 ;
        RECT 524.010 2726.160 524.330 2726.220 ;
      LAYER via ;
        RECT 2801.500 2727.520 2801.760 2727.780 ;
        RECT 2815.760 2727.520 2816.020 2727.780 ;
        RECT 1510.740 2727.180 1511.000 2727.440 ;
        RECT 1545.240 2727.180 1545.500 2727.440 ;
        RECT 2863.140 2727.180 2863.400 2727.440 ;
        RECT 2897.640 2727.180 2897.900 2727.440 ;
        RECT 579.700 2726.840 579.960 2727.100 ;
        RECT 627.080 2726.840 627.340 2727.100 ;
        RECT 676.300 2726.840 676.560 2727.100 ;
        RECT 724.140 2726.840 724.400 2727.100 ;
        RECT 979.440 2726.840 979.700 2727.100 ;
        RECT 1007.040 2726.840 1007.300 2727.100 ;
        RECT 1062.700 2726.840 1062.960 2727.100 ;
        RECT 1110.080 2726.840 1110.340 2727.100 ;
        RECT 1159.300 2726.840 1159.560 2727.100 ;
        RECT 1207.140 2726.840 1207.400 2727.100 ;
        RECT 1255.900 2726.840 1256.160 2727.100 ;
        RECT 1303.740 2726.840 1304.000 2727.100 ;
        RECT 2415.100 2726.840 2415.360 2727.100 ;
        RECT 2429.360 2726.840 2429.620 2727.100 ;
        RECT 2704.900 2726.840 2705.160 2727.100 ;
        RECT 2743.080 2726.840 2743.340 2727.100 ;
        RECT 427.900 2726.500 428.160 2726.760 ;
        RECT 475.280 2726.500 475.540 2726.760 ;
        RECT 834.540 2726.500 834.800 2726.760 ;
        RECT 886.520 2726.500 886.780 2726.760 ;
        RECT 1607.340 2726.500 1607.600 2726.760 ;
        RECT 1641.840 2726.500 1642.100 2726.760 ;
        RECT 483.100 2726.160 483.360 2726.420 ;
        RECT 524.040 2726.160 524.300 2726.420 ;
      LAYER met2 ;
        RECT 1037.850 2728.315 1038.130 2728.685 ;
        RECT 1037.920 2727.325 1038.060 2728.315 ;
        RECT 1545.230 2727.635 1545.510 2728.005 ;
        RECT 1859.410 2727.635 1859.690 2728.005 ;
        RECT 2766.530 2727.890 2766.810 2728.005 ;
        RECT 2767.450 2727.890 2767.730 2728.005 ;
        RECT 2766.530 2727.750 2767.730 2727.890 ;
        RECT 2766.530 2727.635 2766.810 2727.750 ;
        RECT 2767.450 2727.635 2767.730 2727.750 ;
        RECT 2801.490 2727.635 2801.770 2728.005 ;
        RECT 1545.300 2727.470 1545.440 2727.635 ;
        RECT 1510.740 2727.325 1511.000 2727.470 ;
        RECT 579.690 2726.955 579.970 2727.325 ;
        RECT 579.700 2726.810 579.960 2726.955 ;
        RECT 627.080 2726.810 627.340 2727.130 ;
        RECT 676.290 2726.955 676.570 2727.325 ;
        RECT 676.300 2726.810 676.560 2726.955 ;
        RECT 724.140 2726.810 724.400 2727.130 ;
        RECT 979.430 2726.955 979.710 2727.325 ;
        RECT 1007.030 2726.955 1007.310 2727.325 ;
        RECT 1037.850 2726.955 1038.130 2727.325 ;
        RECT 1062.690 2726.955 1062.970 2727.325 ;
        RECT 979.440 2726.810 979.700 2726.955 ;
        RECT 1007.040 2726.810 1007.300 2726.955 ;
        RECT 1062.700 2726.810 1062.960 2726.955 ;
        RECT 1110.080 2726.810 1110.340 2727.130 ;
        RECT 1159.290 2726.955 1159.570 2727.325 ;
        RECT 1159.300 2726.810 1159.560 2726.955 ;
        RECT 1207.140 2726.810 1207.400 2727.130 ;
        RECT 1255.890 2726.955 1256.170 2727.325 ;
        RECT 1255.900 2726.810 1256.160 2726.955 ;
        RECT 1303.740 2726.810 1304.000 2727.130 ;
        RECT 1510.730 2726.955 1511.010 2727.325 ;
        RECT 1545.240 2727.150 1545.500 2727.470 ;
        RECT 1641.830 2726.955 1642.110 2727.325 ;
        RECT 1738.430 2726.955 1738.710 2727.325 ;
        RECT 427.900 2726.645 428.160 2726.790 ;
        RECT 475.280 2726.645 475.540 2726.790 ;
        RECT 427.890 2726.275 428.170 2726.645 ;
        RECT 475.270 2726.275 475.550 2726.645 ;
        RECT 483.090 2726.275 483.370 2726.645 ;
        RECT 483.100 2726.130 483.360 2726.275 ;
        RECT 524.040 2726.130 524.300 2726.450 ;
        RECT 524.100 2725.965 524.240 2726.130 ;
        RECT 627.140 2725.965 627.280 2726.810 ;
        RECT 724.200 2725.965 724.340 2726.810 ;
        RECT 834.540 2726.645 834.800 2726.790 ;
        RECT 886.520 2726.645 886.780 2726.790 ;
        RECT 834.530 2726.275 834.810 2726.645 ;
        RECT 886.510 2726.275 886.790 2726.645 ;
        RECT 1110.140 2725.965 1110.280 2726.810 ;
        RECT 1207.200 2725.965 1207.340 2726.810 ;
        RECT 1303.800 2725.965 1303.940 2726.810 ;
        RECT 1641.900 2726.790 1642.040 2726.955 ;
        RECT 1607.340 2726.645 1607.600 2726.790 ;
        RECT 1607.330 2726.275 1607.610 2726.645 ;
        RECT 1641.840 2726.470 1642.100 2726.790 ;
        RECT 1738.500 2726.645 1738.640 2726.955 ;
        RECT 1738.430 2726.275 1738.710 2726.645 ;
        RECT 1835.030 2726.275 1835.310 2726.645 ;
        RECT 403.510 2725.595 403.790 2725.965 ;
        RECT 524.030 2725.595 524.310 2725.965 ;
        RECT 627.070 2725.595 627.350 2725.965 ;
        RECT 724.130 2725.595 724.410 2725.965 ;
        RECT 1110.070 2725.595 1110.350 2725.965 ;
        RECT 1207.130 2725.595 1207.410 2725.965 ;
        RECT 1303.730 2725.595 1304.010 2725.965 ;
        RECT 403.580 2724.605 403.720 2725.595 ;
        RECT 1835.100 2724.605 1835.240 2726.275 ;
        RECT 1859.480 2725.965 1859.620 2727.635 ;
        RECT 2801.500 2727.490 2801.760 2727.635 ;
        RECT 2815.760 2727.490 2816.020 2727.810 ;
        RECT 2897.630 2727.635 2897.910 2728.005 ;
        RECT 2415.090 2726.955 2415.370 2727.325 ;
        RECT 2415.100 2726.810 2415.360 2726.955 ;
        RECT 2429.360 2726.810 2429.620 2727.130 ;
        RECT 2704.890 2726.955 2705.170 2727.325 ;
        RECT 2704.900 2726.810 2705.160 2726.955 ;
        RECT 2743.080 2726.810 2743.340 2727.130 ;
        RECT 2429.420 2725.965 2429.560 2726.810 ;
        RECT 2743.140 2725.965 2743.280 2726.810 ;
        RECT 2815.820 2726.645 2815.960 2727.490 ;
        RECT 2897.700 2727.470 2897.840 2727.635 ;
        RECT 2863.140 2727.325 2863.400 2727.470 ;
        RECT 2863.130 2726.955 2863.410 2727.325 ;
        RECT 2897.640 2727.150 2897.900 2727.470 ;
        RECT 2815.750 2726.275 2816.030 2726.645 ;
        RECT 1859.410 2725.595 1859.690 2725.965 ;
        RECT 2429.350 2725.595 2429.630 2725.965 ;
        RECT 2743.070 2725.595 2743.350 2725.965 ;
        RECT 403.510 2724.235 403.790 2724.605 ;
        RECT 1835.030 2724.235 1835.310 2724.605 ;
      LAYER via2 ;
        RECT 1037.850 2728.360 1038.130 2728.640 ;
        RECT 1545.230 2727.680 1545.510 2727.960 ;
        RECT 1859.410 2727.680 1859.690 2727.960 ;
        RECT 2766.530 2727.680 2766.810 2727.960 ;
        RECT 2767.450 2727.680 2767.730 2727.960 ;
        RECT 2801.490 2727.680 2801.770 2727.960 ;
        RECT 579.690 2727.000 579.970 2727.280 ;
        RECT 676.290 2727.000 676.570 2727.280 ;
        RECT 979.430 2727.000 979.710 2727.280 ;
        RECT 1007.030 2727.000 1007.310 2727.280 ;
        RECT 1037.850 2727.000 1038.130 2727.280 ;
        RECT 1062.690 2727.000 1062.970 2727.280 ;
        RECT 1159.290 2727.000 1159.570 2727.280 ;
        RECT 1255.890 2727.000 1256.170 2727.280 ;
        RECT 1510.730 2727.000 1511.010 2727.280 ;
        RECT 1641.830 2727.000 1642.110 2727.280 ;
        RECT 1738.430 2727.000 1738.710 2727.280 ;
        RECT 427.890 2726.320 428.170 2726.600 ;
        RECT 475.270 2726.320 475.550 2726.600 ;
        RECT 483.090 2726.320 483.370 2726.600 ;
        RECT 834.530 2726.320 834.810 2726.600 ;
        RECT 886.510 2726.320 886.790 2726.600 ;
        RECT 1607.330 2726.320 1607.610 2726.600 ;
        RECT 1738.430 2726.320 1738.710 2726.600 ;
        RECT 1835.030 2726.320 1835.310 2726.600 ;
        RECT 403.510 2725.640 403.790 2725.920 ;
        RECT 524.030 2725.640 524.310 2725.920 ;
        RECT 627.070 2725.640 627.350 2725.920 ;
        RECT 724.130 2725.640 724.410 2725.920 ;
        RECT 1110.070 2725.640 1110.350 2725.920 ;
        RECT 1207.130 2725.640 1207.410 2725.920 ;
        RECT 1303.730 2725.640 1304.010 2725.920 ;
        RECT 2897.630 2727.680 2897.910 2727.960 ;
        RECT 2415.090 2727.000 2415.370 2727.280 ;
        RECT 2704.890 2727.000 2705.170 2727.280 ;
        RECT 2863.130 2727.000 2863.410 2727.280 ;
        RECT 2815.750 2726.320 2816.030 2726.600 ;
        RECT 1859.410 2725.640 1859.690 2725.920 ;
        RECT 2429.350 2725.640 2429.630 2725.920 ;
        RECT 2743.070 2725.640 2743.350 2725.920 ;
        RECT 403.510 2724.280 403.790 2724.560 ;
        RECT 1835.030 2724.280 1835.310 2724.560 ;
      LAYER met3 ;
        RECT 1037.825 2728.650 1038.155 2728.665 ;
        RECT 1014.150 2728.350 1038.155 2728.650 ;
        RECT 287.310 2727.970 287.690 2727.980 ;
        RECT 287.310 2727.670 304.210 2727.970 ;
        RECT 287.310 2727.660 287.690 2727.670 ;
        RECT 303.910 2726.610 304.210 2727.670 ;
        RECT 579.665 2727.290 579.995 2727.305 ;
        RECT 676.265 2727.290 676.595 2727.305 ;
        RECT 979.405 2727.290 979.735 2727.305 ;
        RECT 544.950 2726.990 579.995 2727.290 ;
        RECT 427.865 2726.610 428.195 2726.625 ;
        RECT 303.910 2726.310 362.170 2726.610 ;
        RECT 361.870 2725.930 362.170 2726.310 ;
        RECT 427.190 2726.310 428.195 2726.610 ;
        RECT 379.310 2725.930 379.690 2725.940 ;
        RECT 361.870 2725.630 379.690 2725.930 ;
        RECT 379.310 2725.620 379.690 2725.630 ;
        RECT 403.485 2725.930 403.815 2725.945 ;
        RECT 427.190 2725.930 427.490 2726.310 ;
        RECT 427.865 2726.295 428.195 2726.310 ;
        RECT 475.245 2726.610 475.575 2726.625 ;
        RECT 483.065 2726.610 483.395 2726.625 ;
        RECT 475.245 2726.310 483.395 2726.610 ;
        RECT 475.245 2726.295 475.575 2726.310 ;
        RECT 483.065 2726.295 483.395 2726.310 ;
        RECT 403.485 2725.630 427.490 2725.930 ;
        RECT 524.005 2725.930 524.335 2725.945 ;
        RECT 544.950 2725.930 545.250 2726.990 ;
        RECT 579.665 2726.975 579.995 2726.990 ;
        RECT 641.550 2726.990 676.595 2727.290 ;
        RECT 524.005 2725.630 545.250 2725.930 ;
        RECT 627.045 2725.930 627.375 2725.945 ;
        RECT 641.550 2725.930 641.850 2726.990 ;
        RECT 676.265 2726.975 676.595 2726.990 ;
        RECT 738.150 2726.990 787.210 2727.290 ;
        RECT 627.045 2725.630 641.850 2725.930 ;
        RECT 724.105 2725.930 724.435 2725.945 ;
        RECT 738.150 2725.930 738.450 2726.990 ;
        RECT 786.910 2726.610 787.210 2726.990 ;
        RECT 958.950 2726.990 979.735 2727.290 ;
        RECT 834.505 2726.610 834.835 2726.625 ;
        RECT 786.910 2726.310 834.835 2726.610 ;
        RECT 834.505 2726.295 834.835 2726.310 ;
        RECT 886.485 2726.610 886.815 2726.625 ;
        RECT 958.950 2726.610 959.250 2726.990 ;
        RECT 979.405 2726.975 979.735 2726.990 ;
        RECT 1007.005 2727.290 1007.335 2727.305 ;
        RECT 1014.150 2727.290 1014.450 2728.350 ;
        RECT 1037.825 2728.335 1038.155 2728.350 ;
        RECT 1545.205 2727.970 1545.535 2727.985 ;
        RECT 1859.385 2727.970 1859.715 2727.985 ;
        RECT 1545.205 2727.670 1560.010 2727.970 ;
        RECT 1545.205 2727.655 1545.535 2727.670 ;
        RECT 1007.005 2726.990 1014.450 2727.290 ;
        RECT 1037.825 2727.290 1038.155 2727.305 ;
        RECT 1062.665 2727.290 1062.995 2727.305 ;
        RECT 1159.265 2727.290 1159.595 2727.305 ;
        RECT 1255.865 2727.290 1256.195 2727.305 ;
        RECT 1510.705 2727.290 1511.035 2727.305 ;
        RECT 1037.825 2726.990 1062.995 2727.290 ;
        RECT 1007.005 2726.975 1007.335 2726.990 ;
        RECT 1037.825 2726.975 1038.155 2726.990 ;
        RECT 1062.665 2726.975 1062.995 2726.990 ;
        RECT 1124.550 2726.990 1159.595 2727.290 ;
        RECT 886.485 2726.310 959.250 2726.610 ;
        RECT 886.485 2726.295 886.815 2726.310 ;
        RECT 724.105 2725.630 738.450 2725.930 ;
        RECT 1110.045 2725.930 1110.375 2725.945 ;
        RECT 1124.550 2725.930 1124.850 2726.990 ;
        RECT 1159.265 2726.975 1159.595 2726.990 ;
        RECT 1221.150 2726.990 1256.195 2727.290 ;
        RECT 1110.045 2725.630 1124.850 2725.930 ;
        RECT 1207.105 2725.930 1207.435 2725.945 ;
        RECT 1221.150 2725.930 1221.450 2726.990 ;
        RECT 1255.865 2726.975 1256.195 2726.990 ;
        RECT 1317.750 2726.990 1414.650 2727.290 ;
        RECT 1207.105 2725.630 1221.450 2725.930 ;
        RECT 1303.705 2725.930 1304.035 2725.945 ;
        RECT 1317.750 2725.930 1318.050 2726.990 ;
        RECT 1414.350 2726.610 1414.650 2726.990 ;
        RECT 1463.110 2726.990 1511.035 2727.290 ;
        RECT 1414.350 2726.310 1462.490 2726.610 ;
        RECT 1303.705 2725.630 1318.050 2725.930 ;
        RECT 1462.190 2725.930 1462.490 2726.310 ;
        RECT 1463.110 2725.930 1463.410 2726.990 ;
        RECT 1510.705 2726.975 1511.035 2726.990 ;
        RECT 1559.710 2726.610 1560.010 2727.670 ;
        RECT 1835.710 2727.670 1859.715 2727.970 ;
        RECT 1641.805 2727.290 1642.135 2727.305 ;
        RECT 1738.405 2727.290 1738.735 2727.305 ;
        RECT 1739.070 2727.290 1739.450 2727.300 ;
        RECT 1641.805 2726.990 1656.610 2727.290 ;
        RECT 1641.805 2726.975 1642.135 2726.990 ;
        RECT 1607.305 2726.610 1607.635 2726.625 ;
        RECT 1559.710 2726.310 1607.635 2726.610 ;
        RECT 1656.310 2726.610 1656.610 2726.990 ;
        RECT 1738.405 2726.990 1739.450 2727.290 ;
        RECT 1738.405 2726.975 1738.735 2726.990 ;
        RECT 1739.070 2726.980 1739.450 2726.990 ;
        RECT 1738.405 2726.610 1738.735 2726.625 ;
        RECT 1656.310 2726.310 1738.735 2726.610 ;
        RECT 1607.305 2726.295 1607.635 2726.310 ;
        RECT 1738.405 2726.295 1738.735 2726.310 ;
        RECT 1835.005 2726.610 1835.335 2726.625 ;
        RECT 1835.710 2726.610 1836.010 2727.670 ;
        RECT 1859.385 2727.655 1859.715 2727.670 ;
        RECT 2752.910 2727.970 2753.290 2727.980 ;
        RECT 2766.505 2727.970 2766.835 2727.985 ;
        RECT 2752.910 2727.670 2766.835 2727.970 ;
        RECT 2752.910 2727.660 2753.290 2727.670 ;
        RECT 2766.505 2727.655 2766.835 2727.670 ;
        RECT 2767.425 2727.970 2767.755 2727.985 ;
        RECT 2801.465 2727.970 2801.795 2727.985 ;
        RECT 2767.425 2727.670 2801.795 2727.970 ;
        RECT 2767.425 2727.655 2767.755 2727.670 ;
        RECT 2801.465 2727.655 2801.795 2727.670 ;
        RECT 2897.605 2727.970 2897.935 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2897.605 2727.670 2924.800 2727.970 ;
        RECT 2897.605 2727.655 2897.935 2727.670 ;
        RECT 1883.510 2727.290 1883.890 2727.300 ;
        RECT 2415.065 2727.290 2415.395 2727.305 ;
        RECT 1883.510 2726.990 1966.650 2727.290 ;
        RECT 1883.510 2726.980 1883.890 2726.990 ;
        RECT 1835.005 2726.310 1836.010 2726.610 ;
        RECT 1966.350 2726.610 1966.650 2726.990 ;
        RECT 2015.110 2726.990 2138.690 2727.290 ;
        RECT 1966.350 2726.310 2014.490 2726.610 ;
        RECT 1835.005 2726.295 1835.335 2726.310 ;
        RECT 1462.190 2725.630 1463.410 2725.930 ;
        RECT 1739.070 2725.930 1739.450 2725.940 ;
        RECT 1786.910 2725.930 1787.290 2725.940 ;
        RECT 1739.070 2725.630 1787.290 2725.930 ;
        RECT 403.485 2725.615 403.815 2725.630 ;
        RECT 524.005 2725.615 524.335 2725.630 ;
        RECT 627.045 2725.615 627.375 2725.630 ;
        RECT 724.105 2725.615 724.435 2725.630 ;
        RECT 1110.045 2725.615 1110.375 2725.630 ;
        RECT 1207.105 2725.615 1207.435 2725.630 ;
        RECT 1303.705 2725.615 1304.035 2725.630 ;
        RECT 1739.070 2725.620 1739.450 2725.630 ;
        RECT 1786.910 2725.620 1787.290 2725.630 ;
        RECT 1859.385 2725.930 1859.715 2725.945 ;
        RECT 1883.510 2725.930 1883.890 2725.940 ;
        RECT 1859.385 2725.630 1883.890 2725.930 ;
        RECT 2014.190 2725.930 2014.490 2726.310 ;
        RECT 2015.110 2725.930 2015.410 2726.990 ;
        RECT 2014.190 2725.630 2015.410 2725.930 ;
        RECT 1859.385 2725.615 1859.715 2725.630 ;
        RECT 1883.510 2725.620 1883.890 2725.630 ;
        RECT 2138.390 2725.250 2138.690 2726.990 ;
        RECT 2208.310 2726.990 2256.450 2727.290 ;
        RECT 2208.310 2725.930 2208.610 2726.990 ;
        RECT 2256.150 2726.610 2256.450 2726.990 ;
        RECT 2304.910 2726.990 2353.050 2727.290 ;
        RECT 2256.150 2726.310 2304.290 2726.610 ;
        RECT 2173.350 2725.630 2208.610 2725.930 ;
        RECT 2303.990 2725.930 2304.290 2726.310 ;
        RECT 2304.910 2725.930 2305.210 2726.990 ;
        RECT 2352.750 2726.610 2353.050 2726.990 ;
        RECT 2401.510 2726.990 2415.395 2727.290 ;
        RECT 2352.750 2726.310 2400.890 2726.610 ;
        RECT 2303.990 2725.630 2305.210 2725.930 ;
        RECT 2400.590 2725.930 2400.890 2726.310 ;
        RECT 2401.510 2725.930 2401.810 2726.990 ;
        RECT 2415.065 2726.975 2415.395 2726.990 ;
        RECT 2463.110 2727.290 2463.490 2727.300 ;
        RECT 2704.865 2727.290 2705.195 2727.305 ;
        RECT 2863.105 2727.290 2863.435 2727.305 ;
        RECT 2463.110 2726.990 2546.250 2727.290 ;
        RECT 2463.110 2726.980 2463.490 2726.990 ;
        RECT 2545.950 2726.610 2546.250 2726.990 ;
        RECT 2594.710 2726.990 2642.850 2727.290 ;
        RECT 2545.950 2726.310 2594.090 2726.610 ;
        RECT 2400.590 2725.630 2401.810 2725.930 ;
        RECT 2429.325 2725.930 2429.655 2725.945 ;
        RECT 2463.110 2725.930 2463.490 2725.940 ;
        RECT 2429.325 2725.630 2463.490 2725.930 ;
        RECT 2593.790 2725.930 2594.090 2726.310 ;
        RECT 2594.710 2725.930 2595.010 2726.990 ;
        RECT 2642.550 2726.610 2642.850 2726.990 ;
        RECT 2691.310 2726.990 2705.195 2727.290 ;
        RECT 2642.550 2726.310 2690.690 2726.610 ;
        RECT 2593.790 2725.630 2595.010 2725.930 ;
        RECT 2690.390 2725.930 2690.690 2726.310 ;
        RECT 2691.310 2725.930 2691.610 2726.990 ;
        RECT 2704.865 2726.975 2705.195 2726.990 ;
        RECT 2849.550 2726.990 2863.435 2727.290 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2815.725 2726.610 2816.055 2726.625 ;
        RECT 2849.550 2726.610 2849.850 2726.990 ;
        RECT 2863.105 2726.975 2863.435 2726.990 ;
        RECT 2815.725 2726.310 2849.850 2726.610 ;
        RECT 2815.725 2726.295 2816.055 2726.310 ;
        RECT 2690.390 2725.630 2691.610 2725.930 ;
        RECT 2743.045 2725.930 2743.375 2725.945 ;
        RECT 2752.910 2725.930 2753.290 2725.940 ;
        RECT 2743.045 2725.630 2753.290 2725.930 ;
        RECT 2173.350 2725.250 2173.650 2725.630 ;
        RECT 2429.325 2725.615 2429.655 2725.630 ;
        RECT 2463.110 2725.620 2463.490 2725.630 ;
        RECT 2743.045 2725.615 2743.375 2725.630 ;
        RECT 2752.910 2725.620 2753.290 2725.630 ;
        RECT 2138.390 2724.950 2173.650 2725.250 ;
        RECT 379.310 2724.570 379.690 2724.580 ;
        RECT 403.485 2724.570 403.815 2724.585 ;
        RECT 379.310 2724.270 403.815 2724.570 ;
        RECT 379.310 2724.260 379.690 2724.270 ;
        RECT 403.485 2724.255 403.815 2724.270 ;
        RECT 1786.910 2724.570 1787.290 2724.580 ;
        RECT 1835.005 2724.570 1835.335 2724.585 ;
        RECT 1786.910 2724.270 1835.335 2724.570 ;
        RECT 1786.910 2724.260 1787.290 2724.270 ;
        RECT 1835.005 2724.255 1835.335 2724.270 ;
        RECT 287.310 1942.570 287.690 1942.580 ;
        RECT 300.000 1942.570 304.000 1942.680 ;
        RECT 287.310 1942.270 304.000 1942.570 ;
        RECT 287.310 1942.260 287.690 1942.270 ;
        RECT 300.000 1942.080 304.000 1942.270 ;
      LAYER via3 ;
        RECT 287.340 2727.660 287.660 2727.980 ;
        RECT 379.340 2725.620 379.660 2725.940 ;
        RECT 1739.100 2726.980 1739.420 2727.300 ;
        RECT 2752.940 2727.660 2753.260 2727.980 ;
        RECT 1883.540 2726.980 1883.860 2727.300 ;
        RECT 1739.100 2725.620 1739.420 2725.940 ;
        RECT 1786.940 2725.620 1787.260 2725.940 ;
        RECT 1883.540 2725.620 1883.860 2725.940 ;
        RECT 2463.140 2726.980 2463.460 2727.300 ;
        RECT 2463.140 2725.620 2463.460 2725.940 ;
        RECT 2752.940 2725.620 2753.260 2725.940 ;
        RECT 379.340 2724.260 379.660 2724.580 ;
        RECT 1786.940 2724.260 1787.260 2724.580 ;
        RECT 287.340 1942.260 287.660 1942.580 ;
      LAYER met4 ;
        RECT 287.335 2727.655 287.665 2727.985 ;
        RECT 2752.935 2727.655 2753.265 2727.985 ;
        RECT 287.350 1942.585 287.650 2727.655 ;
        RECT 1739.095 2726.975 1739.425 2727.305 ;
        RECT 1883.535 2726.975 1883.865 2727.305 ;
        RECT 2463.135 2726.975 2463.465 2727.305 ;
        RECT 1739.110 2725.945 1739.410 2726.975 ;
        RECT 1883.550 2725.945 1883.850 2726.975 ;
        RECT 2463.150 2725.945 2463.450 2726.975 ;
        RECT 2752.950 2725.945 2753.250 2727.655 ;
        RECT 379.335 2725.615 379.665 2725.945 ;
        RECT 1739.095 2725.615 1739.425 2725.945 ;
        RECT 1786.935 2725.615 1787.265 2725.945 ;
        RECT 1883.535 2725.615 1883.865 2725.945 ;
        RECT 2463.135 2725.615 2463.465 2725.945 ;
        RECT 2752.935 2725.615 2753.265 2725.945 ;
        RECT 379.350 2724.585 379.650 2725.615 ;
        RECT 1786.950 2724.585 1787.250 2725.615 ;
        RECT 379.335 2724.255 379.665 2724.585 ;
        RECT 1786.935 2724.255 1787.265 2724.585 ;
        RECT 287.335 1942.255 287.665 1942.585 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2903.150 2962.235 2903.430 2962.605 ;
        RECT 2903.220 2701.485 2903.360 2962.235 ;
        RECT 2903.150 2701.115 2903.430 2701.485 ;
      LAYER via2 ;
        RECT 2903.150 2962.280 2903.430 2962.560 ;
        RECT 2903.150 2701.160 2903.430 2701.440 ;
      LAYER met3 ;
        RECT 2903.125 2962.570 2903.455 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2903.125 2962.270 2924.800 2962.570 ;
        RECT 2903.125 2962.255 2903.455 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 286.390 2701.450 286.770 2701.460 ;
        RECT 2903.125 2701.450 2903.455 2701.465 ;
        RECT 286.390 2701.150 2903.455 2701.450 ;
        RECT 286.390 2701.140 286.770 2701.150 ;
        RECT 2903.125 2701.135 2903.455 2701.150 ;
        RECT 286.390 1971.810 286.770 1971.820 ;
        RECT 300.000 1971.810 304.000 1971.920 ;
        RECT 286.390 1971.510 304.000 1971.810 ;
        RECT 286.390 1971.500 286.770 1971.510 ;
        RECT 300.000 1971.320 304.000 1971.510 ;
      LAYER via3 ;
        RECT 286.420 2701.140 286.740 2701.460 ;
        RECT 286.420 1971.500 286.740 1971.820 ;
      LAYER met4 ;
        RECT 286.415 2701.135 286.745 2701.465 ;
        RECT 286.430 1971.825 286.730 2701.135 ;
        RECT 286.415 1971.495 286.745 1971.825 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 290.330 2701.540 290.650 2701.600 ;
        RECT 2901.290 2701.540 2901.610 2701.600 ;
        RECT 290.330 2701.400 2901.610 2701.540 ;
        RECT 290.330 2701.340 290.650 2701.400 ;
        RECT 2901.290 2701.340 2901.610 2701.400 ;
      LAYER via ;
        RECT 290.360 2701.340 290.620 2701.600 ;
        RECT 2901.320 2701.340 2901.580 2701.600 ;
      LAYER met2 ;
        RECT 2901.310 3196.835 2901.590 3197.205 ;
        RECT 2901.380 2701.630 2901.520 3196.835 ;
        RECT 290.360 2701.310 290.620 2701.630 ;
        RECT 2901.320 2701.310 2901.580 2701.630 ;
        RECT 290.420 2000.405 290.560 2701.310 ;
        RECT 290.350 2000.035 290.630 2000.405 ;
      LAYER via2 ;
        RECT 2901.310 3196.880 2901.590 3197.160 ;
        RECT 290.350 2000.080 290.630 2000.360 ;
      LAYER met3 ;
        RECT 2901.285 3197.170 2901.615 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2901.285 3196.870 2924.800 3197.170 ;
        RECT 2901.285 3196.855 2901.615 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 290.325 2000.370 290.655 2000.385 ;
        RECT 300.000 2000.370 304.000 2000.480 ;
        RECT 290.325 2000.070 304.000 2000.370 ;
        RECT 290.325 2000.055 290.655 2000.070 ;
        RECT 300.000 1999.880 304.000 2000.070 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 869.470 3431.520 869.790 3431.580 ;
        RECT 893.850 3431.520 894.170 3431.580 ;
        RECT 869.470 3431.380 894.170 3431.520 ;
        RECT 869.470 3431.320 869.790 3431.380 ;
        RECT 893.850 3431.320 894.170 3431.380 ;
        RECT 1835.470 3431.520 1835.790 3431.580 ;
        RECT 1859.850 3431.520 1860.170 3431.580 ;
        RECT 1835.470 3431.380 1860.170 3431.520 ;
        RECT 1835.470 3431.320 1835.790 3431.380 ;
        RECT 1859.850 3431.320 1860.170 3431.380 ;
        RECT 2801.470 3431.520 2801.790 3431.580 ;
        RECT 2825.850 3431.520 2826.170 3431.580 ;
        RECT 2801.470 3431.380 2826.170 3431.520 ;
        RECT 2801.470 3431.320 2801.790 3431.380 ;
        RECT 2825.850 3431.320 2826.170 3431.380 ;
        RECT 772.870 3430.840 773.190 3430.900 ;
        RECT 811.050 3430.840 811.370 3430.900 ;
        RECT 772.870 3430.700 811.370 3430.840 ;
        RECT 772.870 3430.640 773.190 3430.700 ;
        RECT 811.050 3430.640 811.370 3430.700 ;
        RECT 1449.070 3430.840 1449.390 3430.900 ;
        RECT 1472.530 3430.840 1472.850 3430.900 ;
        RECT 1449.070 3430.700 1472.850 3430.840 ;
        RECT 1449.070 3430.640 1449.390 3430.700 ;
        RECT 1472.530 3430.640 1472.850 3430.700 ;
        RECT 1738.870 3430.840 1739.190 3430.900 ;
        RECT 1777.050 3430.840 1777.370 3430.900 ;
        RECT 1738.870 3430.700 1777.370 3430.840 ;
        RECT 1738.870 3430.640 1739.190 3430.700 ;
        RECT 1777.050 3430.640 1777.370 3430.700 ;
        RECT 2704.870 3430.840 2705.190 3430.900 ;
        RECT 2743.050 3430.840 2743.370 3430.900 ;
        RECT 2704.870 3430.700 2743.370 3430.840 ;
        RECT 2704.870 3430.640 2705.190 3430.700 ;
        RECT 2743.050 3430.640 2743.370 3430.700 ;
      LAYER via ;
        RECT 869.500 3431.320 869.760 3431.580 ;
        RECT 893.880 3431.320 894.140 3431.580 ;
        RECT 1835.500 3431.320 1835.760 3431.580 ;
        RECT 1859.880 3431.320 1860.140 3431.580 ;
        RECT 2801.500 3431.320 2801.760 3431.580 ;
        RECT 2825.880 3431.320 2826.140 3431.580 ;
        RECT 772.900 3430.640 773.160 3430.900 ;
        RECT 811.080 3430.640 811.340 3430.900 ;
        RECT 1449.100 3430.640 1449.360 3430.900 ;
        RECT 1472.560 3430.640 1472.820 3430.900 ;
        RECT 1738.900 3430.640 1739.160 3430.900 ;
        RECT 1777.080 3430.640 1777.340 3430.900 ;
        RECT 2704.900 3430.640 2705.160 3430.900 ;
        RECT 2743.080 3430.640 2743.340 3430.900 ;
      LAYER met2 ;
        RECT 941.710 3432.115 941.990 3432.485 ;
        RECT 1897.590 3432.115 1897.870 3432.485 ;
        RECT 2207.630 3432.115 2207.910 3432.485 ;
        RECT 834.530 3431.690 834.810 3431.805 ;
        RECT 835.450 3431.690 835.730 3431.805 ;
        RECT 834.530 3431.550 835.730 3431.690 ;
        RECT 834.530 3431.435 834.810 3431.550 ;
        RECT 835.450 3431.435 835.730 3431.550 ;
        RECT 869.490 3431.435 869.770 3431.805 ;
        RECT 869.500 3431.290 869.760 3431.435 ;
        RECT 893.880 3431.290 894.140 3431.610 ;
        RECT 893.940 3431.125 894.080 3431.290 ;
        RECT 941.780 3431.125 941.920 3432.115 ;
        RECT 1800.530 3431.690 1800.810 3431.805 ;
        RECT 1801.450 3431.690 1801.730 3431.805 ;
        RECT 1800.530 3431.550 1801.730 3431.690 ;
        RECT 1800.530 3431.435 1800.810 3431.550 ;
        RECT 1801.450 3431.435 1801.730 3431.550 ;
        RECT 1835.490 3431.435 1835.770 3431.805 ;
        RECT 1835.500 3431.290 1835.760 3431.435 ;
        RECT 1859.880 3431.290 1860.140 3431.610 ;
        RECT 1859.940 3431.125 1860.080 3431.290 ;
        RECT 1897.660 3431.125 1897.800 3432.115 ;
        RECT 2207.700 3431.125 2207.840 3432.115 ;
        RECT 2766.530 3431.690 2766.810 3431.805 ;
        RECT 2767.450 3431.690 2767.730 3431.805 ;
        RECT 2766.530 3431.550 2767.730 3431.690 ;
        RECT 2766.530 3431.435 2766.810 3431.550 ;
        RECT 2767.450 3431.435 2767.730 3431.550 ;
        RECT 2801.490 3431.435 2801.770 3431.805 ;
        RECT 2801.500 3431.290 2801.760 3431.435 ;
        RECT 2825.880 3431.290 2826.140 3431.610 ;
        RECT 2825.940 3431.125 2826.080 3431.290 ;
        RECT 772.890 3430.755 773.170 3431.125 ;
        RECT 772.900 3430.610 773.160 3430.755 ;
        RECT 811.080 3430.610 811.340 3430.930 ;
        RECT 893.870 3430.755 894.150 3431.125 ;
        RECT 941.710 3430.755 941.990 3431.125 ;
        RECT 1449.090 3430.755 1449.370 3431.125 ;
        RECT 1449.100 3430.610 1449.360 3430.755 ;
        RECT 1472.560 3430.610 1472.820 3430.930 ;
        RECT 1738.890 3430.755 1739.170 3431.125 ;
        RECT 1738.900 3430.610 1739.160 3430.755 ;
        RECT 1777.080 3430.610 1777.340 3430.930 ;
        RECT 1859.870 3430.755 1860.150 3431.125 ;
        RECT 1897.590 3430.755 1897.870 3431.125 ;
        RECT 2137.710 3431.010 2137.990 3431.125 ;
        RECT 2138.630 3431.010 2138.910 3431.125 ;
        RECT 2137.710 3430.870 2138.910 3431.010 ;
        RECT 2137.710 3430.755 2137.990 3430.870 ;
        RECT 2138.630 3430.755 2138.910 3430.870 ;
        RECT 2207.630 3430.755 2207.910 3431.125 ;
        RECT 2704.890 3430.755 2705.170 3431.125 ;
        RECT 2704.900 3430.610 2705.160 3430.755 ;
        RECT 2743.080 3430.610 2743.340 3430.930 ;
        RECT 2825.870 3430.755 2826.150 3431.125 ;
        RECT 2863.590 3431.010 2863.870 3431.125 ;
        RECT 2863.200 3430.870 2863.870 3431.010 ;
        RECT 811.140 3429.765 811.280 3430.610 ;
        RECT 1472.620 3429.765 1472.760 3430.610 ;
        RECT 1777.140 3429.765 1777.280 3430.610 ;
        RECT 2743.140 3429.765 2743.280 3430.610 ;
        RECT 2863.200 3430.445 2863.340 3430.870 ;
        RECT 2863.590 3430.755 2863.870 3430.870 ;
        RECT 2863.130 3430.075 2863.410 3430.445 ;
        RECT 811.070 3429.395 811.350 3429.765 ;
        RECT 1472.550 3429.395 1472.830 3429.765 ;
        RECT 1777.070 3429.395 1777.350 3429.765 ;
        RECT 2743.070 3429.395 2743.350 3429.765 ;
      LAYER via2 ;
        RECT 941.710 3432.160 941.990 3432.440 ;
        RECT 1897.590 3432.160 1897.870 3432.440 ;
        RECT 2207.630 3432.160 2207.910 3432.440 ;
        RECT 834.530 3431.480 834.810 3431.760 ;
        RECT 835.450 3431.480 835.730 3431.760 ;
        RECT 869.490 3431.480 869.770 3431.760 ;
        RECT 1800.530 3431.480 1800.810 3431.760 ;
        RECT 1801.450 3431.480 1801.730 3431.760 ;
        RECT 1835.490 3431.480 1835.770 3431.760 ;
        RECT 2766.530 3431.480 2766.810 3431.760 ;
        RECT 2767.450 3431.480 2767.730 3431.760 ;
        RECT 2801.490 3431.480 2801.770 3431.760 ;
        RECT 772.890 3430.800 773.170 3431.080 ;
        RECT 893.870 3430.800 894.150 3431.080 ;
        RECT 941.710 3430.800 941.990 3431.080 ;
        RECT 1449.090 3430.800 1449.370 3431.080 ;
        RECT 1738.890 3430.800 1739.170 3431.080 ;
        RECT 1859.870 3430.800 1860.150 3431.080 ;
        RECT 1897.590 3430.800 1897.870 3431.080 ;
        RECT 2137.710 3430.800 2137.990 3431.080 ;
        RECT 2138.630 3430.800 2138.910 3431.080 ;
        RECT 2207.630 3430.800 2207.910 3431.080 ;
        RECT 2704.890 3430.800 2705.170 3431.080 ;
        RECT 2825.870 3430.800 2826.150 3431.080 ;
        RECT 2863.590 3430.800 2863.870 3431.080 ;
        RECT 2863.130 3430.120 2863.410 3430.400 ;
        RECT 811.070 3429.440 811.350 3429.720 ;
        RECT 1472.550 3429.440 1472.830 3429.720 ;
        RECT 1777.070 3429.440 1777.350 3429.720 ;
        RECT 2743.070 3429.440 2743.350 3429.720 ;
      LAYER met3 ;
        RECT 917.510 3432.450 917.890 3432.460 ;
        RECT 941.685 3432.450 942.015 3432.465 ;
        RECT 917.510 3432.150 942.015 3432.450 ;
        RECT 917.510 3432.140 917.890 3432.150 ;
        RECT 941.685 3432.135 942.015 3432.150 ;
        RECT 1883.510 3432.450 1883.890 3432.460 ;
        RECT 1897.565 3432.450 1897.895 3432.465 ;
        RECT 1883.510 3432.150 1897.895 3432.450 ;
        RECT 1883.510 3432.140 1883.890 3432.150 ;
        RECT 1897.565 3432.135 1897.895 3432.150 ;
        RECT 2173.310 3432.450 2173.690 3432.460 ;
        RECT 2207.605 3432.450 2207.935 3432.465 ;
        RECT 2173.310 3432.150 2207.935 3432.450 ;
        RECT 2173.310 3432.140 2173.690 3432.150 ;
        RECT 2207.605 3432.135 2207.935 3432.150 ;
        RECT 820.910 3431.770 821.290 3431.780 ;
        RECT 834.505 3431.770 834.835 3431.785 ;
        RECT 820.910 3431.470 834.835 3431.770 ;
        RECT 820.910 3431.460 821.290 3431.470 ;
        RECT 834.505 3431.455 834.835 3431.470 ;
        RECT 835.425 3431.770 835.755 3431.785 ;
        RECT 869.465 3431.770 869.795 3431.785 ;
        RECT 835.425 3431.470 869.795 3431.770 ;
        RECT 835.425 3431.455 835.755 3431.470 ;
        RECT 869.465 3431.455 869.795 3431.470 ;
        RECT 1786.910 3431.770 1787.290 3431.780 ;
        RECT 1800.505 3431.770 1800.835 3431.785 ;
        RECT 1786.910 3431.470 1800.835 3431.770 ;
        RECT 1786.910 3431.460 1787.290 3431.470 ;
        RECT 1800.505 3431.455 1800.835 3431.470 ;
        RECT 1801.425 3431.770 1801.755 3431.785 ;
        RECT 1835.465 3431.770 1835.795 3431.785 ;
        RECT 1801.425 3431.470 1835.795 3431.770 ;
        RECT 1801.425 3431.455 1801.755 3431.470 ;
        RECT 1835.465 3431.455 1835.795 3431.470 ;
        RECT 2752.910 3431.770 2753.290 3431.780 ;
        RECT 2766.505 3431.770 2766.835 3431.785 ;
        RECT 2752.910 3431.470 2766.835 3431.770 ;
        RECT 2752.910 3431.460 2753.290 3431.470 ;
        RECT 2766.505 3431.455 2766.835 3431.470 ;
        RECT 2767.425 3431.770 2767.755 3431.785 ;
        RECT 2801.465 3431.770 2801.795 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2767.425 3431.470 2801.795 3431.770 ;
        RECT 2767.425 3431.455 2767.755 3431.470 ;
        RECT 2801.465 3431.455 2801.795 3431.470 ;
        RECT 2916.710 3431.470 2924.800 3431.770 ;
        RECT 288.230 3431.090 288.610 3431.100 ;
        RECT 772.865 3431.090 773.195 3431.105 ;
        RECT 288.230 3430.790 324.450 3431.090 ;
        RECT 288.230 3430.780 288.610 3430.790 ;
        RECT 324.150 3430.410 324.450 3430.790 ;
        RECT 372.910 3430.790 421.050 3431.090 ;
        RECT 324.150 3430.110 372.290 3430.410 ;
        RECT 371.990 3429.730 372.290 3430.110 ;
        RECT 372.910 3429.730 373.210 3430.790 ;
        RECT 420.750 3430.410 421.050 3430.790 ;
        RECT 469.510 3430.790 517.650 3431.090 ;
        RECT 420.750 3430.110 468.890 3430.410 ;
        RECT 371.990 3429.430 373.210 3429.730 ;
        RECT 468.590 3429.730 468.890 3430.110 ;
        RECT 469.510 3429.730 469.810 3430.790 ;
        RECT 517.350 3430.410 517.650 3430.790 ;
        RECT 566.110 3430.790 614.250 3431.090 ;
        RECT 517.350 3430.110 565.490 3430.410 ;
        RECT 468.590 3429.430 469.810 3429.730 ;
        RECT 565.190 3429.730 565.490 3430.110 ;
        RECT 566.110 3429.730 566.410 3430.790 ;
        RECT 613.950 3430.410 614.250 3430.790 ;
        RECT 662.710 3430.790 710.850 3431.090 ;
        RECT 613.950 3430.110 662.090 3430.410 ;
        RECT 565.190 3429.430 566.410 3429.730 ;
        RECT 661.790 3429.730 662.090 3430.110 ;
        RECT 662.710 3429.730 663.010 3430.790 ;
        RECT 710.550 3430.410 710.850 3430.790 ;
        RECT 759.310 3430.790 773.195 3431.090 ;
        RECT 710.550 3430.110 758.690 3430.410 ;
        RECT 661.790 3429.430 663.010 3429.730 ;
        RECT 758.390 3429.730 758.690 3430.110 ;
        RECT 759.310 3429.730 759.610 3430.790 ;
        RECT 772.865 3430.775 773.195 3430.790 ;
        RECT 893.845 3431.090 894.175 3431.105 ;
        RECT 917.510 3431.090 917.890 3431.100 ;
        RECT 893.845 3430.790 917.890 3431.090 ;
        RECT 893.845 3430.775 894.175 3430.790 ;
        RECT 917.510 3430.780 917.890 3430.790 ;
        RECT 941.685 3431.090 942.015 3431.105 ;
        RECT 1449.065 3431.090 1449.395 3431.105 ;
        RECT 941.685 3430.790 1000.650 3431.090 ;
        RECT 941.685 3430.775 942.015 3430.790 ;
        RECT 1000.350 3430.410 1000.650 3430.790 ;
        RECT 1049.110 3430.790 1097.250 3431.090 ;
        RECT 1000.350 3430.110 1048.490 3430.410 ;
        RECT 758.390 3429.430 759.610 3429.730 ;
        RECT 811.045 3429.730 811.375 3429.745 ;
        RECT 820.910 3429.730 821.290 3429.740 ;
        RECT 811.045 3429.430 821.290 3429.730 ;
        RECT 1048.190 3429.730 1048.490 3430.110 ;
        RECT 1049.110 3429.730 1049.410 3430.790 ;
        RECT 1096.950 3430.410 1097.250 3430.790 ;
        RECT 1145.710 3430.790 1193.850 3431.090 ;
        RECT 1096.950 3430.110 1145.090 3430.410 ;
        RECT 1048.190 3429.430 1049.410 3429.730 ;
        RECT 1144.790 3429.730 1145.090 3430.110 ;
        RECT 1145.710 3429.730 1146.010 3430.790 ;
        RECT 1193.550 3430.410 1193.850 3430.790 ;
        RECT 1242.310 3430.790 1290.450 3431.090 ;
        RECT 1193.550 3430.110 1241.690 3430.410 ;
        RECT 1144.790 3429.430 1146.010 3429.730 ;
        RECT 1241.390 3429.730 1241.690 3430.110 ;
        RECT 1242.310 3429.730 1242.610 3430.790 ;
        RECT 1290.150 3430.410 1290.450 3430.790 ;
        RECT 1338.910 3430.790 1387.050 3431.090 ;
        RECT 1290.150 3430.110 1338.290 3430.410 ;
        RECT 1241.390 3429.430 1242.610 3429.730 ;
        RECT 1337.990 3429.730 1338.290 3430.110 ;
        RECT 1338.910 3429.730 1339.210 3430.790 ;
        RECT 1386.750 3430.410 1387.050 3430.790 ;
        RECT 1435.510 3430.790 1449.395 3431.090 ;
        RECT 1386.750 3430.110 1434.890 3430.410 ;
        RECT 1337.990 3429.430 1339.210 3429.730 ;
        RECT 1434.590 3429.730 1434.890 3430.110 ;
        RECT 1435.510 3429.730 1435.810 3430.790 ;
        RECT 1449.065 3430.775 1449.395 3430.790 ;
        RECT 1497.110 3431.090 1497.490 3431.100 ;
        RECT 1738.865 3431.090 1739.195 3431.105 ;
        RECT 1497.110 3430.790 1580.250 3431.090 ;
        RECT 1497.110 3430.780 1497.490 3430.790 ;
        RECT 1579.950 3430.410 1580.250 3430.790 ;
        RECT 1628.710 3430.790 1676.850 3431.090 ;
        RECT 1579.950 3430.110 1628.090 3430.410 ;
        RECT 1434.590 3429.430 1435.810 3429.730 ;
        RECT 1472.525 3429.730 1472.855 3429.745 ;
        RECT 1497.110 3429.730 1497.490 3429.740 ;
        RECT 1472.525 3429.430 1497.490 3429.730 ;
        RECT 1627.790 3429.730 1628.090 3430.110 ;
        RECT 1628.710 3429.730 1629.010 3430.790 ;
        RECT 1676.550 3430.410 1676.850 3430.790 ;
        RECT 1725.310 3430.790 1739.195 3431.090 ;
        RECT 1676.550 3430.110 1724.690 3430.410 ;
        RECT 1627.790 3429.430 1629.010 3429.730 ;
        RECT 1724.390 3429.730 1724.690 3430.110 ;
        RECT 1725.310 3429.730 1725.610 3430.790 ;
        RECT 1738.865 3430.775 1739.195 3430.790 ;
        RECT 1859.845 3431.090 1860.175 3431.105 ;
        RECT 1883.510 3431.090 1883.890 3431.100 ;
        RECT 1859.845 3430.790 1883.890 3431.090 ;
        RECT 1859.845 3430.775 1860.175 3430.790 ;
        RECT 1883.510 3430.780 1883.890 3430.790 ;
        RECT 1897.565 3431.090 1897.895 3431.105 ;
        RECT 2137.685 3431.090 2138.015 3431.105 ;
        RECT 1897.565 3430.790 1966.650 3431.090 ;
        RECT 1897.565 3430.775 1897.895 3430.790 ;
        RECT 1966.350 3430.410 1966.650 3430.790 ;
        RECT 2015.110 3430.790 2138.015 3431.090 ;
        RECT 1966.350 3430.110 2014.490 3430.410 ;
        RECT 1724.390 3429.430 1725.610 3429.730 ;
        RECT 1777.045 3429.730 1777.375 3429.745 ;
        RECT 1786.910 3429.730 1787.290 3429.740 ;
        RECT 1777.045 3429.430 1787.290 3429.730 ;
        RECT 2014.190 3429.730 2014.490 3430.110 ;
        RECT 2015.110 3429.730 2015.410 3430.790 ;
        RECT 2137.685 3430.775 2138.015 3430.790 ;
        RECT 2138.605 3431.090 2138.935 3431.105 ;
        RECT 2207.605 3431.090 2207.935 3431.105 ;
        RECT 2704.865 3431.090 2705.195 3431.105 ;
        RECT 2138.605 3430.790 2148.810 3431.090 ;
        RECT 2138.605 3430.775 2138.935 3430.790 ;
        RECT 2148.510 3430.410 2148.810 3430.790 ;
        RECT 2207.605 3430.790 2256.450 3431.090 ;
        RECT 2207.605 3430.775 2207.935 3430.790 ;
        RECT 2173.310 3430.410 2173.690 3430.420 ;
        RECT 2148.510 3430.110 2173.690 3430.410 ;
        RECT 2256.150 3430.410 2256.450 3430.790 ;
        RECT 2304.910 3430.790 2353.050 3431.090 ;
        RECT 2256.150 3430.110 2304.290 3430.410 ;
        RECT 2173.310 3430.100 2173.690 3430.110 ;
        RECT 2014.190 3429.430 2015.410 3429.730 ;
        RECT 2303.990 3429.730 2304.290 3430.110 ;
        RECT 2304.910 3429.730 2305.210 3430.790 ;
        RECT 2352.750 3430.410 2353.050 3430.790 ;
        RECT 2401.510 3430.790 2449.650 3431.090 ;
        RECT 2352.750 3430.110 2400.890 3430.410 ;
        RECT 2303.990 3429.430 2305.210 3429.730 ;
        RECT 2400.590 3429.730 2400.890 3430.110 ;
        RECT 2401.510 3429.730 2401.810 3430.790 ;
        RECT 2449.350 3430.410 2449.650 3430.790 ;
        RECT 2498.110 3430.790 2546.250 3431.090 ;
        RECT 2449.350 3430.110 2497.490 3430.410 ;
        RECT 2400.590 3429.430 2401.810 3429.730 ;
        RECT 2497.190 3429.730 2497.490 3430.110 ;
        RECT 2498.110 3429.730 2498.410 3430.790 ;
        RECT 2545.950 3430.410 2546.250 3430.790 ;
        RECT 2594.710 3430.790 2642.850 3431.090 ;
        RECT 2545.950 3430.110 2594.090 3430.410 ;
        RECT 2497.190 3429.430 2498.410 3429.730 ;
        RECT 2593.790 3429.730 2594.090 3430.110 ;
        RECT 2594.710 3429.730 2595.010 3430.790 ;
        RECT 2642.550 3430.410 2642.850 3430.790 ;
        RECT 2691.310 3430.790 2705.195 3431.090 ;
        RECT 2642.550 3430.110 2690.690 3430.410 ;
        RECT 2593.790 3429.430 2595.010 3429.730 ;
        RECT 2690.390 3429.730 2690.690 3430.110 ;
        RECT 2691.310 3429.730 2691.610 3430.790 ;
        RECT 2704.865 3430.775 2705.195 3430.790 ;
        RECT 2825.845 3431.090 2826.175 3431.105 ;
        RECT 2863.565 3431.090 2863.895 3431.105 ;
        RECT 2825.845 3430.790 2849.850 3431.090 ;
        RECT 2825.845 3430.775 2826.175 3430.790 ;
        RECT 2849.550 3430.410 2849.850 3430.790 ;
        RECT 2863.565 3430.790 2884.810 3431.090 ;
        RECT 2863.565 3430.775 2863.895 3430.790 ;
        RECT 2863.105 3430.410 2863.435 3430.425 ;
        RECT 2849.550 3430.110 2863.435 3430.410 ;
        RECT 2884.510 3430.410 2884.810 3430.790 ;
        RECT 2916.710 3430.410 2917.010 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2884.510 3430.110 2917.010 3430.410 ;
        RECT 2863.105 3430.095 2863.435 3430.110 ;
        RECT 2690.390 3429.430 2691.610 3429.730 ;
        RECT 2743.045 3429.730 2743.375 3429.745 ;
        RECT 2752.910 3429.730 2753.290 3429.740 ;
        RECT 2743.045 3429.430 2753.290 3429.730 ;
        RECT 811.045 3429.415 811.375 3429.430 ;
        RECT 820.910 3429.420 821.290 3429.430 ;
        RECT 1472.525 3429.415 1472.855 3429.430 ;
        RECT 1497.110 3429.420 1497.490 3429.430 ;
        RECT 1777.045 3429.415 1777.375 3429.430 ;
        RECT 1786.910 3429.420 1787.290 3429.430 ;
        RECT 2743.045 3429.415 2743.375 3429.430 ;
        RECT 2752.910 3429.420 2753.290 3429.430 ;
        RECT 288.230 2029.610 288.610 2029.620 ;
        RECT 300.000 2029.610 304.000 2029.720 ;
        RECT 288.230 2029.310 304.000 2029.610 ;
        RECT 288.230 2029.300 288.610 2029.310 ;
        RECT 300.000 2029.120 304.000 2029.310 ;
      LAYER via3 ;
        RECT 917.540 3432.140 917.860 3432.460 ;
        RECT 1883.540 3432.140 1883.860 3432.460 ;
        RECT 2173.340 3432.140 2173.660 3432.460 ;
        RECT 820.940 3431.460 821.260 3431.780 ;
        RECT 1786.940 3431.460 1787.260 3431.780 ;
        RECT 2752.940 3431.460 2753.260 3431.780 ;
        RECT 288.260 3430.780 288.580 3431.100 ;
        RECT 917.540 3430.780 917.860 3431.100 ;
        RECT 820.940 3429.420 821.260 3429.740 ;
        RECT 1497.140 3430.780 1497.460 3431.100 ;
        RECT 1497.140 3429.420 1497.460 3429.740 ;
        RECT 1883.540 3430.780 1883.860 3431.100 ;
        RECT 1786.940 3429.420 1787.260 3429.740 ;
        RECT 2173.340 3430.100 2173.660 3430.420 ;
        RECT 2752.940 3429.420 2753.260 3429.740 ;
        RECT 288.260 2029.300 288.580 2029.620 ;
      LAYER met4 ;
        RECT 917.535 3432.135 917.865 3432.465 ;
        RECT 1883.535 3432.135 1883.865 3432.465 ;
        RECT 2173.335 3432.135 2173.665 3432.465 ;
        RECT 820.935 3431.455 821.265 3431.785 ;
        RECT 288.255 3430.775 288.585 3431.105 ;
        RECT 288.270 2029.625 288.570 3430.775 ;
        RECT 820.950 3429.745 821.250 3431.455 ;
        RECT 917.550 3431.105 917.850 3432.135 ;
        RECT 1786.935 3431.455 1787.265 3431.785 ;
        RECT 917.535 3430.775 917.865 3431.105 ;
        RECT 1497.135 3430.775 1497.465 3431.105 ;
        RECT 1497.150 3429.745 1497.450 3430.775 ;
        RECT 1786.950 3429.745 1787.250 3431.455 ;
        RECT 1883.550 3431.105 1883.850 3432.135 ;
        RECT 1883.535 3430.775 1883.865 3431.105 ;
        RECT 2173.350 3430.425 2173.650 3432.135 ;
        RECT 2752.935 3431.455 2753.265 3431.785 ;
        RECT 2173.335 3430.095 2173.665 3430.425 ;
        RECT 2752.950 3429.745 2753.250 3431.455 ;
        RECT 820.935 3429.415 821.265 3429.745 ;
        RECT 1497.135 3429.415 1497.465 3429.745 ;
        RECT 1786.935 3429.415 1787.265 3429.745 ;
        RECT 2752.935 3429.415 2753.265 3429.745 ;
        RECT 288.255 2029.295 288.585 2029.625 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.845 2717.520 3517.600 ;
        RECT 2717.310 3501.475 2717.590 3501.845 ;
      LAYER via2 ;
        RECT 2717.310 3501.520 2717.590 3501.800 ;
      LAYER met3 ;
        RECT 289.150 3501.810 289.530 3501.820 ;
        RECT 2717.285 3501.810 2717.615 3501.825 ;
        RECT 289.150 3501.510 2717.615 3501.810 ;
        RECT 289.150 3501.500 289.530 3501.510 ;
        RECT 2717.285 3501.495 2717.615 3501.510 ;
        RECT 289.150 2058.850 289.530 2058.860 ;
        RECT 300.000 2058.850 304.000 2058.960 ;
        RECT 289.150 2058.550 304.000 2058.850 ;
        RECT 289.150 2058.540 289.530 2058.550 ;
        RECT 300.000 2058.360 304.000 2058.550 ;
      LAYER via3 ;
        RECT 289.180 3501.500 289.500 3501.820 ;
        RECT 289.180 2058.540 289.500 2058.860 ;
      LAYER met4 ;
        RECT 289.175 3501.495 289.505 3501.825 ;
        RECT 289.190 2058.865 289.490 3501.495 ;
        RECT 289.175 2058.535 289.505 2058.865 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 296.310 3501.900 296.630 3501.960 ;
        RECT 2392.530 3501.900 2392.850 3501.960 ;
        RECT 296.310 3501.760 2392.850 3501.900 ;
        RECT 296.310 3501.700 296.630 3501.760 ;
        RECT 2392.530 3501.700 2392.850 3501.760 ;
      LAYER via ;
        RECT 296.340 3501.700 296.600 3501.960 ;
        RECT 2392.560 3501.700 2392.820 3501.960 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3501.990 2392.760 3517.600 ;
        RECT 296.340 3501.670 296.600 3501.990 ;
        RECT 2392.560 3501.670 2392.820 3501.990 ;
        RECT 296.400 2087.445 296.540 3501.670 ;
        RECT 296.330 2087.075 296.610 2087.445 ;
      LAYER via2 ;
        RECT 296.330 2087.120 296.610 2087.400 ;
      LAYER met3 ;
        RECT 296.305 2087.410 296.635 2087.425 ;
        RECT 300.000 2087.410 304.000 2087.520 ;
        RECT 296.305 2087.110 304.000 2087.410 ;
        RECT 296.305 2087.095 296.635 2087.110 ;
        RECT 300.000 2086.920 304.000 2087.110 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 295.390 3502.240 295.710 3502.300 ;
        RECT 2068.230 3502.240 2068.550 3502.300 ;
        RECT 295.390 3502.100 2068.550 3502.240 ;
        RECT 295.390 3502.040 295.710 3502.100 ;
        RECT 2068.230 3502.040 2068.550 3502.100 ;
      LAYER via ;
        RECT 295.420 3502.040 295.680 3502.300 ;
        RECT 2068.260 3502.040 2068.520 3502.300 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3502.330 2068.460 3517.600 ;
        RECT 295.420 3502.010 295.680 3502.330 ;
        RECT 2068.260 3502.010 2068.520 3502.330 ;
        RECT 295.480 2116.685 295.620 3502.010 ;
        RECT 295.410 2116.315 295.690 2116.685 ;
      LAYER via2 ;
        RECT 295.410 2116.360 295.690 2116.640 ;
      LAYER met3 ;
        RECT 295.385 2116.650 295.715 2116.665 ;
        RECT 300.000 2116.650 304.000 2116.760 ;
        RECT 295.385 2116.350 304.000 2116.650 ;
        RECT 295.385 2116.335 295.715 2116.350 ;
        RECT 300.000 2116.160 304.000 2116.350 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 3502.920 289.730 3502.980 ;
        RECT 1743.930 3502.920 1744.250 3502.980 ;
        RECT 289.410 3502.780 1744.250 3502.920 ;
        RECT 289.410 3502.720 289.730 3502.780 ;
        RECT 1743.930 3502.720 1744.250 3502.780 ;
      LAYER via ;
        RECT 289.440 3502.720 289.700 3502.980 ;
        RECT 1743.960 3502.720 1744.220 3502.980 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3503.010 1744.160 3517.600 ;
        RECT 289.440 3502.690 289.700 3503.010 ;
        RECT 1743.960 3502.690 1744.220 3503.010 ;
        RECT 289.500 2145.245 289.640 3502.690 ;
        RECT 289.430 2144.875 289.710 2145.245 ;
      LAYER via2 ;
        RECT 289.430 2144.920 289.710 2145.200 ;
      LAYER met3 ;
        RECT 289.405 2145.210 289.735 2145.225 ;
        RECT 300.000 2145.210 304.000 2145.320 ;
        RECT 289.405 2144.910 304.000 2145.210 ;
        RECT 289.405 2144.895 289.735 2144.910 ;
        RECT 300.000 2144.720 304.000 2144.910 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 294.010 3503.600 294.330 3503.660 ;
        RECT 1419.170 3503.600 1419.490 3503.660 ;
        RECT 294.010 3503.460 1419.490 3503.600 ;
        RECT 294.010 3503.400 294.330 3503.460 ;
        RECT 1419.170 3503.400 1419.490 3503.460 ;
      LAYER via ;
        RECT 294.040 3503.400 294.300 3503.660 ;
        RECT 1419.200 3503.400 1419.460 3503.660 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3503.690 1419.400 3517.600 ;
        RECT 294.040 3503.370 294.300 3503.690 ;
        RECT 1419.200 3503.370 1419.460 3503.690 ;
        RECT 294.100 2174.485 294.240 3503.370 ;
        RECT 294.030 2174.115 294.310 2174.485 ;
      LAYER via2 ;
        RECT 294.030 2174.160 294.310 2174.440 ;
      LAYER met3 ;
        RECT 294.005 2174.450 294.335 2174.465 ;
        RECT 300.000 2174.450 304.000 2174.560 ;
        RECT 294.005 2174.150 304.000 2174.450 ;
        RECT 294.005 2174.135 294.335 2174.150 ;
        RECT 300.000 2173.960 304.000 2174.150 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.110 380.700 448.430 380.760 ;
        RECT 458.690 380.700 459.010 380.760 ;
        RECT 448.110 380.560 459.010 380.700 ;
        RECT 448.110 380.500 448.430 380.560 ;
        RECT 458.690 380.500 459.010 380.560 ;
        RECT 737.910 380.700 738.230 380.760 ;
        RECT 772.410 380.700 772.730 380.760 ;
        RECT 737.910 380.560 772.730 380.700 ;
        RECT 737.910 380.500 738.230 380.560 ;
        RECT 772.410 380.500 772.730 380.560 ;
        RECT 579.670 380.020 579.990 380.080 ;
        RECT 593.930 380.020 594.250 380.080 ;
        RECT 579.670 379.880 594.250 380.020 ;
        RECT 579.670 379.820 579.990 379.880 ;
        RECT 593.930 379.820 594.250 379.880 ;
      LAYER via ;
        RECT 448.140 380.500 448.400 380.760 ;
        RECT 458.720 380.500 458.980 380.760 ;
        RECT 737.940 380.500 738.200 380.760 ;
        RECT 772.440 380.500 772.700 380.760 ;
        RECT 579.700 379.820 579.960 380.080 ;
        RECT 593.960 379.820 594.220 380.080 ;
      LAYER met2 ;
        RECT 675.830 382.315 676.110 382.685 ;
        RECT 386.030 380.955 386.310 381.325 ;
        RECT 593.950 380.955 594.230 381.325 ;
        RECT 386.100 380.645 386.240 380.955 ;
        RECT 448.140 380.645 448.400 380.790 ;
        RECT 458.720 380.645 458.980 380.790 ;
        RECT 386.030 380.275 386.310 380.645 ;
        RECT 448.130 380.275 448.410 380.645 ;
        RECT 458.710 380.275 458.990 380.645 ;
        RECT 594.020 380.110 594.160 380.955 ;
        RECT 675.900 380.645 676.040 382.315 ;
        RECT 700.210 381.635 700.490 382.005 ;
        RECT 675.830 380.275 676.110 380.645 ;
        RECT 579.700 379.965 579.960 380.110 ;
        RECT 579.690 379.595 579.970 379.965 ;
        RECT 593.960 379.790 594.220 380.110 ;
        RECT 700.280 379.965 700.420 381.635 ;
        RECT 772.430 380.955 772.710 381.325 ;
        RECT 772.500 380.790 772.640 380.955 ;
        RECT 737.940 380.645 738.200 380.790 ;
        RECT 737.930 380.275 738.210 380.645 ;
        RECT 772.440 380.470 772.700 380.790 ;
        RECT 700.210 379.595 700.490 379.965 ;
      LAYER via2 ;
        RECT 675.830 382.360 676.110 382.640 ;
        RECT 386.030 381.000 386.310 381.280 ;
        RECT 593.950 381.000 594.230 381.280 ;
        RECT 386.030 380.320 386.310 380.600 ;
        RECT 448.130 380.320 448.410 380.600 ;
        RECT 458.710 380.320 458.990 380.600 ;
        RECT 700.210 381.680 700.490 381.960 ;
        RECT 675.830 380.320 676.110 380.600 ;
        RECT 579.690 379.640 579.970 379.920 ;
        RECT 772.430 381.000 772.710 381.280 ;
        RECT 737.930 380.320 738.210 380.600 ;
        RECT 700.210 379.640 700.490 379.920 ;
      LAYER met3 ;
        RECT 289.150 1652.890 289.530 1652.900 ;
        RECT 300.000 1652.890 304.000 1653.000 ;
        RECT 289.150 1652.590 304.000 1652.890 ;
        RECT 289.150 1652.580 289.530 1652.590 ;
        RECT 300.000 1652.400 304.000 1652.590 ;
        RECT 627.710 382.650 628.090 382.660 ;
        RECT 675.805 382.650 676.135 382.665 ;
        RECT 627.710 382.350 676.135 382.650 ;
        RECT 627.710 382.340 628.090 382.350 ;
        RECT 675.805 382.335 676.135 382.350 ;
        RECT 700.185 381.970 700.515 381.985 ;
        RECT 676.510 381.670 700.515 381.970 ;
        RECT 289.150 381.290 289.530 381.300 ;
        RECT 386.005 381.290 386.335 381.305 ;
        RECT 593.925 381.290 594.255 381.305 ;
        RECT 627.710 381.290 628.090 381.300 ;
        RECT 289.150 380.990 304.210 381.290 ;
        RECT 289.150 380.980 289.530 380.990 ;
        RECT 303.910 380.610 304.210 380.990 ;
        RECT 386.005 380.990 400.810 381.290 ;
        RECT 386.005 380.975 386.335 380.990 ;
        RECT 386.005 380.610 386.335 380.625 ;
        RECT 303.910 380.310 386.335 380.610 ;
        RECT 400.510 380.610 400.810 380.990 ;
        RECT 482.390 380.990 545.250 381.290 ;
        RECT 448.105 380.610 448.435 380.625 ;
        RECT 400.510 380.310 448.435 380.610 ;
        RECT 386.005 380.295 386.335 380.310 ;
        RECT 448.105 380.295 448.435 380.310 ;
        RECT 458.685 380.610 459.015 380.625 ;
        RECT 482.390 380.610 482.690 380.990 ;
        RECT 458.685 380.310 482.690 380.610 ;
        RECT 458.685 380.295 459.015 380.310 ;
        RECT 544.950 379.930 545.250 380.990 ;
        RECT 593.925 380.990 628.090 381.290 ;
        RECT 593.925 380.975 594.255 380.990 ;
        RECT 627.710 380.980 628.090 380.990 ;
        RECT 675.805 380.610 676.135 380.625 ;
        RECT 676.510 380.610 676.810 381.670 ;
        RECT 700.185 381.655 700.515 381.670 ;
        RECT 772.405 381.290 772.735 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 772.405 380.990 807.450 381.290 ;
        RECT 772.405 380.975 772.735 380.990 ;
        RECT 737.905 380.610 738.235 380.625 ;
        RECT 675.805 380.310 676.810 380.610 ;
        RECT 724.350 380.310 738.235 380.610 ;
        RECT 807.150 380.610 807.450 380.990 ;
        RECT 855.910 380.990 904.050 381.290 ;
        RECT 807.150 380.310 855.290 380.610 ;
        RECT 675.805 380.295 676.135 380.310 ;
        RECT 579.665 379.930 579.995 379.945 ;
        RECT 544.950 379.630 579.995 379.930 ;
        RECT 579.665 379.615 579.995 379.630 ;
        RECT 700.185 379.930 700.515 379.945 ;
        RECT 724.350 379.930 724.650 380.310 ;
        RECT 737.905 380.295 738.235 380.310 ;
        RECT 700.185 379.630 724.650 379.930 ;
        RECT 854.990 379.930 855.290 380.310 ;
        RECT 855.910 379.930 856.210 380.990 ;
        RECT 903.750 380.610 904.050 380.990 ;
        RECT 952.510 380.990 1000.650 381.290 ;
        RECT 903.750 380.310 951.890 380.610 ;
        RECT 854.990 379.630 856.210 379.930 ;
        RECT 951.590 379.930 951.890 380.310 ;
        RECT 952.510 379.930 952.810 380.990 ;
        RECT 1000.350 380.610 1000.650 380.990 ;
        RECT 1049.110 380.990 1097.250 381.290 ;
        RECT 1000.350 380.310 1048.490 380.610 ;
        RECT 951.590 379.630 952.810 379.930 ;
        RECT 1048.190 379.930 1048.490 380.310 ;
        RECT 1049.110 379.930 1049.410 380.990 ;
        RECT 1096.950 380.610 1097.250 380.990 ;
        RECT 1145.710 380.990 1193.850 381.290 ;
        RECT 1096.950 380.310 1145.090 380.610 ;
        RECT 1048.190 379.630 1049.410 379.930 ;
        RECT 1144.790 379.930 1145.090 380.310 ;
        RECT 1145.710 379.930 1146.010 380.990 ;
        RECT 1193.550 380.610 1193.850 380.990 ;
        RECT 1242.310 380.990 1290.450 381.290 ;
        RECT 1193.550 380.310 1241.690 380.610 ;
        RECT 1144.790 379.630 1146.010 379.930 ;
        RECT 1241.390 379.930 1241.690 380.310 ;
        RECT 1242.310 379.930 1242.610 380.990 ;
        RECT 1290.150 380.610 1290.450 380.990 ;
        RECT 1338.910 380.990 1387.050 381.290 ;
        RECT 1290.150 380.310 1338.290 380.610 ;
        RECT 1241.390 379.630 1242.610 379.930 ;
        RECT 1337.990 379.930 1338.290 380.310 ;
        RECT 1338.910 379.930 1339.210 380.990 ;
        RECT 1386.750 380.610 1387.050 380.990 ;
        RECT 1435.510 380.990 1483.650 381.290 ;
        RECT 1386.750 380.310 1434.890 380.610 ;
        RECT 1337.990 379.630 1339.210 379.930 ;
        RECT 1434.590 379.930 1434.890 380.310 ;
        RECT 1435.510 379.930 1435.810 380.990 ;
        RECT 1483.350 380.610 1483.650 380.990 ;
        RECT 1532.110 380.990 1580.250 381.290 ;
        RECT 1483.350 380.310 1531.490 380.610 ;
        RECT 1434.590 379.630 1435.810 379.930 ;
        RECT 1531.190 379.930 1531.490 380.310 ;
        RECT 1532.110 379.930 1532.410 380.990 ;
        RECT 1579.950 380.610 1580.250 380.990 ;
        RECT 1628.710 380.990 1676.850 381.290 ;
        RECT 1579.950 380.310 1628.090 380.610 ;
        RECT 1531.190 379.630 1532.410 379.930 ;
        RECT 1627.790 379.930 1628.090 380.310 ;
        RECT 1628.710 379.930 1629.010 380.990 ;
        RECT 1676.550 380.610 1676.850 380.990 ;
        RECT 1725.310 380.990 1773.450 381.290 ;
        RECT 1676.550 380.310 1724.690 380.610 ;
        RECT 1627.790 379.630 1629.010 379.930 ;
        RECT 1724.390 379.930 1724.690 380.310 ;
        RECT 1725.310 379.930 1725.610 380.990 ;
        RECT 1773.150 380.610 1773.450 380.990 ;
        RECT 1821.910 380.990 1870.050 381.290 ;
        RECT 1773.150 380.310 1821.290 380.610 ;
        RECT 1724.390 379.630 1725.610 379.930 ;
        RECT 1820.990 379.930 1821.290 380.310 ;
        RECT 1821.910 379.930 1822.210 380.990 ;
        RECT 1869.750 380.610 1870.050 380.990 ;
        RECT 1918.510 380.990 1966.650 381.290 ;
        RECT 1869.750 380.310 1917.890 380.610 ;
        RECT 1820.990 379.630 1822.210 379.930 ;
        RECT 1917.590 379.930 1917.890 380.310 ;
        RECT 1918.510 379.930 1918.810 380.990 ;
        RECT 1966.350 380.610 1966.650 380.990 ;
        RECT 2015.110 380.990 2063.250 381.290 ;
        RECT 1966.350 380.310 2014.490 380.610 ;
        RECT 1917.590 379.630 1918.810 379.930 ;
        RECT 2014.190 379.930 2014.490 380.310 ;
        RECT 2015.110 379.930 2015.410 380.990 ;
        RECT 2062.950 380.610 2063.250 380.990 ;
        RECT 2111.710 380.990 2159.850 381.290 ;
        RECT 2062.950 380.310 2111.090 380.610 ;
        RECT 2014.190 379.630 2015.410 379.930 ;
        RECT 2110.790 379.930 2111.090 380.310 ;
        RECT 2111.710 379.930 2112.010 380.990 ;
        RECT 2159.550 380.610 2159.850 380.990 ;
        RECT 2208.310 380.990 2256.450 381.290 ;
        RECT 2159.550 380.310 2207.690 380.610 ;
        RECT 2110.790 379.630 2112.010 379.930 ;
        RECT 2207.390 379.930 2207.690 380.310 ;
        RECT 2208.310 379.930 2208.610 380.990 ;
        RECT 2256.150 380.610 2256.450 380.990 ;
        RECT 2304.910 380.990 2353.050 381.290 ;
        RECT 2256.150 380.310 2304.290 380.610 ;
        RECT 2207.390 379.630 2208.610 379.930 ;
        RECT 2303.990 379.930 2304.290 380.310 ;
        RECT 2304.910 379.930 2305.210 380.990 ;
        RECT 2352.750 380.610 2353.050 380.990 ;
        RECT 2401.510 380.990 2449.650 381.290 ;
        RECT 2352.750 380.310 2400.890 380.610 ;
        RECT 2303.990 379.630 2305.210 379.930 ;
        RECT 2400.590 379.930 2400.890 380.310 ;
        RECT 2401.510 379.930 2401.810 380.990 ;
        RECT 2449.350 380.610 2449.650 380.990 ;
        RECT 2498.110 380.990 2546.250 381.290 ;
        RECT 2449.350 380.310 2497.490 380.610 ;
        RECT 2400.590 379.630 2401.810 379.930 ;
        RECT 2497.190 379.930 2497.490 380.310 ;
        RECT 2498.110 379.930 2498.410 380.990 ;
        RECT 2545.950 380.610 2546.250 380.990 ;
        RECT 2594.710 380.990 2642.850 381.290 ;
        RECT 2545.950 380.310 2594.090 380.610 ;
        RECT 2497.190 379.630 2498.410 379.930 ;
        RECT 2593.790 379.930 2594.090 380.310 ;
        RECT 2594.710 379.930 2595.010 380.990 ;
        RECT 2642.550 380.610 2642.850 380.990 ;
        RECT 2691.310 380.990 2739.450 381.290 ;
        RECT 2642.550 380.310 2690.690 380.610 ;
        RECT 2593.790 379.630 2595.010 379.930 ;
        RECT 2690.390 379.930 2690.690 380.310 ;
        RECT 2691.310 379.930 2691.610 380.990 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2690.390 379.630 2691.610 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 700.185 379.615 700.515 379.630 ;
      LAYER via3 ;
        RECT 289.180 1652.580 289.500 1652.900 ;
        RECT 627.740 382.340 628.060 382.660 ;
        RECT 289.180 380.980 289.500 381.300 ;
        RECT 627.740 380.980 628.060 381.300 ;
      LAYER met4 ;
        RECT 289.175 1652.575 289.505 1652.905 ;
        RECT 289.190 381.305 289.490 1652.575 ;
        RECT 627.735 382.335 628.065 382.665 ;
        RECT 627.750 381.305 628.050 382.335 ;
        RECT 289.175 380.975 289.505 381.305 ;
        RECT 627.735 380.975 628.065 381.305 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 3504.280 289.270 3504.340 ;
        RECT 1094.870 3504.280 1095.190 3504.340 ;
        RECT 288.950 3504.140 1095.190 3504.280 ;
        RECT 288.950 3504.080 289.270 3504.140 ;
        RECT 1094.870 3504.080 1095.190 3504.140 ;
      LAYER via ;
        RECT 288.980 3504.080 289.240 3504.340 ;
        RECT 1094.900 3504.080 1095.160 3504.340 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3504.370 1095.100 3517.600 ;
        RECT 288.980 3504.050 289.240 3504.370 ;
        RECT 1094.900 3504.050 1095.160 3504.370 ;
        RECT 289.040 2203.045 289.180 3504.050 ;
        RECT 288.970 2202.675 289.250 2203.045 ;
      LAYER via2 ;
        RECT 288.970 2202.720 289.250 2203.000 ;
      LAYER met3 ;
        RECT 288.945 2203.010 289.275 2203.025 ;
        RECT 300.000 2203.010 304.000 2203.120 ;
        RECT 288.945 2202.710 304.000 2203.010 ;
        RECT 288.945 2202.695 289.275 2202.710 ;
        RECT 300.000 2202.520 304.000 2202.710 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 292.630 3501.220 292.950 3501.280 ;
        RECT 770.570 3501.220 770.890 3501.280 ;
        RECT 292.630 3501.080 770.890 3501.220 ;
        RECT 292.630 3501.020 292.950 3501.080 ;
        RECT 770.570 3501.020 770.890 3501.080 ;
      LAYER via ;
        RECT 292.660 3501.020 292.920 3501.280 ;
        RECT 770.600 3501.020 770.860 3501.280 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3501.310 770.800 3517.600 ;
        RECT 292.660 3500.990 292.920 3501.310 ;
        RECT 770.600 3500.990 770.860 3501.310 ;
        RECT 292.720 2232.285 292.860 3500.990 ;
        RECT 292.650 2231.915 292.930 2232.285 ;
      LAYER via2 ;
        RECT 292.650 2231.960 292.930 2232.240 ;
      LAYER met3 ;
        RECT 292.625 2232.250 292.955 2232.265 ;
        RECT 300.000 2232.250 304.000 2232.360 ;
        RECT 292.625 2231.950 304.000 2232.250 ;
        RECT 292.625 2231.935 292.955 2231.950 ;
        RECT 300.000 2231.760 304.000 2231.950 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 291.710 3500.880 292.030 3500.940 ;
        RECT 445.810 3500.880 446.130 3500.940 ;
        RECT 291.710 3500.740 446.130 3500.880 ;
        RECT 291.710 3500.680 292.030 3500.740 ;
        RECT 445.810 3500.680 446.130 3500.740 ;
      LAYER via ;
        RECT 291.740 3500.680 292.000 3500.940 ;
        RECT 445.840 3500.680 446.100 3500.940 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3500.970 446.040 3517.600 ;
        RECT 291.740 3500.650 292.000 3500.970 ;
        RECT 445.840 3500.650 446.100 3500.970 ;
        RECT 291.800 2261.525 291.940 3500.650 ;
        RECT 291.730 2261.155 292.010 2261.525 ;
      LAYER via2 ;
        RECT 291.730 2261.200 292.010 2261.480 ;
      LAYER met3 ;
        RECT 291.705 2261.490 292.035 2261.505 ;
        RECT 300.000 2261.490 304.000 2261.600 ;
        RECT 291.705 2261.190 304.000 2261.490 ;
        RECT 291.705 2261.175 292.035 2261.190 ;
        RECT 300.000 2261.000 304.000 2261.190 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 2290.820 124.130 2290.880 ;
        RECT 282.970 2290.820 283.290 2290.880 ;
        RECT 123.810 2290.680 283.290 2290.820 ;
        RECT 123.810 2290.620 124.130 2290.680 ;
        RECT 282.970 2290.620 283.290 2290.680 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 2290.620 124.100 2290.880 ;
        RECT 283.000 2290.620 283.260 2290.880 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 2290.910 124.040 3498.270 ;
        RECT 123.840 2290.590 124.100 2290.910 ;
        RECT 283.000 2290.590 283.260 2290.910 ;
        RECT 283.060 2290.085 283.200 2290.590 ;
        RECT 282.990 2289.715 283.270 2290.085 ;
      LAYER via2 ;
        RECT 282.990 2289.760 283.270 2290.040 ;
      LAYER met3 ;
        RECT 282.965 2290.050 283.295 2290.065 ;
        RECT 300.000 2290.050 304.000 2290.160 ;
        RECT 282.965 2289.750 304.000 2290.050 ;
        RECT 282.965 2289.735 283.295 2289.750 ;
        RECT 300.000 2289.560 304.000 2289.750 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 3339.720 17.870 3339.780 ;
        RECT 106.790 3339.720 107.110 3339.780 ;
        RECT 17.550 3339.580 107.110 3339.720 ;
        RECT 17.550 3339.520 17.870 3339.580 ;
        RECT 106.790 3339.520 107.110 3339.580 ;
        RECT 106.790 2325.160 107.110 2325.220 ;
        RECT 282.510 2325.160 282.830 2325.220 ;
        RECT 106.790 2325.020 282.830 2325.160 ;
        RECT 106.790 2324.960 107.110 2325.020 ;
        RECT 282.510 2324.960 282.830 2325.020 ;
      LAYER via ;
        RECT 17.580 3339.520 17.840 3339.780 ;
        RECT 106.820 3339.520 107.080 3339.780 ;
        RECT 106.820 2324.960 107.080 2325.220 ;
        RECT 282.540 2324.960 282.800 2325.220 ;
      LAYER met2 ;
        RECT 17.570 3339.635 17.850 3340.005 ;
        RECT 17.580 3339.490 17.840 3339.635 ;
        RECT 106.820 3339.490 107.080 3339.810 ;
        RECT 106.880 2325.250 107.020 3339.490 ;
        RECT 106.820 2324.930 107.080 2325.250 ;
        RECT 282.540 2324.930 282.800 2325.250 ;
        RECT 282.600 2319.325 282.740 2324.930 ;
        RECT 282.530 2318.955 282.810 2319.325 ;
      LAYER via2 ;
        RECT 17.570 3339.680 17.850 3339.960 ;
        RECT 282.530 2319.000 282.810 2319.280 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.545 3339.970 17.875 3339.985 ;
        RECT -4.800 3339.670 17.875 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.545 3339.655 17.875 3339.670 ;
        RECT 282.505 2319.290 282.835 2319.305 ;
        RECT 300.000 2319.290 304.000 2319.400 ;
        RECT 282.505 2318.990 304.000 2319.290 ;
        RECT 282.505 2318.975 282.835 2318.990 ;
        RECT 300.000 2318.800 304.000 2318.990 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 3050.040 18.330 3050.100 ;
        RECT 155.090 3050.040 155.410 3050.100 ;
        RECT 18.010 3049.900 155.410 3050.040 ;
        RECT 18.010 3049.840 18.330 3049.900 ;
        RECT 155.090 3049.840 155.410 3049.900 ;
        RECT 155.090 2352.700 155.410 2352.760 ;
        RECT 282.510 2352.700 282.830 2352.760 ;
        RECT 155.090 2352.560 282.830 2352.700 ;
        RECT 155.090 2352.500 155.410 2352.560 ;
        RECT 282.510 2352.500 282.830 2352.560 ;
      LAYER via ;
        RECT 18.040 3049.840 18.300 3050.100 ;
        RECT 155.120 3049.840 155.380 3050.100 ;
        RECT 155.120 2352.500 155.380 2352.760 ;
        RECT 282.540 2352.500 282.800 2352.760 ;
      LAYER met2 ;
        RECT 18.030 3051.995 18.310 3052.365 ;
        RECT 18.100 3050.130 18.240 3051.995 ;
        RECT 18.040 3049.810 18.300 3050.130 ;
        RECT 155.120 3049.810 155.380 3050.130 ;
        RECT 155.180 2352.790 155.320 3049.810 ;
        RECT 155.120 2352.470 155.380 2352.790 ;
        RECT 282.540 2352.470 282.800 2352.790 ;
        RECT 282.600 2347.885 282.740 2352.470 ;
        RECT 282.530 2347.515 282.810 2347.885 ;
      LAYER via2 ;
        RECT 18.030 3052.040 18.310 3052.320 ;
        RECT 282.530 2347.560 282.810 2347.840 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 18.005 3052.330 18.335 3052.345 ;
        RECT -4.800 3052.030 18.335 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 18.005 3052.015 18.335 3052.030 ;
        RECT 282.505 2347.850 282.835 2347.865 ;
        RECT 300.000 2347.850 304.000 2347.960 ;
        RECT 282.505 2347.550 304.000 2347.850 ;
        RECT 282.505 2347.535 282.835 2347.550 ;
        RECT 300.000 2347.360 304.000 2347.550 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2380.240 18.790 2380.300 ;
        RECT 282.510 2380.240 282.830 2380.300 ;
        RECT 18.470 2380.100 282.830 2380.240 ;
        RECT 18.470 2380.040 18.790 2380.100 ;
        RECT 282.510 2380.040 282.830 2380.100 ;
      LAYER via ;
        RECT 18.500 2380.040 18.760 2380.300 ;
        RECT 282.540 2380.040 282.800 2380.300 ;
      LAYER met2 ;
        RECT 18.490 2765.035 18.770 2765.405 ;
        RECT 18.560 2380.330 18.700 2765.035 ;
        RECT 18.500 2380.010 18.760 2380.330 ;
        RECT 282.540 2380.010 282.800 2380.330 ;
        RECT 282.600 2377.125 282.740 2380.010 ;
        RECT 282.530 2376.755 282.810 2377.125 ;
      LAYER via2 ;
        RECT 18.490 2765.080 18.770 2765.360 ;
        RECT 282.530 2376.800 282.810 2377.080 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.465 2765.370 18.795 2765.385 ;
        RECT -4.800 2765.070 18.795 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.465 2765.055 18.795 2765.070 ;
        RECT 282.505 2377.090 282.835 2377.105 ;
        RECT 300.000 2377.090 304.000 2377.200 ;
        RECT 282.505 2376.790 304.000 2377.090 ;
        RECT 282.505 2376.775 282.835 2376.790 ;
        RECT 300.000 2376.600 304.000 2376.790 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 2477.480 20.170 2477.540 ;
        RECT 25.830 2477.480 26.150 2477.540 ;
        RECT 19.850 2477.340 26.150 2477.480 ;
        RECT 19.850 2477.280 20.170 2477.340 ;
        RECT 25.830 2477.280 26.150 2477.340 ;
        RECT 25.830 2408.120 26.150 2408.180 ;
        RECT 283.430 2408.120 283.750 2408.180 ;
        RECT 25.830 2407.980 283.750 2408.120 ;
        RECT 25.830 2407.920 26.150 2407.980 ;
        RECT 283.430 2407.920 283.750 2407.980 ;
      LAYER via ;
        RECT 19.880 2477.280 20.140 2477.540 ;
        RECT 25.860 2477.280 26.120 2477.540 ;
        RECT 25.860 2407.920 26.120 2408.180 ;
        RECT 283.460 2407.920 283.720 2408.180 ;
      LAYER met2 ;
        RECT 19.870 2477.395 20.150 2477.765 ;
        RECT 19.880 2477.250 20.140 2477.395 ;
        RECT 25.860 2477.250 26.120 2477.570 ;
        RECT 25.920 2408.210 26.060 2477.250 ;
        RECT 25.860 2407.890 26.120 2408.210 ;
        RECT 283.460 2407.890 283.720 2408.210 ;
        RECT 283.520 2406.365 283.660 2407.890 ;
        RECT 283.450 2405.995 283.730 2406.365 ;
      LAYER via2 ;
        RECT 19.870 2477.440 20.150 2477.720 ;
        RECT 283.450 2406.040 283.730 2406.320 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 19.845 2477.730 20.175 2477.745 ;
        RECT -4.800 2477.430 20.175 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 19.845 2477.415 20.175 2477.430 ;
        RECT 283.425 2406.330 283.755 2406.345 ;
        RECT 300.000 2406.330 304.000 2406.440 ;
        RECT 283.425 2406.030 304.000 2406.330 ;
        RECT 283.425 2406.015 283.755 2406.030 ;
        RECT 300.000 2405.840 304.000 2406.030 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 2429.200 20.170 2429.260 ;
        RECT 283.430 2429.200 283.750 2429.260 ;
        RECT 19.850 2429.060 283.750 2429.200 ;
        RECT 19.850 2429.000 20.170 2429.060 ;
        RECT 283.430 2429.000 283.750 2429.060 ;
      LAYER via ;
        RECT 19.880 2429.000 20.140 2429.260 ;
        RECT 283.460 2429.000 283.720 2429.260 ;
      LAYER met2 ;
        RECT 283.450 2434.555 283.730 2434.925 ;
        RECT 283.520 2429.290 283.660 2434.555 ;
        RECT 19.880 2428.970 20.140 2429.290 ;
        RECT 283.460 2428.970 283.720 2429.290 ;
        RECT 19.940 2190.125 20.080 2428.970 ;
        RECT 19.870 2189.755 20.150 2190.125 ;
      LAYER via2 ;
        RECT 283.450 2434.600 283.730 2434.880 ;
        RECT 19.870 2189.800 20.150 2190.080 ;
      LAYER met3 ;
        RECT 283.425 2434.890 283.755 2434.905 ;
        RECT 300.000 2434.890 304.000 2435.000 ;
        RECT 283.425 2434.590 304.000 2434.890 ;
        RECT 283.425 2434.575 283.755 2434.590 ;
        RECT 300.000 2434.400 304.000 2434.590 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 19.845 2190.090 20.175 2190.105 ;
        RECT -4.800 2189.790 20.175 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 19.845 2189.775 20.175 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 285.270 1904.240 285.590 1904.300 ;
        RECT 16.170 1904.100 285.590 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 285.270 1904.040 285.590 1904.100 ;
      LAYER via ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 285.300 1904.040 285.560 1904.300 ;
      LAYER met2 ;
        RECT 285.290 2463.795 285.570 2464.165 ;
        RECT 285.360 1904.330 285.500 2463.795 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 285.300 1904.010 285.560 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 285.290 2463.840 285.570 2464.120 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 285.265 2464.130 285.595 2464.145 ;
        RECT 300.000 2464.130 304.000 2464.240 ;
        RECT 285.265 2463.830 304.000 2464.130 ;
        RECT 285.265 2463.815 285.595 2463.830 ;
        RECT 300.000 2463.640 304.000 2463.830 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.810 1646.860 285.130 1646.920 ;
        RECT 288.950 1646.860 289.270 1646.920 ;
        RECT 284.810 1646.720 289.270 1646.860 ;
        RECT 284.810 1646.660 285.130 1646.720 ;
        RECT 288.950 1646.660 289.270 1646.720 ;
        RECT 284.810 620.740 285.130 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 284.810 620.600 2901.150 620.740 ;
        RECT 284.810 620.540 285.130 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 284.840 1646.660 285.100 1646.920 ;
        RECT 288.980 1646.660 289.240 1646.920 ;
        RECT 284.840 620.540 285.100 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 288.970 1681.795 289.250 1682.165 ;
        RECT 289.040 1646.950 289.180 1681.795 ;
        RECT 284.840 1646.630 285.100 1646.950 ;
        RECT 288.980 1646.630 289.240 1646.950 ;
        RECT 284.900 620.830 285.040 1646.630 ;
        RECT 284.840 620.510 285.100 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 288.970 1681.840 289.250 1682.120 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 288.945 1682.130 289.275 1682.145 ;
        RECT 300.000 1682.130 304.000 1682.240 ;
        RECT 288.945 1681.830 304.000 1682.130 ;
        RECT 288.945 1681.815 289.275 1681.830 ;
        RECT 300.000 1681.640 304.000 1681.830 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 161.990 2491.080 162.310 2491.140 ;
        RECT 287.110 2491.080 287.430 2491.140 ;
        RECT 161.990 2490.940 287.430 2491.080 ;
        RECT 161.990 2490.880 162.310 2490.940 ;
        RECT 287.110 2490.880 287.430 2490.940 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 161.990 1621.360 162.310 1621.420 ;
        RECT 16.170 1621.220 162.310 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 161.990 1621.160 162.310 1621.220 ;
      LAYER via ;
        RECT 162.020 2490.880 162.280 2491.140 ;
        RECT 287.140 2490.880 287.400 2491.140 ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 162.020 1621.160 162.280 1621.420 ;
      LAYER met2 ;
        RECT 287.130 2492.355 287.410 2492.725 ;
        RECT 287.200 2491.170 287.340 2492.355 ;
        RECT 162.020 2490.850 162.280 2491.170 ;
        RECT 287.140 2490.850 287.400 2491.170 ;
        RECT 162.080 1621.450 162.220 2490.850 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 162.020 1621.130 162.280 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 287.130 2492.400 287.410 2492.680 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT 287.105 2492.690 287.435 2492.705 ;
        RECT 300.000 2492.690 304.000 2492.800 ;
        RECT 287.105 2492.390 304.000 2492.690 ;
        RECT 287.105 2492.375 287.435 2492.390 ;
        RECT 300.000 2492.200 304.000 2492.390 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 189.590 2518.620 189.910 2518.680 ;
        RECT 287.110 2518.620 287.430 2518.680 ;
        RECT 189.590 2518.480 287.430 2518.620 ;
        RECT 189.590 2518.420 189.910 2518.480 ;
        RECT 287.110 2518.420 287.430 2518.480 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 189.590 1400.700 189.910 1400.760 ;
        RECT 17.090 1400.560 189.910 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 189.590 1400.500 189.910 1400.560 ;
      LAYER via ;
        RECT 189.620 2518.420 189.880 2518.680 ;
        RECT 287.140 2518.420 287.400 2518.680 ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 189.620 1400.500 189.880 1400.760 ;
      LAYER met2 ;
        RECT 287.130 2521.595 287.410 2521.965 ;
        RECT 287.200 2518.710 287.340 2521.595 ;
        RECT 189.620 2518.390 189.880 2518.710 ;
        RECT 287.140 2518.390 287.400 2518.710 ;
        RECT 189.680 1400.790 189.820 2518.390 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 189.620 1400.470 189.880 1400.790 ;
      LAYER via2 ;
        RECT 287.130 2521.640 287.410 2521.920 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 287.105 2521.930 287.435 2521.945 ;
        RECT 300.000 2521.930 304.000 2522.040 ;
        RECT 287.105 2521.630 304.000 2521.930 ;
        RECT 287.105 2521.615 287.435 2521.630 ;
        RECT 300.000 2521.440 304.000 2521.630 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.950 2546.500 197.270 2546.560 ;
        RECT 287.110 2546.500 287.430 2546.560 ;
        RECT 196.950 2546.360 287.430 2546.500 ;
        RECT 196.950 2546.300 197.270 2546.360 ;
        RECT 287.110 2546.300 287.430 2546.360 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 196.950 1186.840 197.270 1186.900 ;
        RECT 17.090 1186.700 197.270 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 196.950 1186.640 197.270 1186.700 ;
      LAYER via ;
        RECT 196.980 2546.300 197.240 2546.560 ;
        RECT 287.140 2546.300 287.400 2546.560 ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 196.980 1186.640 197.240 1186.900 ;
      LAYER met2 ;
        RECT 287.130 2550.155 287.410 2550.525 ;
        RECT 287.200 2546.590 287.340 2550.155 ;
        RECT 196.980 2546.270 197.240 2546.590 ;
        RECT 287.140 2546.270 287.400 2546.590 ;
        RECT 197.040 1186.930 197.180 2546.270 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 196.980 1186.610 197.240 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 287.130 2550.200 287.410 2550.480 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 287.105 2550.490 287.435 2550.505 ;
        RECT 300.000 2550.490 304.000 2550.600 ;
        RECT 287.105 2550.190 304.000 2550.490 ;
        RECT 287.105 2550.175 287.435 2550.190 ;
        RECT 300.000 2550.000 304.000 2550.190 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 251.690 2574.040 252.010 2574.100 ;
        RECT 287.110 2574.040 287.430 2574.100 ;
        RECT 251.690 2573.900 287.430 2574.040 ;
        RECT 251.690 2573.840 252.010 2573.900 ;
        RECT 287.110 2573.840 287.430 2573.900 ;
        RECT 14.330 972.640 14.650 972.700 ;
        RECT 251.690 972.640 252.010 972.700 ;
        RECT 14.330 972.500 252.010 972.640 ;
        RECT 14.330 972.440 14.650 972.500 ;
        RECT 251.690 972.440 252.010 972.500 ;
      LAYER via ;
        RECT 251.720 2573.840 251.980 2574.100 ;
        RECT 287.140 2573.840 287.400 2574.100 ;
        RECT 14.360 972.440 14.620 972.700 ;
        RECT 251.720 972.440 251.980 972.700 ;
      LAYER met2 ;
        RECT 287.130 2579.395 287.410 2579.765 ;
        RECT 287.200 2574.130 287.340 2579.395 ;
        RECT 251.720 2573.810 251.980 2574.130 ;
        RECT 287.140 2573.810 287.400 2574.130 ;
        RECT 251.780 972.730 251.920 2573.810 ;
        RECT 14.360 972.410 14.620 972.730 ;
        RECT 251.720 972.410 251.980 972.730 ;
        RECT 14.420 969.525 14.560 972.410 ;
        RECT 14.350 969.155 14.630 969.525 ;
      LAYER via2 ;
        RECT 287.130 2579.440 287.410 2579.720 ;
        RECT 14.350 969.200 14.630 969.480 ;
      LAYER met3 ;
        RECT 287.105 2579.730 287.435 2579.745 ;
        RECT 300.000 2579.730 304.000 2579.840 ;
        RECT 287.105 2579.430 304.000 2579.730 ;
        RECT 287.105 2579.415 287.435 2579.430 ;
        RECT 300.000 2579.240 304.000 2579.430 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 14.325 969.490 14.655 969.505 ;
        RECT -4.800 969.190 14.655 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 14.325 969.175 14.655 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 258.590 2608.720 258.910 2608.780 ;
        RECT 287.110 2608.720 287.430 2608.780 ;
        RECT 258.590 2608.580 287.430 2608.720 ;
        RECT 258.590 2608.520 258.910 2608.580 ;
        RECT 287.110 2608.520 287.430 2608.580 ;
        RECT 15.710 758.780 16.030 758.840 ;
        RECT 258.590 758.780 258.910 758.840 ;
        RECT 15.710 758.640 258.910 758.780 ;
        RECT 15.710 758.580 16.030 758.640 ;
        RECT 258.590 758.580 258.910 758.640 ;
      LAYER via ;
        RECT 258.620 2608.520 258.880 2608.780 ;
        RECT 287.140 2608.520 287.400 2608.780 ;
        RECT 15.740 758.580 16.000 758.840 ;
        RECT 258.620 758.580 258.880 758.840 ;
      LAYER met2 ;
        RECT 258.620 2608.490 258.880 2608.810 ;
        RECT 287.130 2608.635 287.410 2609.005 ;
        RECT 287.140 2608.490 287.400 2608.635 ;
        RECT 258.680 758.870 258.820 2608.490 ;
        RECT 15.740 758.550 16.000 758.870 ;
        RECT 258.620 758.550 258.880 758.870 ;
        RECT 15.800 753.965 15.940 758.550 ;
        RECT 15.730 753.595 16.010 753.965 ;
      LAYER via2 ;
        RECT 287.130 2608.680 287.410 2608.960 ;
        RECT 15.730 753.640 16.010 753.920 ;
      LAYER met3 ;
        RECT 287.105 2608.970 287.435 2608.985 ;
        RECT 300.000 2608.970 304.000 2609.080 ;
        RECT 287.105 2608.670 304.000 2608.970 ;
        RECT 287.105 2608.655 287.435 2608.670 ;
        RECT 300.000 2608.480 304.000 2608.670 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 15.705 753.930 16.035 753.945 ;
        RECT -4.800 753.630 16.035 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 15.705 753.615 16.035 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 265.490 2635.920 265.810 2635.980 ;
        RECT 287.110 2635.920 287.430 2635.980 ;
        RECT 265.490 2635.780 287.430 2635.920 ;
        RECT 265.490 2635.720 265.810 2635.780 ;
        RECT 287.110 2635.720 287.430 2635.780 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 265.490 544.920 265.810 544.980 ;
        RECT 16.170 544.780 265.810 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 265.490 544.720 265.810 544.780 ;
      LAYER via ;
        RECT 265.520 2635.720 265.780 2635.980 ;
        RECT 287.140 2635.720 287.400 2635.980 ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 265.520 544.720 265.780 544.980 ;
      LAYER met2 ;
        RECT 287.130 2637.195 287.410 2637.565 ;
        RECT 287.200 2636.010 287.340 2637.195 ;
        RECT 265.520 2635.690 265.780 2636.010 ;
        RECT 287.140 2635.690 287.400 2636.010 ;
        RECT 265.580 545.010 265.720 2635.690 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 265.520 544.690 265.780 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 287.130 2637.240 287.410 2637.520 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 287.105 2637.530 287.435 2637.545 ;
        RECT 300.000 2637.530 304.000 2637.640 ;
        RECT 287.105 2637.230 304.000 2637.530 ;
        RECT 287.105 2637.215 287.435 2637.230 ;
        RECT 300.000 2637.040 304.000 2637.230 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 141.290 2663.800 141.610 2663.860 ;
        RECT 287.110 2663.800 287.430 2663.860 ;
        RECT 141.290 2663.660 287.430 2663.800 ;
        RECT 141.290 2663.600 141.610 2663.660 ;
        RECT 287.110 2663.600 287.430 2663.660 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 141.290 324.260 141.610 324.320 ;
        RECT 16.630 324.120 141.610 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 141.290 324.060 141.610 324.120 ;
      LAYER via ;
        RECT 141.320 2663.600 141.580 2663.860 ;
        RECT 287.140 2663.600 287.400 2663.860 ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 141.320 324.060 141.580 324.320 ;
      LAYER met2 ;
        RECT 287.130 2666.435 287.410 2666.805 ;
        RECT 287.200 2663.890 287.340 2666.435 ;
        RECT 141.320 2663.570 141.580 2663.890 ;
        RECT 287.140 2663.570 287.400 2663.890 ;
        RECT 141.380 324.350 141.520 2663.570 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 141.320 324.030 141.580 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 287.130 2666.480 287.410 2666.760 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 287.105 2666.770 287.435 2666.785 ;
        RECT 300.000 2666.770 304.000 2666.880 ;
        RECT 287.105 2666.470 304.000 2666.770 ;
        RECT 287.105 2666.455 287.435 2666.470 ;
        RECT 300.000 2666.280 304.000 2666.470 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 168.890 2691.340 169.210 2691.400 ;
        RECT 287.110 2691.340 287.430 2691.400 ;
        RECT 168.890 2691.200 287.430 2691.340 ;
        RECT 168.890 2691.140 169.210 2691.200 ;
        RECT 287.110 2691.140 287.430 2691.200 ;
        RECT 14.330 110.400 14.650 110.460 ;
        RECT 168.890 110.400 169.210 110.460 ;
        RECT 14.330 110.260 169.210 110.400 ;
        RECT 14.330 110.200 14.650 110.260 ;
        RECT 168.890 110.200 169.210 110.260 ;
      LAYER via ;
        RECT 168.920 2691.140 169.180 2691.400 ;
        RECT 287.140 2691.140 287.400 2691.400 ;
        RECT 14.360 110.200 14.620 110.460 ;
        RECT 168.920 110.200 169.180 110.460 ;
      LAYER met2 ;
        RECT 287.130 2694.995 287.410 2695.365 ;
        RECT 287.200 2691.430 287.340 2694.995 ;
        RECT 168.920 2691.110 169.180 2691.430 ;
        RECT 287.140 2691.110 287.400 2691.430 ;
        RECT 168.980 110.490 169.120 2691.110 ;
        RECT 14.360 110.170 14.620 110.490 ;
        RECT 168.920 110.170 169.180 110.490 ;
        RECT 14.420 107.285 14.560 110.170 ;
        RECT 14.350 106.915 14.630 107.285 ;
      LAYER via2 ;
        RECT 287.130 2695.040 287.410 2695.320 ;
        RECT 14.350 106.960 14.630 107.240 ;
      LAYER met3 ;
        RECT 287.105 2695.330 287.435 2695.345 ;
        RECT 300.000 2695.330 304.000 2695.440 ;
        RECT 287.105 2695.030 304.000 2695.330 ;
        RECT 287.105 2695.015 287.435 2695.030 ;
        RECT 300.000 2694.840 304.000 2695.030 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 14.325 107.250 14.655 107.265 ;
        RECT -4.800 106.950 14.655 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 14.325 106.935 14.655 106.950 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 331.270 850.240 331.590 850.300 ;
        RECT 379.110 850.240 379.430 850.300 ;
        RECT 331.270 850.100 379.430 850.240 ;
        RECT 331.270 850.040 331.590 850.100 ;
        RECT 379.110 850.040 379.430 850.100 ;
        RECT 737.910 849.900 738.230 849.960 ;
        RECT 772.410 849.900 772.730 849.960 ;
        RECT 737.910 849.760 772.730 849.900 ;
        RECT 737.910 849.700 738.230 849.760 ;
        RECT 772.410 849.700 772.730 849.760 ;
        RECT 579.670 849.220 579.990 849.280 ;
        RECT 593.930 849.220 594.250 849.280 ;
        RECT 579.670 849.080 594.250 849.220 ;
        RECT 579.670 849.020 579.990 849.080 ;
        RECT 593.930 849.020 594.250 849.080 ;
      LAYER via ;
        RECT 331.300 850.040 331.560 850.300 ;
        RECT 379.140 850.040 379.400 850.300 ;
        RECT 737.940 849.700 738.200 849.960 ;
        RECT 772.440 849.700 772.700 849.960 ;
        RECT 579.700 849.020 579.960 849.280 ;
        RECT 593.960 849.020 594.220 849.280 ;
      LAYER met2 ;
        RECT 555.310 852.195 555.590 852.565 ;
        RECT 331.300 850.010 331.560 850.330 ;
        RECT 379.130 850.155 379.410 850.525 ;
        RECT 447.670 850.155 447.950 850.525 ;
        RECT 379.140 850.010 379.400 850.155 ;
        RECT 331.360 849.845 331.500 850.010 ;
        RECT 331.290 849.475 331.570 849.845 ;
        RECT 447.740 849.165 447.880 850.155 ;
        RECT 555.380 849.165 555.520 852.195 ;
        RECT 675.830 851.515 676.110 851.885 ;
        RECT 593.950 850.155 594.230 850.525 ;
        RECT 594.020 849.310 594.160 850.155 ;
        RECT 675.900 849.845 676.040 851.515 ;
        RECT 700.210 850.835 700.490 851.205 ;
        RECT 675.830 849.475 676.110 849.845 ;
        RECT 579.700 849.165 579.960 849.310 ;
        RECT 447.670 848.795 447.950 849.165 ;
        RECT 555.310 848.795 555.590 849.165 ;
        RECT 579.690 848.795 579.970 849.165 ;
        RECT 593.960 848.990 594.220 849.310 ;
        RECT 700.280 849.165 700.420 850.835 ;
        RECT 772.430 850.155 772.710 850.525 ;
        RECT 772.500 849.990 772.640 850.155 ;
        RECT 737.940 849.845 738.200 849.990 ;
        RECT 737.930 849.475 738.210 849.845 ;
        RECT 772.440 849.670 772.700 849.990 ;
        RECT 700.210 848.795 700.490 849.165 ;
      LAYER via2 ;
        RECT 555.310 852.240 555.590 852.520 ;
        RECT 379.130 850.200 379.410 850.480 ;
        RECT 447.670 850.200 447.950 850.480 ;
        RECT 331.290 849.520 331.570 849.800 ;
        RECT 675.830 851.560 676.110 851.840 ;
        RECT 593.950 850.200 594.230 850.480 ;
        RECT 700.210 850.880 700.490 851.160 ;
        RECT 675.830 849.520 676.110 849.800 ;
        RECT 447.670 848.840 447.950 849.120 ;
        RECT 555.310 848.840 555.590 849.120 ;
        RECT 579.690 848.840 579.970 849.120 ;
        RECT 772.430 850.200 772.710 850.480 ;
        RECT 737.930 849.520 738.210 849.800 ;
        RECT 700.210 848.840 700.490 849.120 ;
      LAYER met3 ;
        RECT 288.230 1711.370 288.610 1711.380 ;
        RECT 300.000 1711.370 304.000 1711.480 ;
        RECT 288.230 1711.070 304.000 1711.370 ;
        RECT 288.230 1711.060 288.610 1711.070 ;
        RECT 300.000 1710.880 304.000 1711.070 ;
        RECT 531.110 852.530 531.490 852.540 ;
        RECT 555.285 852.530 555.615 852.545 ;
        RECT 531.110 852.230 555.615 852.530 ;
        RECT 531.110 852.220 531.490 852.230 ;
        RECT 555.285 852.215 555.615 852.230 ;
        RECT 627.710 851.850 628.090 851.860 ;
        RECT 675.805 851.850 676.135 851.865 ;
        RECT 627.710 851.550 676.135 851.850 ;
        RECT 627.710 851.540 628.090 851.550 ;
        RECT 675.805 851.535 676.135 851.550 ;
        RECT 531.110 851.170 531.490 851.180 ;
        RECT 700.185 851.170 700.515 851.185 ;
        RECT 497.110 850.870 531.490 851.170 ;
        RECT 288.230 850.490 288.610 850.500 ;
        RECT 379.105 850.490 379.435 850.505 ;
        RECT 447.645 850.490 447.975 850.505 ;
        RECT 288.230 850.190 304.210 850.490 ;
        RECT 288.230 850.180 288.610 850.190 ;
        RECT 303.910 849.810 304.210 850.190 ;
        RECT 379.105 850.190 410.930 850.490 ;
        RECT 379.105 850.175 379.435 850.190 ;
        RECT 331.265 849.810 331.595 849.825 ;
        RECT 303.910 849.510 331.595 849.810 ;
        RECT 331.265 849.495 331.595 849.510 ;
        RECT 410.630 849.130 410.930 850.190 ;
        RECT 447.645 850.190 482.690 850.490 ;
        RECT 447.645 850.175 447.975 850.190 ;
        RECT 482.390 849.810 482.690 850.190 ;
        RECT 497.110 849.810 497.410 850.870 ;
        RECT 531.110 850.860 531.490 850.870 ;
        RECT 676.510 850.870 700.515 851.170 ;
        RECT 593.925 850.490 594.255 850.505 ;
        RECT 627.710 850.490 628.090 850.500 ;
        RECT 593.925 850.190 628.090 850.490 ;
        RECT 593.925 850.175 594.255 850.190 ;
        RECT 627.710 850.180 628.090 850.190 ;
        RECT 482.390 849.510 497.410 849.810 ;
        RECT 675.805 849.810 676.135 849.825 ;
        RECT 676.510 849.810 676.810 850.870 ;
        RECT 700.185 850.855 700.515 850.870 ;
        RECT 772.405 850.490 772.735 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 772.405 850.190 807.450 850.490 ;
        RECT 772.405 850.175 772.735 850.190 ;
        RECT 737.905 849.810 738.235 849.825 ;
        RECT 675.805 849.510 676.810 849.810 ;
        RECT 724.350 849.510 738.235 849.810 ;
        RECT 807.150 849.810 807.450 850.190 ;
        RECT 855.910 850.190 904.050 850.490 ;
        RECT 807.150 849.510 855.290 849.810 ;
        RECT 675.805 849.495 676.135 849.510 ;
        RECT 447.645 849.130 447.975 849.145 ;
        RECT 410.630 848.830 447.975 849.130 ;
        RECT 447.645 848.815 447.975 848.830 ;
        RECT 555.285 849.130 555.615 849.145 ;
        RECT 579.665 849.130 579.995 849.145 ;
        RECT 555.285 848.830 579.995 849.130 ;
        RECT 555.285 848.815 555.615 848.830 ;
        RECT 579.665 848.815 579.995 848.830 ;
        RECT 700.185 849.130 700.515 849.145 ;
        RECT 724.350 849.130 724.650 849.510 ;
        RECT 737.905 849.495 738.235 849.510 ;
        RECT 700.185 848.830 724.650 849.130 ;
        RECT 854.990 849.130 855.290 849.510 ;
        RECT 855.910 849.130 856.210 850.190 ;
        RECT 903.750 849.810 904.050 850.190 ;
        RECT 952.510 850.190 1000.650 850.490 ;
        RECT 903.750 849.510 951.890 849.810 ;
        RECT 854.990 848.830 856.210 849.130 ;
        RECT 951.590 849.130 951.890 849.510 ;
        RECT 952.510 849.130 952.810 850.190 ;
        RECT 1000.350 849.810 1000.650 850.190 ;
        RECT 1049.110 850.190 1097.250 850.490 ;
        RECT 1000.350 849.510 1048.490 849.810 ;
        RECT 951.590 848.830 952.810 849.130 ;
        RECT 1048.190 849.130 1048.490 849.510 ;
        RECT 1049.110 849.130 1049.410 850.190 ;
        RECT 1096.950 849.810 1097.250 850.190 ;
        RECT 1145.710 850.190 1193.850 850.490 ;
        RECT 1096.950 849.510 1145.090 849.810 ;
        RECT 1048.190 848.830 1049.410 849.130 ;
        RECT 1144.790 849.130 1145.090 849.510 ;
        RECT 1145.710 849.130 1146.010 850.190 ;
        RECT 1193.550 849.810 1193.850 850.190 ;
        RECT 1242.310 850.190 1290.450 850.490 ;
        RECT 1193.550 849.510 1241.690 849.810 ;
        RECT 1144.790 848.830 1146.010 849.130 ;
        RECT 1241.390 849.130 1241.690 849.510 ;
        RECT 1242.310 849.130 1242.610 850.190 ;
        RECT 1290.150 849.810 1290.450 850.190 ;
        RECT 1338.910 850.190 1387.050 850.490 ;
        RECT 1290.150 849.510 1338.290 849.810 ;
        RECT 1241.390 848.830 1242.610 849.130 ;
        RECT 1337.990 849.130 1338.290 849.510 ;
        RECT 1338.910 849.130 1339.210 850.190 ;
        RECT 1386.750 849.810 1387.050 850.190 ;
        RECT 1435.510 850.190 1483.650 850.490 ;
        RECT 1386.750 849.510 1434.890 849.810 ;
        RECT 1337.990 848.830 1339.210 849.130 ;
        RECT 1434.590 849.130 1434.890 849.510 ;
        RECT 1435.510 849.130 1435.810 850.190 ;
        RECT 1483.350 849.810 1483.650 850.190 ;
        RECT 1532.110 850.190 1580.250 850.490 ;
        RECT 1483.350 849.510 1531.490 849.810 ;
        RECT 1434.590 848.830 1435.810 849.130 ;
        RECT 1531.190 849.130 1531.490 849.510 ;
        RECT 1532.110 849.130 1532.410 850.190 ;
        RECT 1579.950 849.810 1580.250 850.190 ;
        RECT 1628.710 850.190 1676.850 850.490 ;
        RECT 1579.950 849.510 1628.090 849.810 ;
        RECT 1531.190 848.830 1532.410 849.130 ;
        RECT 1627.790 849.130 1628.090 849.510 ;
        RECT 1628.710 849.130 1629.010 850.190 ;
        RECT 1676.550 849.810 1676.850 850.190 ;
        RECT 1725.310 850.190 1773.450 850.490 ;
        RECT 1676.550 849.510 1724.690 849.810 ;
        RECT 1627.790 848.830 1629.010 849.130 ;
        RECT 1724.390 849.130 1724.690 849.510 ;
        RECT 1725.310 849.130 1725.610 850.190 ;
        RECT 1773.150 849.810 1773.450 850.190 ;
        RECT 1821.910 850.190 1870.050 850.490 ;
        RECT 1773.150 849.510 1821.290 849.810 ;
        RECT 1724.390 848.830 1725.610 849.130 ;
        RECT 1820.990 849.130 1821.290 849.510 ;
        RECT 1821.910 849.130 1822.210 850.190 ;
        RECT 1869.750 849.810 1870.050 850.190 ;
        RECT 1918.510 850.190 1966.650 850.490 ;
        RECT 1869.750 849.510 1917.890 849.810 ;
        RECT 1820.990 848.830 1822.210 849.130 ;
        RECT 1917.590 849.130 1917.890 849.510 ;
        RECT 1918.510 849.130 1918.810 850.190 ;
        RECT 1966.350 849.810 1966.650 850.190 ;
        RECT 2015.110 850.190 2063.250 850.490 ;
        RECT 1966.350 849.510 2014.490 849.810 ;
        RECT 1917.590 848.830 1918.810 849.130 ;
        RECT 2014.190 849.130 2014.490 849.510 ;
        RECT 2015.110 849.130 2015.410 850.190 ;
        RECT 2062.950 849.810 2063.250 850.190 ;
        RECT 2111.710 850.190 2159.850 850.490 ;
        RECT 2062.950 849.510 2111.090 849.810 ;
        RECT 2014.190 848.830 2015.410 849.130 ;
        RECT 2110.790 849.130 2111.090 849.510 ;
        RECT 2111.710 849.130 2112.010 850.190 ;
        RECT 2159.550 849.810 2159.850 850.190 ;
        RECT 2208.310 850.190 2256.450 850.490 ;
        RECT 2159.550 849.510 2207.690 849.810 ;
        RECT 2110.790 848.830 2112.010 849.130 ;
        RECT 2207.390 849.130 2207.690 849.510 ;
        RECT 2208.310 849.130 2208.610 850.190 ;
        RECT 2256.150 849.810 2256.450 850.190 ;
        RECT 2304.910 850.190 2353.050 850.490 ;
        RECT 2256.150 849.510 2304.290 849.810 ;
        RECT 2207.390 848.830 2208.610 849.130 ;
        RECT 2303.990 849.130 2304.290 849.510 ;
        RECT 2304.910 849.130 2305.210 850.190 ;
        RECT 2352.750 849.810 2353.050 850.190 ;
        RECT 2401.510 850.190 2449.650 850.490 ;
        RECT 2352.750 849.510 2400.890 849.810 ;
        RECT 2303.990 848.830 2305.210 849.130 ;
        RECT 2400.590 849.130 2400.890 849.510 ;
        RECT 2401.510 849.130 2401.810 850.190 ;
        RECT 2449.350 849.810 2449.650 850.190 ;
        RECT 2498.110 850.190 2546.250 850.490 ;
        RECT 2449.350 849.510 2497.490 849.810 ;
        RECT 2400.590 848.830 2401.810 849.130 ;
        RECT 2497.190 849.130 2497.490 849.510 ;
        RECT 2498.110 849.130 2498.410 850.190 ;
        RECT 2545.950 849.810 2546.250 850.190 ;
        RECT 2594.710 850.190 2642.850 850.490 ;
        RECT 2545.950 849.510 2594.090 849.810 ;
        RECT 2497.190 848.830 2498.410 849.130 ;
        RECT 2593.790 849.130 2594.090 849.510 ;
        RECT 2594.710 849.130 2595.010 850.190 ;
        RECT 2642.550 849.810 2642.850 850.190 ;
        RECT 2691.310 850.190 2739.450 850.490 ;
        RECT 2642.550 849.510 2690.690 849.810 ;
        RECT 2593.790 848.830 2595.010 849.130 ;
        RECT 2690.390 849.130 2690.690 849.510 ;
        RECT 2691.310 849.130 2691.610 850.190 ;
        RECT 2739.150 849.810 2739.450 850.190 ;
        RECT 2787.910 850.190 2836.050 850.490 ;
        RECT 2739.150 849.510 2787.290 849.810 ;
        RECT 2690.390 848.830 2691.610 849.130 ;
        RECT 2786.990 849.130 2787.290 849.510 ;
        RECT 2787.910 849.130 2788.210 850.190 ;
        RECT 2835.750 849.810 2836.050 850.190 ;
        RECT 2916.710 850.190 2924.800 850.490 ;
        RECT 2916.710 849.810 2917.010 850.190 ;
        RECT 2835.750 849.510 2883.890 849.810 ;
        RECT 2786.990 848.830 2788.210 849.130 ;
        RECT 2883.590 849.130 2883.890 849.510 ;
        RECT 2884.510 849.510 2917.010 849.810 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
        RECT 2884.510 849.130 2884.810 849.510 ;
        RECT 2883.590 848.830 2884.810 849.130 ;
        RECT 700.185 848.815 700.515 848.830 ;
      LAYER via3 ;
        RECT 288.260 1711.060 288.580 1711.380 ;
        RECT 531.140 852.220 531.460 852.540 ;
        RECT 627.740 851.540 628.060 851.860 ;
        RECT 288.260 850.180 288.580 850.500 ;
        RECT 531.140 850.860 531.460 851.180 ;
        RECT 627.740 850.180 628.060 850.500 ;
      LAYER met4 ;
        RECT 288.255 1711.055 288.585 1711.385 ;
        RECT 288.270 850.505 288.570 1711.055 ;
        RECT 531.135 852.215 531.465 852.545 ;
        RECT 531.150 851.185 531.450 852.215 ;
        RECT 627.735 851.535 628.065 851.865 ;
        RECT 531.135 850.855 531.465 851.185 ;
        RECT 627.750 850.505 628.050 851.535 ;
        RECT 288.255 850.175 288.585 850.505 ;
        RECT 627.735 850.175 628.065 850.505 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 346.910 1084.840 347.230 1084.900 ;
        RECT 386.010 1084.840 386.330 1084.900 ;
        RECT 346.910 1084.700 386.330 1084.840 ;
        RECT 346.910 1084.640 347.230 1084.700 ;
        RECT 386.010 1084.640 386.330 1084.700 ;
        RECT 447.650 1084.500 447.970 1084.560 ;
        RECT 458.690 1084.500 459.010 1084.560 ;
        RECT 447.650 1084.360 459.010 1084.500 ;
        RECT 447.650 1084.300 447.970 1084.360 ;
        RECT 458.690 1084.300 459.010 1084.360 ;
        RECT 737.910 1084.500 738.230 1084.560 ;
        RECT 772.410 1084.500 772.730 1084.560 ;
        RECT 737.910 1084.360 772.730 1084.500 ;
        RECT 737.910 1084.300 738.230 1084.360 ;
        RECT 772.410 1084.300 772.730 1084.360 ;
        RECT 579.670 1083.820 579.990 1083.880 ;
        RECT 593.930 1083.820 594.250 1083.880 ;
        RECT 579.670 1083.680 594.250 1083.820 ;
        RECT 579.670 1083.620 579.990 1083.680 ;
        RECT 593.930 1083.620 594.250 1083.680 ;
      LAYER via ;
        RECT 346.940 1084.640 347.200 1084.900 ;
        RECT 386.040 1084.640 386.300 1084.900 ;
        RECT 447.680 1084.300 447.940 1084.560 ;
        RECT 458.720 1084.300 458.980 1084.560 ;
        RECT 737.940 1084.300 738.200 1084.560 ;
        RECT 772.440 1084.300 772.700 1084.560 ;
        RECT 579.700 1083.620 579.960 1083.880 ;
        RECT 593.960 1083.620 594.220 1083.880 ;
      LAYER met2 ;
        RECT 675.830 1086.115 676.110 1086.485 ;
        RECT 346.940 1084.610 347.200 1084.930 ;
        RECT 386.030 1084.755 386.310 1085.125 ;
        RECT 593.950 1084.755 594.230 1085.125 ;
        RECT 386.040 1084.610 386.300 1084.755 ;
        RECT 347.000 1084.445 347.140 1084.610 ;
        RECT 447.680 1084.445 447.940 1084.590 ;
        RECT 458.720 1084.445 458.980 1084.590 ;
        RECT 346.930 1084.075 347.210 1084.445 ;
        RECT 447.670 1084.075 447.950 1084.445 ;
        RECT 458.710 1084.075 458.990 1084.445 ;
        RECT 594.020 1083.910 594.160 1084.755 ;
        RECT 675.900 1084.445 676.040 1086.115 ;
        RECT 700.210 1085.435 700.490 1085.805 ;
        RECT 675.830 1084.075 676.110 1084.445 ;
        RECT 579.700 1083.765 579.960 1083.910 ;
        RECT 579.690 1083.395 579.970 1083.765 ;
        RECT 593.960 1083.590 594.220 1083.910 ;
        RECT 700.280 1083.765 700.420 1085.435 ;
        RECT 772.430 1084.755 772.710 1085.125 ;
        RECT 772.500 1084.590 772.640 1084.755 ;
        RECT 737.940 1084.445 738.200 1084.590 ;
        RECT 737.930 1084.075 738.210 1084.445 ;
        RECT 772.440 1084.270 772.700 1084.590 ;
        RECT 700.210 1083.395 700.490 1083.765 ;
      LAYER via2 ;
        RECT 675.830 1086.160 676.110 1086.440 ;
        RECT 386.030 1084.800 386.310 1085.080 ;
        RECT 593.950 1084.800 594.230 1085.080 ;
        RECT 346.930 1084.120 347.210 1084.400 ;
        RECT 447.670 1084.120 447.950 1084.400 ;
        RECT 458.710 1084.120 458.990 1084.400 ;
        RECT 700.210 1085.480 700.490 1085.760 ;
        RECT 675.830 1084.120 676.110 1084.400 ;
        RECT 579.690 1083.440 579.970 1083.720 ;
        RECT 772.430 1084.800 772.710 1085.080 ;
        RECT 737.930 1084.120 738.210 1084.400 ;
        RECT 700.210 1083.440 700.490 1083.720 ;
      LAYER met3 ;
        RECT 286.390 1739.930 286.770 1739.940 ;
        RECT 300.000 1739.930 304.000 1740.040 ;
        RECT 286.390 1739.630 304.000 1739.930 ;
        RECT 286.390 1739.620 286.770 1739.630 ;
        RECT 300.000 1739.440 304.000 1739.630 ;
        RECT 627.710 1086.450 628.090 1086.460 ;
        RECT 675.805 1086.450 676.135 1086.465 ;
        RECT 627.710 1086.150 676.135 1086.450 ;
        RECT 627.710 1086.140 628.090 1086.150 ;
        RECT 675.805 1086.135 676.135 1086.150 ;
        RECT 700.185 1085.770 700.515 1085.785 ;
        RECT 676.510 1085.470 700.515 1085.770 ;
        RECT 286.390 1085.090 286.770 1085.100 ;
        RECT 386.005 1085.090 386.335 1085.105 ;
        RECT 593.925 1085.090 594.255 1085.105 ;
        RECT 627.710 1085.090 628.090 1085.100 ;
        RECT 286.390 1084.790 304.210 1085.090 ;
        RECT 286.390 1084.780 286.770 1084.790 ;
        RECT 303.910 1084.410 304.210 1084.790 ;
        RECT 386.005 1084.790 400.810 1085.090 ;
        RECT 386.005 1084.775 386.335 1084.790 ;
        RECT 346.905 1084.410 347.235 1084.425 ;
        RECT 303.910 1084.110 347.235 1084.410 ;
        RECT 400.510 1084.410 400.810 1084.790 ;
        RECT 482.390 1084.790 545.250 1085.090 ;
        RECT 447.645 1084.410 447.975 1084.425 ;
        RECT 400.510 1084.110 447.975 1084.410 ;
        RECT 346.905 1084.095 347.235 1084.110 ;
        RECT 447.645 1084.095 447.975 1084.110 ;
        RECT 458.685 1084.410 459.015 1084.425 ;
        RECT 482.390 1084.410 482.690 1084.790 ;
        RECT 458.685 1084.110 482.690 1084.410 ;
        RECT 458.685 1084.095 459.015 1084.110 ;
        RECT 544.950 1083.730 545.250 1084.790 ;
        RECT 593.925 1084.790 628.090 1085.090 ;
        RECT 593.925 1084.775 594.255 1084.790 ;
        RECT 627.710 1084.780 628.090 1084.790 ;
        RECT 675.805 1084.410 676.135 1084.425 ;
        RECT 676.510 1084.410 676.810 1085.470 ;
        RECT 700.185 1085.455 700.515 1085.470 ;
        RECT 772.405 1085.090 772.735 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 772.405 1084.790 807.450 1085.090 ;
        RECT 772.405 1084.775 772.735 1084.790 ;
        RECT 737.905 1084.410 738.235 1084.425 ;
        RECT 675.805 1084.110 676.810 1084.410 ;
        RECT 724.350 1084.110 738.235 1084.410 ;
        RECT 807.150 1084.410 807.450 1084.790 ;
        RECT 855.910 1084.790 904.050 1085.090 ;
        RECT 807.150 1084.110 855.290 1084.410 ;
        RECT 675.805 1084.095 676.135 1084.110 ;
        RECT 579.665 1083.730 579.995 1083.745 ;
        RECT 544.950 1083.430 579.995 1083.730 ;
        RECT 579.665 1083.415 579.995 1083.430 ;
        RECT 700.185 1083.730 700.515 1083.745 ;
        RECT 724.350 1083.730 724.650 1084.110 ;
        RECT 737.905 1084.095 738.235 1084.110 ;
        RECT 700.185 1083.430 724.650 1083.730 ;
        RECT 854.990 1083.730 855.290 1084.110 ;
        RECT 855.910 1083.730 856.210 1084.790 ;
        RECT 903.750 1084.410 904.050 1084.790 ;
        RECT 952.510 1084.790 1000.650 1085.090 ;
        RECT 903.750 1084.110 951.890 1084.410 ;
        RECT 854.990 1083.430 856.210 1083.730 ;
        RECT 951.590 1083.730 951.890 1084.110 ;
        RECT 952.510 1083.730 952.810 1084.790 ;
        RECT 1000.350 1084.410 1000.650 1084.790 ;
        RECT 1049.110 1084.790 1097.250 1085.090 ;
        RECT 1000.350 1084.110 1048.490 1084.410 ;
        RECT 951.590 1083.430 952.810 1083.730 ;
        RECT 1048.190 1083.730 1048.490 1084.110 ;
        RECT 1049.110 1083.730 1049.410 1084.790 ;
        RECT 1096.950 1084.410 1097.250 1084.790 ;
        RECT 1145.710 1084.790 1193.850 1085.090 ;
        RECT 1096.950 1084.110 1145.090 1084.410 ;
        RECT 1048.190 1083.430 1049.410 1083.730 ;
        RECT 1144.790 1083.730 1145.090 1084.110 ;
        RECT 1145.710 1083.730 1146.010 1084.790 ;
        RECT 1193.550 1084.410 1193.850 1084.790 ;
        RECT 1242.310 1084.790 1290.450 1085.090 ;
        RECT 1193.550 1084.110 1241.690 1084.410 ;
        RECT 1144.790 1083.430 1146.010 1083.730 ;
        RECT 1241.390 1083.730 1241.690 1084.110 ;
        RECT 1242.310 1083.730 1242.610 1084.790 ;
        RECT 1290.150 1084.410 1290.450 1084.790 ;
        RECT 1338.910 1084.790 1387.050 1085.090 ;
        RECT 1290.150 1084.110 1338.290 1084.410 ;
        RECT 1241.390 1083.430 1242.610 1083.730 ;
        RECT 1337.990 1083.730 1338.290 1084.110 ;
        RECT 1338.910 1083.730 1339.210 1084.790 ;
        RECT 1386.750 1084.410 1387.050 1084.790 ;
        RECT 1435.510 1084.790 1483.650 1085.090 ;
        RECT 1386.750 1084.110 1434.890 1084.410 ;
        RECT 1337.990 1083.430 1339.210 1083.730 ;
        RECT 1434.590 1083.730 1434.890 1084.110 ;
        RECT 1435.510 1083.730 1435.810 1084.790 ;
        RECT 1483.350 1084.410 1483.650 1084.790 ;
        RECT 1532.110 1084.790 1580.250 1085.090 ;
        RECT 1483.350 1084.110 1531.490 1084.410 ;
        RECT 1434.590 1083.430 1435.810 1083.730 ;
        RECT 1531.190 1083.730 1531.490 1084.110 ;
        RECT 1532.110 1083.730 1532.410 1084.790 ;
        RECT 1579.950 1084.410 1580.250 1084.790 ;
        RECT 1628.710 1084.790 1676.850 1085.090 ;
        RECT 1579.950 1084.110 1628.090 1084.410 ;
        RECT 1531.190 1083.430 1532.410 1083.730 ;
        RECT 1627.790 1083.730 1628.090 1084.110 ;
        RECT 1628.710 1083.730 1629.010 1084.790 ;
        RECT 1676.550 1084.410 1676.850 1084.790 ;
        RECT 1725.310 1084.790 1773.450 1085.090 ;
        RECT 1676.550 1084.110 1724.690 1084.410 ;
        RECT 1627.790 1083.430 1629.010 1083.730 ;
        RECT 1724.390 1083.730 1724.690 1084.110 ;
        RECT 1725.310 1083.730 1725.610 1084.790 ;
        RECT 1773.150 1084.410 1773.450 1084.790 ;
        RECT 1821.910 1084.790 1870.050 1085.090 ;
        RECT 1773.150 1084.110 1821.290 1084.410 ;
        RECT 1724.390 1083.430 1725.610 1083.730 ;
        RECT 1820.990 1083.730 1821.290 1084.110 ;
        RECT 1821.910 1083.730 1822.210 1084.790 ;
        RECT 1869.750 1084.410 1870.050 1084.790 ;
        RECT 1918.510 1084.790 1966.650 1085.090 ;
        RECT 1869.750 1084.110 1917.890 1084.410 ;
        RECT 1820.990 1083.430 1822.210 1083.730 ;
        RECT 1917.590 1083.730 1917.890 1084.110 ;
        RECT 1918.510 1083.730 1918.810 1084.790 ;
        RECT 1966.350 1084.410 1966.650 1084.790 ;
        RECT 2015.110 1084.790 2063.250 1085.090 ;
        RECT 1966.350 1084.110 2014.490 1084.410 ;
        RECT 1917.590 1083.430 1918.810 1083.730 ;
        RECT 2014.190 1083.730 2014.490 1084.110 ;
        RECT 2015.110 1083.730 2015.410 1084.790 ;
        RECT 2062.950 1084.410 2063.250 1084.790 ;
        RECT 2111.710 1084.790 2159.850 1085.090 ;
        RECT 2062.950 1084.110 2111.090 1084.410 ;
        RECT 2014.190 1083.430 2015.410 1083.730 ;
        RECT 2110.790 1083.730 2111.090 1084.110 ;
        RECT 2111.710 1083.730 2112.010 1084.790 ;
        RECT 2159.550 1084.410 2159.850 1084.790 ;
        RECT 2208.310 1084.790 2256.450 1085.090 ;
        RECT 2159.550 1084.110 2207.690 1084.410 ;
        RECT 2110.790 1083.430 2112.010 1083.730 ;
        RECT 2207.390 1083.730 2207.690 1084.110 ;
        RECT 2208.310 1083.730 2208.610 1084.790 ;
        RECT 2256.150 1084.410 2256.450 1084.790 ;
        RECT 2304.910 1084.790 2353.050 1085.090 ;
        RECT 2256.150 1084.110 2304.290 1084.410 ;
        RECT 2207.390 1083.430 2208.610 1083.730 ;
        RECT 2303.990 1083.730 2304.290 1084.110 ;
        RECT 2304.910 1083.730 2305.210 1084.790 ;
        RECT 2352.750 1084.410 2353.050 1084.790 ;
        RECT 2401.510 1084.790 2449.650 1085.090 ;
        RECT 2352.750 1084.110 2400.890 1084.410 ;
        RECT 2303.990 1083.430 2305.210 1083.730 ;
        RECT 2400.590 1083.730 2400.890 1084.110 ;
        RECT 2401.510 1083.730 2401.810 1084.790 ;
        RECT 2449.350 1084.410 2449.650 1084.790 ;
        RECT 2498.110 1084.790 2546.250 1085.090 ;
        RECT 2449.350 1084.110 2497.490 1084.410 ;
        RECT 2400.590 1083.430 2401.810 1083.730 ;
        RECT 2497.190 1083.730 2497.490 1084.110 ;
        RECT 2498.110 1083.730 2498.410 1084.790 ;
        RECT 2545.950 1084.410 2546.250 1084.790 ;
        RECT 2594.710 1084.790 2642.850 1085.090 ;
        RECT 2545.950 1084.110 2594.090 1084.410 ;
        RECT 2497.190 1083.430 2498.410 1083.730 ;
        RECT 2593.790 1083.730 2594.090 1084.110 ;
        RECT 2594.710 1083.730 2595.010 1084.790 ;
        RECT 2642.550 1084.410 2642.850 1084.790 ;
        RECT 2691.310 1084.790 2739.450 1085.090 ;
        RECT 2642.550 1084.110 2690.690 1084.410 ;
        RECT 2593.790 1083.430 2595.010 1083.730 ;
        RECT 2690.390 1083.730 2690.690 1084.110 ;
        RECT 2691.310 1083.730 2691.610 1084.790 ;
        RECT 2739.150 1084.410 2739.450 1084.790 ;
        RECT 2787.910 1084.790 2836.050 1085.090 ;
        RECT 2739.150 1084.110 2787.290 1084.410 ;
        RECT 2690.390 1083.430 2691.610 1083.730 ;
        RECT 2786.990 1083.730 2787.290 1084.110 ;
        RECT 2787.910 1083.730 2788.210 1084.790 ;
        RECT 2835.750 1084.410 2836.050 1084.790 ;
        RECT 2916.710 1084.790 2924.800 1085.090 ;
        RECT 2916.710 1084.410 2917.010 1084.790 ;
        RECT 2835.750 1084.110 2883.890 1084.410 ;
        RECT 2786.990 1083.430 2788.210 1083.730 ;
        RECT 2883.590 1083.730 2883.890 1084.110 ;
        RECT 2884.510 1084.110 2917.010 1084.410 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
        RECT 2884.510 1083.730 2884.810 1084.110 ;
        RECT 2883.590 1083.430 2884.810 1083.730 ;
        RECT 700.185 1083.415 700.515 1083.430 ;
      LAYER via3 ;
        RECT 286.420 1739.620 286.740 1739.940 ;
        RECT 627.740 1086.140 628.060 1086.460 ;
        RECT 286.420 1084.780 286.740 1085.100 ;
        RECT 627.740 1084.780 628.060 1085.100 ;
      LAYER met4 ;
        RECT 286.415 1739.615 286.745 1739.945 ;
        RECT 286.430 1085.105 286.730 1739.615 ;
        RECT 627.735 1086.135 628.065 1086.465 ;
        RECT 627.750 1085.105 628.050 1086.135 ;
        RECT 286.415 1084.775 286.745 1085.105 ;
        RECT 627.735 1084.775 628.065 1085.105 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 737.910 1319.100 738.230 1319.160 ;
        RECT 772.410 1319.100 772.730 1319.160 ;
        RECT 737.910 1318.960 772.730 1319.100 ;
        RECT 737.910 1318.900 738.230 1318.960 ;
        RECT 772.410 1318.900 772.730 1318.960 ;
        RECT 579.670 1318.420 579.990 1318.480 ;
        RECT 593.930 1318.420 594.250 1318.480 ;
        RECT 579.670 1318.280 594.250 1318.420 ;
        RECT 579.670 1318.220 579.990 1318.280 ;
        RECT 593.930 1318.220 594.250 1318.280 ;
      LAYER via ;
        RECT 737.940 1318.900 738.200 1319.160 ;
        RECT 772.440 1318.900 772.700 1319.160 ;
        RECT 579.700 1318.220 579.960 1318.480 ;
        RECT 593.960 1318.220 594.220 1318.480 ;
      LAYER met2 ;
        RECT 555.310 1321.395 555.590 1321.765 ;
        RECT 555.380 1318.365 555.520 1321.395 ;
        RECT 675.830 1320.715 676.110 1321.085 ;
        RECT 593.950 1319.355 594.230 1319.725 ;
        RECT 594.020 1318.510 594.160 1319.355 ;
        RECT 675.900 1319.045 676.040 1320.715 ;
        RECT 700.210 1320.035 700.490 1320.405 ;
        RECT 675.830 1318.675 676.110 1319.045 ;
        RECT 579.700 1318.365 579.960 1318.510 ;
        RECT 555.310 1317.995 555.590 1318.365 ;
        RECT 579.690 1317.995 579.970 1318.365 ;
        RECT 593.960 1318.190 594.220 1318.510 ;
        RECT 700.280 1318.365 700.420 1320.035 ;
        RECT 772.430 1319.355 772.710 1319.725 ;
        RECT 772.500 1319.190 772.640 1319.355 ;
        RECT 737.940 1319.045 738.200 1319.190 ;
        RECT 737.930 1318.675 738.210 1319.045 ;
        RECT 772.440 1318.870 772.700 1319.190 ;
        RECT 700.210 1317.995 700.490 1318.365 ;
      LAYER via2 ;
        RECT 555.310 1321.440 555.590 1321.720 ;
        RECT 675.830 1320.760 676.110 1321.040 ;
        RECT 593.950 1319.400 594.230 1319.680 ;
        RECT 700.210 1320.080 700.490 1320.360 ;
        RECT 675.830 1318.720 676.110 1319.000 ;
        RECT 555.310 1318.040 555.590 1318.320 ;
        RECT 579.690 1318.040 579.970 1318.320 ;
        RECT 772.430 1319.400 772.710 1319.680 ;
        RECT 737.930 1318.720 738.210 1319.000 ;
        RECT 700.210 1318.040 700.490 1318.320 ;
      LAYER met3 ;
        RECT 284.550 1769.170 284.930 1769.180 ;
        RECT 300.000 1769.170 304.000 1769.280 ;
        RECT 284.550 1768.870 304.000 1769.170 ;
        RECT 284.550 1768.860 284.930 1768.870 ;
        RECT 300.000 1768.680 304.000 1768.870 ;
        RECT 531.110 1321.730 531.490 1321.740 ;
        RECT 555.285 1321.730 555.615 1321.745 ;
        RECT 531.110 1321.430 555.615 1321.730 ;
        RECT 531.110 1321.420 531.490 1321.430 ;
        RECT 555.285 1321.415 555.615 1321.430 ;
        RECT 627.710 1321.050 628.090 1321.060 ;
        RECT 675.805 1321.050 676.135 1321.065 ;
        RECT 627.710 1320.750 676.135 1321.050 ;
        RECT 627.710 1320.740 628.090 1320.750 ;
        RECT 675.805 1320.735 676.135 1320.750 ;
        RECT 434.510 1320.370 434.890 1320.380 ;
        RECT 482.350 1320.370 482.730 1320.380 ;
        RECT 531.110 1320.370 531.490 1320.380 ;
        RECT 700.185 1320.370 700.515 1320.385 ;
        RECT 434.510 1320.070 482.730 1320.370 ;
        RECT 434.510 1320.060 434.890 1320.070 ;
        RECT 482.350 1320.060 482.730 1320.070 ;
        RECT 497.110 1320.070 531.490 1320.370 ;
        RECT 284.550 1319.690 284.930 1319.700 ;
        RECT 284.550 1319.390 324.450 1319.690 ;
        RECT 284.550 1319.380 284.930 1319.390 ;
        RECT 324.150 1318.330 324.450 1319.390 ;
        RECT 351.750 1319.390 410.930 1319.690 ;
        RECT 351.750 1318.330 352.050 1319.390 ;
        RECT 324.150 1318.030 352.050 1318.330 ;
        RECT 410.630 1318.330 410.930 1319.390 ;
        RECT 482.350 1319.010 482.730 1319.020 ;
        RECT 497.110 1319.010 497.410 1320.070 ;
        RECT 531.110 1320.060 531.490 1320.070 ;
        RECT 676.510 1320.070 700.515 1320.370 ;
        RECT 593.925 1319.690 594.255 1319.705 ;
        RECT 627.710 1319.690 628.090 1319.700 ;
        RECT 593.925 1319.390 628.090 1319.690 ;
        RECT 593.925 1319.375 594.255 1319.390 ;
        RECT 627.710 1319.380 628.090 1319.390 ;
        RECT 482.350 1318.710 497.410 1319.010 ;
        RECT 675.805 1319.010 676.135 1319.025 ;
        RECT 676.510 1319.010 676.810 1320.070 ;
        RECT 700.185 1320.055 700.515 1320.070 ;
        RECT 772.405 1319.690 772.735 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 772.405 1319.390 807.450 1319.690 ;
        RECT 772.405 1319.375 772.735 1319.390 ;
        RECT 737.905 1319.010 738.235 1319.025 ;
        RECT 675.805 1318.710 676.810 1319.010 ;
        RECT 724.350 1318.710 738.235 1319.010 ;
        RECT 807.150 1319.010 807.450 1319.390 ;
        RECT 855.910 1319.390 904.050 1319.690 ;
        RECT 807.150 1318.710 855.290 1319.010 ;
        RECT 482.350 1318.700 482.730 1318.710 ;
        RECT 675.805 1318.695 676.135 1318.710 ;
        RECT 434.510 1318.330 434.890 1318.340 ;
        RECT 410.630 1318.030 434.890 1318.330 ;
        RECT 434.510 1318.020 434.890 1318.030 ;
        RECT 555.285 1318.330 555.615 1318.345 ;
        RECT 579.665 1318.330 579.995 1318.345 ;
        RECT 555.285 1318.030 579.995 1318.330 ;
        RECT 555.285 1318.015 555.615 1318.030 ;
        RECT 579.665 1318.015 579.995 1318.030 ;
        RECT 700.185 1318.330 700.515 1318.345 ;
        RECT 724.350 1318.330 724.650 1318.710 ;
        RECT 737.905 1318.695 738.235 1318.710 ;
        RECT 700.185 1318.030 724.650 1318.330 ;
        RECT 854.990 1318.330 855.290 1318.710 ;
        RECT 855.910 1318.330 856.210 1319.390 ;
        RECT 903.750 1319.010 904.050 1319.390 ;
        RECT 952.510 1319.390 1000.650 1319.690 ;
        RECT 903.750 1318.710 951.890 1319.010 ;
        RECT 854.990 1318.030 856.210 1318.330 ;
        RECT 951.590 1318.330 951.890 1318.710 ;
        RECT 952.510 1318.330 952.810 1319.390 ;
        RECT 1000.350 1319.010 1000.650 1319.390 ;
        RECT 1049.110 1319.390 1097.250 1319.690 ;
        RECT 1000.350 1318.710 1048.490 1319.010 ;
        RECT 951.590 1318.030 952.810 1318.330 ;
        RECT 1048.190 1318.330 1048.490 1318.710 ;
        RECT 1049.110 1318.330 1049.410 1319.390 ;
        RECT 1096.950 1319.010 1097.250 1319.390 ;
        RECT 1145.710 1319.390 1193.850 1319.690 ;
        RECT 1096.950 1318.710 1145.090 1319.010 ;
        RECT 1048.190 1318.030 1049.410 1318.330 ;
        RECT 1144.790 1318.330 1145.090 1318.710 ;
        RECT 1145.710 1318.330 1146.010 1319.390 ;
        RECT 1193.550 1319.010 1193.850 1319.390 ;
        RECT 1242.310 1319.390 1290.450 1319.690 ;
        RECT 1193.550 1318.710 1241.690 1319.010 ;
        RECT 1144.790 1318.030 1146.010 1318.330 ;
        RECT 1241.390 1318.330 1241.690 1318.710 ;
        RECT 1242.310 1318.330 1242.610 1319.390 ;
        RECT 1290.150 1319.010 1290.450 1319.390 ;
        RECT 1338.910 1319.390 1387.050 1319.690 ;
        RECT 1290.150 1318.710 1338.290 1319.010 ;
        RECT 1241.390 1318.030 1242.610 1318.330 ;
        RECT 1337.990 1318.330 1338.290 1318.710 ;
        RECT 1338.910 1318.330 1339.210 1319.390 ;
        RECT 1386.750 1319.010 1387.050 1319.390 ;
        RECT 1435.510 1319.390 1483.650 1319.690 ;
        RECT 1386.750 1318.710 1434.890 1319.010 ;
        RECT 1337.990 1318.030 1339.210 1318.330 ;
        RECT 1434.590 1318.330 1434.890 1318.710 ;
        RECT 1435.510 1318.330 1435.810 1319.390 ;
        RECT 1483.350 1319.010 1483.650 1319.390 ;
        RECT 1532.110 1319.390 1580.250 1319.690 ;
        RECT 1483.350 1318.710 1531.490 1319.010 ;
        RECT 1434.590 1318.030 1435.810 1318.330 ;
        RECT 1531.190 1318.330 1531.490 1318.710 ;
        RECT 1532.110 1318.330 1532.410 1319.390 ;
        RECT 1579.950 1319.010 1580.250 1319.390 ;
        RECT 1628.710 1319.390 1676.850 1319.690 ;
        RECT 1579.950 1318.710 1628.090 1319.010 ;
        RECT 1531.190 1318.030 1532.410 1318.330 ;
        RECT 1627.790 1318.330 1628.090 1318.710 ;
        RECT 1628.710 1318.330 1629.010 1319.390 ;
        RECT 1676.550 1319.010 1676.850 1319.390 ;
        RECT 1725.310 1319.390 1773.450 1319.690 ;
        RECT 1676.550 1318.710 1724.690 1319.010 ;
        RECT 1627.790 1318.030 1629.010 1318.330 ;
        RECT 1724.390 1318.330 1724.690 1318.710 ;
        RECT 1725.310 1318.330 1725.610 1319.390 ;
        RECT 1773.150 1319.010 1773.450 1319.390 ;
        RECT 1821.910 1319.390 1870.050 1319.690 ;
        RECT 1773.150 1318.710 1821.290 1319.010 ;
        RECT 1724.390 1318.030 1725.610 1318.330 ;
        RECT 1820.990 1318.330 1821.290 1318.710 ;
        RECT 1821.910 1318.330 1822.210 1319.390 ;
        RECT 1869.750 1319.010 1870.050 1319.390 ;
        RECT 1918.510 1319.390 1966.650 1319.690 ;
        RECT 1869.750 1318.710 1917.890 1319.010 ;
        RECT 1820.990 1318.030 1822.210 1318.330 ;
        RECT 1917.590 1318.330 1917.890 1318.710 ;
        RECT 1918.510 1318.330 1918.810 1319.390 ;
        RECT 1966.350 1319.010 1966.650 1319.390 ;
        RECT 2015.110 1319.390 2063.250 1319.690 ;
        RECT 1966.350 1318.710 2014.490 1319.010 ;
        RECT 1917.590 1318.030 1918.810 1318.330 ;
        RECT 2014.190 1318.330 2014.490 1318.710 ;
        RECT 2015.110 1318.330 2015.410 1319.390 ;
        RECT 2062.950 1319.010 2063.250 1319.390 ;
        RECT 2111.710 1319.390 2159.850 1319.690 ;
        RECT 2062.950 1318.710 2111.090 1319.010 ;
        RECT 2014.190 1318.030 2015.410 1318.330 ;
        RECT 2110.790 1318.330 2111.090 1318.710 ;
        RECT 2111.710 1318.330 2112.010 1319.390 ;
        RECT 2159.550 1319.010 2159.850 1319.390 ;
        RECT 2208.310 1319.390 2256.450 1319.690 ;
        RECT 2159.550 1318.710 2207.690 1319.010 ;
        RECT 2110.790 1318.030 2112.010 1318.330 ;
        RECT 2207.390 1318.330 2207.690 1318.710 ;
        RECT 2208.310 1318.330 2208.610 1319.390 ;
        RECT 2256.150 1319.010 2256.450 1319.390 ;
        RECT 2304.910 1319.390 2353.050 1319.690 ;
        RECT 2256.150 1318.710 2304.290 1319.010 ;
        RECT 2207.390 1318.030 2208.610 1318.330 ;
        RECT 2303.990 1318.330 2304.290 1318.710 ;
        RECT 2304.910 1318.330 2305.210 1319.390 ;
        RECT 2352.750 1319.010 2353.050 1319.390 ;
        RECT 2401.510 1319.390 2449.650 1319.690 ;
        RECT 2352.750 1318.710 2400.890 1319.010 ;
        RECT 2303.990 1318.030 2305.210 1318.330 ;
        RECT 2400.590 1318.330 2400.890 1318.710 ;
        RECT 2401.510 1318.330 2401.810 1319.390 ;
        RECT 2449.350 1319.010 2449.650 1319.390 ;
        RECT 2498.110 1319.390 2546.250 1319.690 ;
        RECT 2449.350 1318.710 2497.490 1319.010 ;
        RECT 2400.590 1318.030 2401.810 1318.330 ;
        RECT 2497.190 1318.330 2497.490 1318.710 ;
        RECT 2498.110 1318.330 2498.410 1319.390 ;
        RECT 2545.950 1319.010 2546.250 1319.390 ;
        RECT 2594.710 1319.390 2642.850 1319.690 ;
        RECT 2545.950 1318.710 2594.090 1319.010 ;
        RECT 2497.190 1318.030 2498.410 1318.330 ;
        RECT 2593.790 1318.330 2594.090 1318.710 ;
        RECT 2594.710 1318.330 2595.010 1319.390 ;
        RECT 2642.550 1319.010 2642.850 1319.390 ;
        RECT 2691.310 1319.390 2739.450 1319.690 ;
        RECT 2642.550 1318.710 2690.690 1319.010 ;
        RECT 2593.790 1318.030 2595.010 1318.330 ;
        RECT 2690.390 1318.330 2690.690 1318.710 ;
        RECT 2691.310 1318.330 2691.610 1319.390 ;
        RECT 2739.150 1319.010 2739.450 1319.390 ;
        RECT 2787.910 1319.390 2836.050 1319.690 ;
        RECT 2739.150 1318.710 2787.290 1319.010 ;
        RECT 2690.390 1318.030 2691.610 1318.330 ;
        RECT 2786.990 1318.330 2787.290 1318.710 ;
        RECT 2787.910 1318.330 2788.210 1319.390 ;
        RECT 2835.750 1319.010 2836.050 1319.390 ;
        RECT 2916.710 1319.390 2924.800 1319.690 ;
        RECT 2916.710 1319.010 2917.010 1319.390 ;
        RECT 2835.750 1318.710 2883.890 1319.010 ;
        RECT 2786.990 1318.030 2788.210 1318.330 ;
        RECT 2883.590 1318.330 2883.890 1318.710 ;
        RECT 2884.510 1318.710 2917.010 1319.010 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
        RECT 2884.510 1318.330 2884.810 1318.710 ;
        RECT 2883.590 1318.030 2884.810 1318.330 ;
        RECT 700.185 1318.015 700.515 1318.030 ;
      LAYER via3 ;
        RECT 284.580 1768.860 284.900 1769.180 ;
        RECT 531.140 1321.420 531.460 1321.740 ;
        RECT 627.740 1320.740 628.060 1321.060 ;
        RECT 434.540 1320.060 434.860 1320.380 ;
        RECT 482.380 1320.060 482.700 1320.380 ;
        RECT 284.580 1319.380 284.900 1319.700 ;
        RECT 482.380 1318.700 482.700 1319.020 ;
        RECT 531.140 1320.060 531.460 1320.380 ;
        RECT 627.740 1319.380 628.060 1319.700 ;
        RECT 434.540 1318.020 434.860 1318.340 ;
      LAYER met4 ;
        RECT 284.575 1768.855 284.905 1769.185 ;
        RECT 284.590 1319.705 284.890 1768.855 ;
        RECT 531.135 1321.415 531.465 1321.745 ;
        RECT 531.150 1320.385 531.450 1321.415 ;
        RECT 627.735 1320.735 628.065 1321.065 ;
        RECT 434.535 1320.055 434.865 1320.385 ;
        RECT 482.375 1320.055 482.705 1320.385 ;
        RECT 531.135 1320.055 531.465 1320.385 ;
        RECT 284.575 1319.375 284.905 1319.705 ;
        RECT 434.550 1318.345 434.850 1320.055 ;
        RECT 482.390 1319.025 482.690 1320.055 ;
        RECT 627.750 1319.705 628.050 1320.735 ;
        RECT 627.735 1319.375 628.065 1319.705 ;
        RECT 482.375 1318.695 482.705 1319.025 ;
        RECT 434.535 1318.015 434.865 1318.345 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 283.430 1559.140 283.750 1559.200 ;
        RECT 2900.830 1559.140 2901.150 1559.200 ;
        RECT 283.430 1559.000 2901.150 1559.140 ;
        RECT 283.430 1558.940 283.750 1559.000 ;
        RECT 2900.830 1558.940 2901.150 1559.000 ;
      LAYER via ;
        RECT 283.460 1558.940 283.720 1559.200 ;
        RECT 2900.860 1558.940 2901.120 1559.200 ;
      LAYER met2 ;
        RECT 283.450 1797.395 283.730 1797.765 ;
        RECT 283.520 1559.230 283.660 1797.395 ;
        RECT 283.460 1558.910 283.720 1559.230 ;
        RECT 2900.860 1558.910 2901.120 1559.230 ;
        RECT 2900.920 1554.325 2901.060 1558.910 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 283.450 1797.440 283.730 1797.720 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 283.425 1797.730 283.755 1797.745 ;
        RECT 300.000 1797.730 304.000 1797.840 ;
        RECT 283.425 1797.430 304.000 1797.730 ;
        RECT 283.425 1797.415 283.755 1797.430 ;
        RECT 300.000 1797.240 304.000 1797.430 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 282.970 1626.800 283.290 1626.860 ;
        RECT 284.350 1626.800 284.670 1626.860 ;
        RECT 282.970 1626.660 284.670 1626.800 ;
        RECT 282.970 1626.600 283.290 1626.660 ;
        RECT 284.350 1626.600 284.670 1626.660 ;
        RECT 282.970 1604.020 283.290 1604.080 ;
        RECT 2904.510 1604.020 2904.830 1604.080 ;
        RECT 282.970 1603.880 2904.830 1604.020 ;
        RECT 282.970 1603.820 283.290 1603.880 ;
        RECT 2904.510 1603.820 2904.830 1603.880 ;
      LAYER via ;
        RECT 283.000 1626.600 283.260 1626.860 ;
        RECT 284.380 1626.600 284.640 1626.860 ;
        RECT 283.000 1603.820 283.260 1604.080 ;
        RECT 2904.540 1603.820 2904.800 1604.080 ;
      LAYER met2 ;
        RECT 285.290 1826.635 285.570 1827.005 ;
        RECT 285.360 1652.810 285.500 1826.635 ;
        RECT 2904.530 1789.235 2904.810 1789.605 ;
        RECT 284.440 1652.670 285.500 1652.810 ;
        RECT 284.440 1626.890 284.580 1652.670 ;
        RECT 283.000 1626.570 283.260 1626.890 ;
        RECT 284.380 1626.570 284.640 1626.890 ;
        RECT 283.060 1604.110 283.200 1626.570 ;
        RECT 2904.600 1604.110 2904.740 1789.235 ;
        RECT 283.000 1603.790 283.260 1604.110 ;
        RECT 2904.540 1603.790 2904.800 1604.110 ;
      LAYER via2 ;
        RECT 285.290 1826.680 285.570 1826.960 ;
        RECT 2904.530 1789.280 2904.810 1789.560 ;
      LAYER met3 ;
        RECT 285.265 1826.970 285.595 1826.985 ;
        RECT 300.000 1826.970 304.000 1827.080 ;
        RECT 285.265 1826.670 304.000 1826.970 ;
        RECT 285.265 1826.655 285.595 1826.670 ;
        RECT 300.000 1826.480 304.000 1826.670 ;
        RECT 2904.505 1789.570 2904.835 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2904.505 1789.270 2924.800 1789.570 ;
        RECT 2904.505 1789.255 2904.835 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 284.810 1654.340 285.130 1654.400 ;
        RECT 299.070 1654.340 299.390 1654.400 ;
        RECT 284.810 1654.200 299.390 1654.340 ;
        RECT 284.810 1654.140 285.130 1654.200 ;
        RECT 299.070 1654.140 299.390 1654.200 ;
        RECT 299.070 1600.280 299.390 1600.340 ;
        RECT 2903.130 1600.280 2903.450 1600.340 ;
        RECT 299.070 1600.140 2903.450 1600.280 ;
        RECT 299.070 1600.080 299.390 1600.140 ;
        RECT 2903.130 1600.080 2903.450 1600.140 ;
      LAYER via ;
        RECT 284.840 1654.140 285.100 1654.400 ;
        RECT 299.100 1654.140 299.360 1654.400 ;
        RECT 299.100 1600.080 299.360 1600.340 ;
        RECT 2903.160 1600.080 2903.420 1600.340 ;
      LAYER met2 ;
        RECT 2903.150 2023.835 2903.430 2024.205 ;
        RECT 284.830 1855.875 285.110 1856.245 ;
        RECT 284.900 1654.430 285.040 1855.875 ;
        RECT 284.840 1654.110 285.100 1654.430 ;
        RECT 299.100 1654.110 299.360 1654.430 ;
        RECT 299.160 1600.370 299.300 1654.110 ;
        RECT 2903.220 1600.370 2903.360 2023.835 ;
        RECT 299.100 1600.050 299.360 1600.370 ;
        RECT 2903.160 1600.050 2903.420 1600.370 ;
      LAYER via2 ;
        RECT 2903.150 2023.880 2903.430 2024.160 ;
        RECT 284.830 1855.920 285.110 1856.200 ;
      LAYER met3 ;
        RECT 2903.125 2024.170 2903.455 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2903.125 2023.870 2924.800 2024.170 ;
        RECT 2903.125 2023.855 2903.455 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 284.805 1856.210 285.135 1856.225 ;
        RECT 300.000 1856.210 304.000 1856.320 ;
        RECT 284.805 1855.910 304.000 1856.210 ;
        RECT 284.805 1855.895 285.135 1855.910 ;
        RECT 300.000 1855.720 304.000 1855.910 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.950 1683.580 289.270 1683.640 ;
        RECT 298.610 1683.580 298.930 1683.640 ;
        RECT 288.950 1683.440 298.930 1683.580 ;
        RECT 288.950 1683.380 289.270 1683.440 ;
        RECT 298.610 1683.380 298.930 1683.440 ;
        RECT 299.530 1599.600 299.850 1599.660 ;
        RECT 2901.750 1599.600 2902.070 1599.660 ;
        RECT 299.530 1599.460 2902.070 1599.600 ;
        RECT 299.530 1599.400 299.850 1599.460 ;
        RECT 2901.750 1599.400 2902.070 1599.460 ;
      LAYER via ;
        RECT 288.980 1683.380 289.240 1683.640 ;
        RECT 298.640 1683.380 298.900 1683.640 ;
        RECT 299.560 1599.400 299.820 1599.660 ;
        RECT 2901.780 1599.400 2902.040 1599.660 ;
      LAYER met2 ;
        RECT 2901.770 2258.435 2902.050 2258.805 ;
        RECT 288.970 1884.435 289.250 1884.805 ;
        RECT 289.040 1683.670 289.180 1884.435 ;
        RECT 288.980 1683.350 289.240 1683.670 ;
        RECT 298.640 1683.410 298.900 1683.670 ;
        RECT 298.640 1683.350 299.760 1683.410 ;
        RECT 298.700 1683.270 299.760 1683.350 ;
        RECT 299.620 1599.690 299.760 1683.270 ;
        RECT 2901.840 1599.690 2901.980 2258.435 ;
        RECT 299.560 1599.370 299.820 1599.690 ;
        RECT 2901.780 1599.370 2902.040 1599.690 ;
      LAYER via2 ;
        RECT 2901.770 2258.480 2902.050 2258.760 ;
        RECT 288.970 1884.480 289.250 1884.760 ;
      LAYER met3 ;
        RECT 2901.745 2258.770 2902.075 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2901.745 2258.470 2924.800 2258.770 ;
        RECT 2901.745 2258.455 2902.075 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 288.945 1884.770 289.275 1884.785 ;
        RECT 300.000 1884.770 304.000 1884.880 ;
        RECT 288.945 1884.470 304.000 1884.770 ;
        RECT 288.945 1884.455 289.275 1884.470 ;
        RECT 300.000 1884.280 304.000 1884.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 687.310 25.740 687.630 25.800 ;
        RECT 1331.770 25.740 1332.090 25.800 ;
        RECT 687.310 25.600 1332.090 25.740 ;
        RECT 687.310 25.540 687.630 25.600 ;
        RECT 1331.770 25.540 1332.090 25.600 ;
        RECT 635.330 24.380 635.650 24.440 ;
        RECT 687.310 24.380 687.630 24.440 ;
        RECT 635.330 24.240 687.630 24.380 ;
        RECT 635.330 24.180 635.650 24.240 ;
        RECT 687.310 24.180 687.630 24.240 ;
      LAYER via ;
        RECT 687.340 25.540 687.600 25.800 ;
        RECT 1331.800 25.540 1332.060 25.800 ;
        RECT 635.360 24.180 635.620 24.440 ;
        RECT 687.340 24.180 687.600 24.440 ;
      LAYER met2 ;
        RECT 1336.010 1600.450 1336.290 1604.000 ;
        RECT 1331.860 1600.310 1336.290 1600.450 ;
        RECT 1331.860 25.830 1332.000 1600.310 ;
        RECT 1336.010 1600.000 1336.290 1600.310 ;
        RECT 687.340 25.510 687.600 25.830 ;
        RECT 1331.800 25.510 1332.060 25.830 ;
        RECT 687.400 24.470 687.540 25.510 ;
        RECT 635.360 24.150 635.620 24.470 ;
        RECT 687.340 24.150 687.600 24.470 ;
        RECT 635.420 23.530 635.560 24.150 ;
        RECT 633.120 23.390 635.560 23.530 ;
        RECT 633.120 2.400 633.260 23.390 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 25.400 651.290 25.460 ;
        RECT 650.970 25.260 686.620 25.400 ;
        RECT 650.970 25.200 651.290 25.260 ;
        RECT 686.480 25.060 686.620 25.260 ;
        RECT 1359.370 25.060 1359.690 25.120 ;
        RECT 686.480 24.920 1359.690 25.060 ;
        RECT 1359.370 24.860 1359.690 24.920 ;
      LAYER via ;
        RECT 651.000 25.200 651.260 25.460 ;
        RECT 1359.400 24.860 1359.660 25.120 ;
      LAYER met2 ;
        RECT 1365.450 1600.450 1365.730 1604.000 ;
        RECT 1359.460 1600.310 1365.730 1600.450 ;
        RECT 651.000 25.170 651.260 25.490 ;
        RECT 651.060 2.400 651.200 25.170 ;
        RECT 1359.460 25.150 1359.600 1600.310 ;
        RECT 1365.450 1600.000 1365.730 1600.310 ;
        RECT 1359.400 24.830 1359.660 25.150 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 639.010 25.740 639.330 25.800 ;
        RECT 639.010 25.600 687.080 25.740 ;
        RECT 639.010 25.540 639.330 25.600 ;
        RECT 686.940 25.400 687.080 25.600 ;
        RECT 1345.570 25.400 1345.890 25.460 ;
        RECT 686.940 25.260 1345.890 25.400 ;
        RECT 1345.570 25.200 1345.890 25.260 ;
      LAYER via ;
        RECT 639.040 25.540 639.300 25.800 ;
        RECT 1345.600 25.200 1345.860 25.460 ;
      LAYER met2 ;
        RECT 1346.130 1600.450 1346.410 1604.000 ;
        RECT 1345.660 1600.310 1346.410 1600.450 ;
        RECT 639.040 25.510 639.300 25.830 ;
        RECT 639.100 2.400 639.240 25.510 ;
        RECT 1345.660 25.490 1345.800 1600.310 ;
        RECT 1346.130 1600.000 1346.410 1600.310 ;
        RECT 1345.600 25.170 1345.860 25.490 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.110 1600.450 1375.390 1604.000 ;
        RECT 1373.260 1600.310 1375.390 1600.450 ;
        RECT 1373.260 24.325 1373.400 1600.310 ;
        RECT 1375.110 1600.000 1375.390 1600.310 ;
        RECT 656.970 23.955 657.250 24.325 ;
        RECT 1373.190 23.955 1373.470 24.325 ;
        RECT 657.040 2.400 657.180 23.955 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 656.970 24.000 657.250 24.280 ;
        RECT 1373.190 24.000 1373.470 24.280 ;
      LAYER met3 ;
        RECT 656.945 24.290 657.275 24.305 ;
        RECT 1373.165 24.290 1373.495 24.305 ;
        RECT 656.945 23.990 1373.495 24.290 ;
        RECT 656.945 23.975 657.275 23.990 ;
        RECT 1373.165 23.975 1373.495 23.990 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 674.430 24.040 674.750 24.100 ;
        RECT 1393.870 24.040 1394.190 24.100 ;
        RECT 674.430 23.900 1394.190 24.040 ;
        RECT 674.430 23.840 674.750 23.900 ;
        RECT 1393.870 23.840 1394.190 23.900 ;
      LAYER via ;
        RECT 674.460 23.840 674.720 24.100 ;
        RECT 1393.900 23.840 1394.160 24.100 ;
      LAYER met2 ;
        RECT 1394.430 1600.450 1394.710 1604.000 ;
        RECT 1393.960 1600.310 1394.710 1600.450 ;
        RECT 1393.960 24.130 1394.100 1600.310 ;
        RECT 1394.430 1600.000 1394.710 1600.310 ;
        RECT 674.460 23.810 674.720 24.130 ;
        RECT 1393.900 23.810 1394.160 24.130 ;
        RECT 674.520 2.400 674.660 23.810 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 644.990 24.720 645.310 24.780 ;
        RECT 1352.470 24.720 1352.790 24.780 ;
        RECT 644.990 24.580 1352.790 24.720 ;
        RECT 644.990 24.520 645.310 24.580 ;
        RECT 1352.470 24.520 1352.790 24.580 ;
      LAYER via ;
        RECT 645.020 24.520 645.280 24.780 ;
        RECT 1352.500 24.520 1352.760 24.780 ;
      LAYER met2 ;
        RECT 1355.790 1600.450 1356.070 1604.000 ;
        RECT 1352.560 1600.310 1356.070 1600.450 ;
        RECT 1352.560 24.810 1352.700 1600.310 ;
        RECT 1355.790 1600.000 1356.070 1600.310 ;
        RECT 645.020 24.490 645.280 24.810 ;
        RECT 1352.500 24.490 1352.760 24.810 ;
        RECT 645.080 2.400 645.220 24.490 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 673.050 25.060 673.370 25.120 ;
        RECT 685.930 25.060 686.250 25.120 ;
        RECT 673.050 24.920 686.250 25.060 ;
        RECT 673.050 24.860 673.370 24.920 ;
        RECT 685.930 24.860 686.250 24.920 ;
        RECT 687.770 24.380 688.090 24.440 ;
        RECT 1380.070 24.380 1380.390 24.440 ;
        RECT 687.770 24.240 1380.390 24.380 ;
        RECT 687.770 24.180 688.090 24.240 ;
        RECT 1380.070 24.180 1380.390 24.240 ;
        RECT 662.930 24.040 663.250 24.100 ;
        RECT 673.050 24.040 673.370 24.100 ;
        RECT 662.930 23.900 673.370 24.040 ;
        RECT 662.930 23.840 663.250 23.900 ;
        RECT 673.050 23.840 673.370 23.900 ;
      LAYER via ;
        RECT 673.080 24.860 673.340 25.120 ;
        RECT 685.960 24.860 686.220 25.120 ;
        RECT 687.800 24.180 688.060 24.440 ;
        RECT 1380.100 24.180 1380.360 24.440 ;
        RECT 662.960 23.840 663.220 24.100 ;
        RECT 673.080 23.840 673.340 24.100 ;
      LAYER met2 ;
        RECT 1384.770 1600.450 1385.050 1604.000 ;
        RECT 1380.160 1600.310 1385.050 1600.450 ;
        RECT 673.080 24.830 673.340 25.150 ;
        RECT 685.960 24.830 686.220 25.150 ;
        RECT 673.140 24.130 673.280 24.830 ;
        RECT 662.960 23.810 663.220 24.130 ;
        RECT 673.080 23.810 673.340 24.130 ;
        RECT 663.020 2.400 663.160 23.810 ;
        RECT 686.020 23.530 686.160 24.830 ;
        RECT 1380.160 24.470 1380.300 1600.310 ;
        RECT 1384.770 1600.000 1385.050 1600.310 ;
        RECT 687.800 24.150 688.060 24.470 ;
        RECT 1380.100 24.150 1380.360 24.470 ;
        RECT 687.860 23.530 688.000 24.150 ;
        RECT 686.020 23.390 688.000 23.530 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1442.630 2790.960 1442.950 2791.020 ;
        RECT 1490.010 2790.960 1490.330 2791.020 ;
        RECT 1442.630 2790.820 1490.330 2790.960 ;
        RECT 1442.630 2790.760 1442.950 2790.820 ;
        RECT 1490.010 2790.760 1490.330 2790.820 ;
        RECT 1511.170 2790.960 1511.490 2791.020 ;
        RECT 1566.830 2790.960 1567.150 2791.020 ;
        RECT 1511.170 2790.820 1567.150 2790.960 ;
        RECT 1511.170 2790.760 1511.490 2790.820 ;
        RECT 1566.830 2790.760 1567.150 2790.820 ;
        RECT 1000.570 2790.280 1000.890 2790.340 ;
        RECT 1068.190 2790.280 1068.510 2790.340 ;
        RECT 1000.570 2790.140 1068.510 2790.280 ;
        RECT 1000.570 2790.080 1000.890 2790.140 ;
        RECT 1068.190 2790.080 1068.510 2790.140 ;
        RECT 972.050 2789.940 972.370 2790.000 ;
        RECT 1000.110 2789.940 1000.430 2790.000 ;
        RECT 972.050 2789.800 1000.430 2789.940 ;
        RECT 972.050 2789.740 972.370 2789.800 ;
        RECT 1000.110 2789.740 1000.430 2789.800 ;
        RECT 1490.010 2789.940 1490.330 2790.000 ;
        RECT 1510.710 2789.940 1511.030 2790.000 ;
        RECT 1490.010 2789.800 1511.030 2789.940 ;
        RECT 1490.010 2789.740 1490.330 2789.800 ;
        RECT 1510.710 2789.740 1511.030 2789.800 ;
        RECT 1442.170 2789.260 1442.490 2789.320 ;
        RECT 1441.800 2789.120 1442.490 2789.260 ;
        RECT 1441.800 2788.980 1441.940 2789.120 ;
        RECT 1442.170 2789.060 1442.490 2789.120 ;
        RECT 1068.190 2788.920 1068.510 2788.980 ;
        RECT 1110.510 2788.920 1110.830 2788.980 ;
        RECT 1068.190 2788.780 1110.830 2788.920 ;
        RECT 1068.190 2788.720 1068.510 2788.780 ;
        RECT 1110.510 2788.720 1110.830 2788.780 ;
        RECT 1110.970 2788.920 1111.290 2788.980 ;
        RECT 1145.470 2788.920 1145.790 2788.980 ;
        RECT 1110.970 2788.780 1145.790 2788.920 ;
        RECT 1110.970 2788.720 1111.290 2788.780 ;
        RECT 1145.470 2788.720 1145.790 2788.780 ;
        RECT 1441.710 2788.720 1442.030 2788.980 ;
        RECT 1510.710 2788.920 1511.030 2788.980 ;
        RECT 1511.170 2788.920 1511.490 2788.980 ;
        RECT 1510.710 2788.780 1511.490 2788.920 ;
        RECT 1510.710 2788.720 1511.030 2788.780 ;
        RECT 1511.170 2788.720 1511.490 2788.780 ;
        RECT 1208.030 2788.580 1208.350 2788.640 ;
        RECT 1200.300 2788.440 1208.350 2788.580 ;
        RECT 1193.310 2788.040 1193.630 2788.300 ;
        RECT 1000.110 2787.900 1000.430 2787.960 ;
        RECT 1000.570 2787.900 1000.890 2787.960 ;
        RECT 1000.110 2787.760 1000.890 2787.900 ;
        RECT 1193.400 2787.900 1193.540 2788.040 ;
        RECT 1200.300 2787.900 1200.440 2788.440 ;
        RECT 1208.030 2788.380 1208.350 2788.440 ;
        RECT 1255.410 2788.240 1255.730 2788.300 ;
        RECT 1269.210 2788.240 1269.530 2788.300 ;
        RECT 1255.410 2788.100 1269.530 2788.240 ;
        RECT 1255.410 2788.040 1255.730 2788.100 ;
        RECT 1269.210 2788.040 1269.530 2788.100 ;
        RECT 1269.670 2788.240 1269.990 2788.300 ;
        RECT 1352.010 2788.240 1352.330 2788.300 ;
        RECT 1365.810 2788.240 1366.130 2788.300 ;
        RECT 1269.670 2788.100 1275.880 2788.240 ;
        RECT 1269.670 2788.040 1269.990 2788.100 ;
        RECT 1193.400 2787.760 1200.440 2787.900 ;
        RECT 1275.740 2787.900 1275.880 2788.100 ;
        RECT 1352.010 2788.100 1366.130 2788.240 ;
        RECT 1352.010 2788.040 1352.330 2788.100 ;
        RECT 1365.810 2788.040 1366.130 2788.100 ;
        RECT 1366.270 2788.240 1366.590 2788.300 ;
        RECT 1366.270 2788.100 1372.480 2788.240 ;
        RECT 1366.270 2788.040 1366.590 2788.100 ;
        RECT 1304.170 2787.900 1304.490 2787.960 ;
        RECT 1275.740 2787.760 1304.490 2787.900 ;
        RECT 1372.340 2787.900 1372.480 2788.100 ;
        RECT 1411.810 2787.900 1412.130 2787.960 ;
        RECT 1441.710 2787.900 1442.030 2787.960 ;
        RECT 1372.340 2787.760 1442.030 2787.900 ;
        RECT 1000.110 2787.700 1000.430 2787.760 ;
        RECT 1000.570 2787.700 1000.890 2787.760 ;
        RECT 1304.170 2787.700 1304.490 2787.760 ;
        RECT 1411.810 2787.700 1412.130 2787.760 ;
        RECT 1441.710 2787.700 1442.030 2787.760 ;
        RECT 1411.810 2746.420 1412.130 2746.480 ;
        RECT 1412.270 2746.420 1412.590 2746.480 ;
        RECT 1411.810 2746.280 1412.590 2746.420 ;
        RECT 1411.810 2746.220 1412.130 2746.280 ;
        RECT 1412.270 2746.220 1412.590 2746.280 ;
        RECT 1412.730 2622.120 1413.050 2622.380 ;
        RECT 1412.820 2621.640 1412.960 2622.120 ;
        RECT 1413.190 2621.640 1413.510 2621.700 ;
        RECT 1412.820 2621.500 1413.510 2621.640 ;
        RECT 1413.190 2621.440 1413.510 2621.500 ;
        RECT 1412.730 2573.840 1413.050 2574.100 ;
        RECT 1412.820 2573.700 1412.960 2573.840 ;
        RECT 1413.190 2573.700 1413.510 2573.760 ;
        RECT 1412.820 2573.560 1413.510 2573.700 ;
        RECT 1413.190 2573.500 1413.510 2573.560 ;
        RECT 1412.730 2560.100 1413.050 2560.160 ;
        RECT 1413.190 2560.100 1413.510 2560.160 ;
        RECT 1412.730 2559.960 1413.510 2560.100 ;
        RECT 1412.730 2559.900 1413.050 2559.960 ;
        RECT 1413.190 2559.900 1413.510 2559.960 ;
        RECT 1412.730 2525.560 1413.050 2525.820 ;
        RECT 1412.820 2525.080 1412.960 2525.560 ;
        RECT 1413.190 2525.080 1413.510 2525.140 ;
        RECT 1412.820 2524.940 1413.510 2525.080 ;
        RECT 1413.190 2524.880 1413.510 2524.940 ;
        RECT 1411.810 2487.680 1412.130 2487.740 ;
        RECT 1412.730 2487.680 1413.050 2487.740 ;
        RECT 1411.810 2487.540 1413.050 2487.680 ;
        RECT 1411.810 2487.480 1412.130 2487.540 ;
        RECT 1412.730 2487.480 1413.050 2487.540 ;
        RECT 1412.730 2429.000 1413.050 2429.260 ;
        RECT 1412.820 2428.520 1412.960 2429.000 ;
        RECT 1413.190 2428.520 1413.510 2428.580 ;
        RECT 1412.820 2428.380 1413.510 2428.520 ;
        RECT 1413.190 2428.320 1413.510 2428.380 ;
        RECT 1411.810 2414.920 1412.130 2414.980 ;
        RECT 1413.190 2414.920 1413.510 2414.980 ;
        RECT 1411.810 2414.780 1413.510 2414.920 ;
        RECT 1411.810 2414.720 1412.130 2414.780 ;
        RECT 1413.190 2414.720 1413.510 2414.780 ;
        RECT 1412.730 2332.100 1413.050 2332.360 ;
        RECT 1412.820 2331.960 1412.960 2332.100 ;
        RECT 1413.190 2331.960 1413.510 2332.020 ;
        RECT 1412.820 2331.820 1413.510 2331.960 ;
        RECT 1413.190 2331.760 1413.510 2331.820 ;
        RECT 1411.810 2318.360 1412.130 2318.420 ;
        RECT 1413.190 2318.360 1413.510 2318.420 ;
        RECT 1411.810 2318.220 1413.510 2318.360 ;
        RECT 1411.810 2318.160 1412.130 2318.220 ;
        RECT 1413.190 2318.160 1413.510 2318.220 ;
        RECT 1412.730 2235.540 1413.050 2235.800 ;
        RECT 1412.820 2235.400 1412.960 2235.540 ;
        RECT 1413.190 2235.400 1413.510 2235.460 ;
        RECT 1412.820 2235.260 1413.510 2235.400 ;
        RECT 1413.190 2235.200 1413.510 2235.260 ;
        RECT 1414.110 2173.520 1414.430 2173.580 ;
        RECT 1415.030 2173.520 1415.350 2173.580 ;
        RECT 1414.110 2173.380 1415.350 2173.520 ;
        RECT 1414.110 2173.320 1414.430 2173.380 ;
        RECT 1415.030 2173.320 1415.350 2173.380 ;
        RECT 1413.190 2069.820 1413.510 2069.880 ;
        RECT 2063.170 2069.820 2063.490 2069.880 ;
        RECT 1413.190 2069.680 2063.490 2069.820 ;
        RECT 1413.190 2069.620 1413.510 2069.680 ;
        RECT 2063.170 2069.620 2063.490 2069.680 ;
        RECT 2.830 16.220 3.150 16.280 ;
        RECT 306.890 16.220 307.210 16.280 ;
        RECT 2.830 16.080 307.210 16.220 ;
        RECT 2.830 16.020 3.150 16.080 ;
        RECT 306.890 16.020 307.210 16.080 ;
      LAYER via ;
        RECT 1442.660 2790.760 1442.920 2791.020 ;
        RECT 1490.040 2790.760 1490.300 2791.020 ;
        RECT 1511.200 2790.760 1511.460 2791.020 ;
        RECT 1566.860 2790.760 1567.120 2791.020 ;
        RECT 1000.600 2790.080 1000.860 2790.340 ;
        RECT 1068.220 2790.080 1068.480 2790.340 ;
        RECT 972.080 2789.740 972.340 2790.000 ;
        RECT 1000.140 2789.740 1000.400 2790.000 ;
        RECT 1490.040 2789.740 1490.300 2790.000 ;
        RECT 1510.740 2789.740 1511.000 2790.000 ;
        RECT 1442.200 2789.060 1442.460 2789.320 ;
        RECT 1068.220 2788.720 1068.480 2788.980 ;
        RECT 1110.540 2788.720 1110.800 2788.980 ;
        RECT 1111.000 2788.720 1111.260 2788.980 ;
        RECT 1145.500 2788.720 1145.760 2788.980 ;
        RECT 1441.740 2788.720 1442.000 2788.980 ;
        RECT 1510.740 2788.720 1511.000 2788.980 ;
        RECT 1511.200 2788.720 1511.460 2788.980 ;
        RECT 1193.340 2788.040 1193.600 2788.300 ;
        RECT 1000.140 2787.700 1000.400 2787.960 ;
        RECT 1000.600 2787.700 1000.860 2787.960 ;
        RECT 1208.060 2788.380 1208.320 2788.640 ;
        RECT 1255.440 2788.040 1255.700 2788.300 ;
        RECT 1269.240 2788.040 1269.500 2788.300 ;
        RECT 1269.700 2788.040 1269.960 2788.300 ;
        RECT 1352.040 2788.040 1352.300 2788.300 ;
        RECT 1365.840 2788.040 1366.100 2788.300 ;
        RECT 1366.300 2788.040 1366.560 2788.300 ;
        RECT 1304.200 2787.700 1304.460 2787.960 ;
        RECT 1411.840 2787.700 1412.100 2787.960 ;
        RECT 1441.740 2787.700 1442.000 2787.960 ;
        RECT 1411.840 2746.220 1412.100 2746.480 ;
        RECT 1412.300 2746.220 1412.560 2746.480 ;
        RECT 1412.760 2622.120 1413.020 2622.380 ;
        RECT 1413.220 2621.440 1413.480 2621.700 ;
        RECT 1412.760 2573.840 1413.020 2574.100 ;
        RECT 1413.220 2573.500 1413.480 2573.760 ;
        RECT 1412.760 2559.900 1413.020 2560.160 ;
        RECT 1413.220 2559.900 1413.480 2560.160 ;
        RECT 1412.760 2525.560 1413.020 2525.820 ;
        RECT 1413.220 2524.880 1413.480 2525.140 ;
        RECT 1411.840 2487.480 1412.100 2487.740 ;
        RECT 1412.760 2487.480 1413.020 2487.740 ;
        RECT 1412.760 2429.000 1413.020 2429.260 ;
        RECT 1413.220 2428.320 1413.480 2428.580 ;
        RECT 1411.840 2414.720 1412.100 2414.980 ;
        RECT 1413.220 2414.720 1413.480 2414.980 ;
        RECT 1412.760 2332.100 1413.020 2332.360 ;
        RECT 1413.220 2331.760 1413.480 2332.020 ;
        RECT 1411.840 2318.160 1412.100 2318.420 ;
        RECT 1413.220 2318.160 1413.480 2318.420 ;
        RECT 1412.760 2235.540 1413.020 2235.800 ;
        RECT 1413.220 2235.200 1413.480 2235.460 ;
        RECT 1414.140 2173.320 1414.400 2173.580 ;
        RECT 1415.060 2173.320 1415.320 2173.580 ;
        RECT 1413.220 2069.620 1413.480 2069.880 ;
        RECT 2063.200 2069.620 2063.460 2069.880 ;
        RECT 2.860 16.020 3.120 16.280 ;
        RECT 306.920 16.020 307.180 16.280 ;
      LAYER met2 ;
        RECT 1566.850 2794.275 1567.130 2794.645 ;
        RECT 972.070 2793.595 972.350 2793.965 ;
        RECT 972.140 2790.030 972.280 2793.595 ;
        RECT 1566.920 2791.050 1567.060 2794.275 ;
        RECT 1442.660 2790.730 1442.920 2791.050 ;
        RECT 1490.040 2790.730 1490.300 2791.050 ;
        RECT 1511.200 2790.730 1511.460 2791.050 ;
        RECT 1566.860 2790.730 1567.120 2791.050 ;
        RECT 1000.600 2790.050 1000.860 2790.370 ;
        RECT 1068.220 2790.050 1068.480 2790.370 ;
        RECT 972.080 2789.710 972.340 2790.030 ;
        RECT 1000.140 2789.710 1000.400 2790.030 ;
        RECT 1000.200 2787.990 1000.340 2789.710 ;
        RECT 1000.660 2787.990 1000.800 2790.050 ;
        RECT 1068.280 2789.010 1068.420 2790.050 ;
        RECT 1110.600 2789.010 1111.200 2789.090 ;
        RECT 1068.220 2788.690 1068.480 2789.010 ;
        RECT 1110.540 2788.950 1111.260 2789.010 ;
        RECT 1110.540 2788.690 1110.800 2788.950 ;
        RECT 1111.000 2788.690 1111.260 2788.950 ;
        RECT 1145.490 2788.835 1145.770 2789.205 ;
        RECT 1193.330 2788.835 1193.610 2789.205 ;
        RECT 1442.200 2789.090 1442.460 2789.350 ;
        RECT 1442.720 2789.090 1442.860 2790.730 ;
        RECT 1490.100 2790.030 1490.240 2790.730 ;
        RECT 1490.040 2789.710 1490.300 2790.030 ;
        RECT 1510.740 2789.710 1511.000 2790.030 ;
        RECT 1442.200 2789.030 1442.860 2789.090 ;
        RECT 1145.500 2788.690 1145.760 2788.835 ;
        RECT 1193.400 2788.330 1193.540 2788.835 ;
        RECT 1441.740 2788.690 1442.000 2789.010 ;
        RECT 1442.260 2788.950 1442.860 2789.030 ;
        RECT 1510.800 2789.010 1510.940 2789.710 ;
        RECT 1511.260 2789.010 1511.400 2790.730 ;
        RECT 1510.740 2788.690 1511.000 2789.010 ;
        RECT 1511.200 2788.690 1511.460 2789.010 ;
        RECT 1208.060 2788.350 1208.320 2788.670 ;
        RECT 1193.340 2788.010 1193.600 2788.330 ;
        RECT 1000.140 2787.670 1000.400 2787.990 ;
        RECT 1000.600 2787.670 1000.860 2787.990 ;
        RECT 1208.120 2787.845 1208.260 2788.350 ;
        RECT 1269.300 2788.330 1269.900 2788.410 ;
        RECT 1365.900 2788.330 1366.500 2788.410 ;
        RECT 1255.440 2788.010 1255.700 2788.330 ;
        RECT 1269.240 2788.270 1269.960 2788.330 ;
        RECT 1269.240 2788.010 1269.500 2788.270 ;
        RECT 1269.700 2788.010 1269.960 2788.270 ;
        RECT 1352.040 2788.010 1352.300 2788.330 ;
        RECT 1365.840 2788.270 1366.560 2788.330 ;
        RECT 1365.840 2788.010 1366.100 2788.270 ;
        RECT 1366.300 2788.010 1366.560 2788.270 ;
        RECT 1255.500 2787.845 1255.640 2788.010 ;
        RECT 1304.200 2787.845 1304.460 2787.990 ;
        RECT 1352.100 2787.845 1352.240 2788.010 ;
        RECT 1441.800 2787.990 1441.940 2788.690 ;
        RECT 1208.050 2787.475 1208.330 2787.845 ;
        RECT 1255.430 2787.475 1255.710 2787.845 ;
        RECT 1304.190 2787.475 1304.470 2787.845 ;
        RECT 1352.030 2787.475 1352.310 2787.845 ;
        RECT 1411.840 2787.670 1412.100 2787.990 ;
        RECT 1441.740 2787.670 1442.000 2787.990 ;
        RECT 1411.900 2746.510 1412.040 2787.670 ;
        RECT 1411.840 2746.190 1412.100 2746.510 ;
        RECT 1412.300 2746.190 1412.560 2746.510 ;
        RECT 1412.360 2697.970 1412.500 2746.190 ;
        RECT 1412.360 2697.830 1412.960 2697.970 ;
        RECT 1412.820 2622.410 1412.960 2697.830 ;
        RECT 1412.760 2622.090 1413.020 2622.410 ;
        RECT 1413.220 2621.410 1413.480 2621.730 ;
        RECT 1413.280 2608.210 1413.420 2621.410 ;
        RECT 1412.820 2608.070 1413.420 2608.210 ;
        RECT 1412.820 2574.130 1412.960 2608.070 ;
        RECT 1412.760 2573.810 1413.020 2574.130 ;
        RECT 1413.220 2573.470 1413.480 2573.790 ;
        RECT 1413.280 2560.190 1413.420 2573.470 ;
        RECT 1412.760 2559.870 1413.020 2560.190 ;
        RECT 1413.220 2559.870 1413.480 2560.190 ;
        RECT 1412.820 2525.850 1412.960 2559.870 ;
        RECT 1412.760 2525.530 1413.020 2525.850 ;
        RECT 1413.220 2524.850 1413.480 2525.170 ;
        RECT 1413.280 2511.650 1413.420 2524.850 ;
        RECT 1412.820 2511.510 1413.420 2511.650 ;
        RECT 1412.820 2487.770 1412.960 2511.510 ;
        RECT 1411.840 2487.450 1412.100 2487.770 ;
        RECT 1412.760 2487.450 1413.020 2487.770 ;
        RECT 1411.900 2463.485 1412.040 2487.450 ;
        RECT 1411.830 2463.115 1412.110 2463.485 ;
        RECT 1412.750 2463.115 1413.030 2463.485 ;
        RECT 1412.820 2429.290 1412.960 2463.115 ;
        RECT 1412.760 2428.970 1413.020 2429.290 ;
        RECT 1413.220 2428.290 1413.480 2428.610 ;
        RECT 1413.280 2415.010 1413.420 2428.290 ;
        RECT 1411.840 2414.690 1412.100 2415.010 ;
        RECT 1413.220 2414.690 1413.480 2415.010 ;
        RECT 1411.900 2366.925 1412.040 2414.690 ;
        RECT 1411.830 2366.555 1412.110 2366.925 ;
        RECT 1412.750 2366.555 1413.030 2366.925 ;
        RECT 1412.820 2332.390 1412.960 2366.555 ;
        RECT 1412.760 2332.070 1413.020 2332.390 ;
        RECT 1413.220 2331.730 1413.480 2332.050 ;
        RECT 1413.280 2318.450 1413.420 2331.730 ;
        RECT 1411.840 2318.130 1412.100 2318.450 ;
        RECT 1413.220 2318.130 1413.480 2318.450 ;
        RECT 1411.900 2270.365 1412.040 2318.130 ;
        RECT 1411.830 2269.995 1412.110 2270.365 ;
        RECT 1412.750 2269.995 1413.030 2270.365 ;
        RECT 1412.820 2235.830 1412.960 2269.995 ;
        RECT 1412.760 2235.510 1413.020 2235.830 ;
        RECT 1413.220 2235.170 1413.480 2235.490 ;
        RECT 1413.280 2187.290 1413.420 2235.170 ;
        RECT 1413.280 2187.150 1414.340 2187.290 ;
        RECT 1414.200 2173.610 1414.340 2187.150 ;
        RECT 1414.140 2173.290 1414.400 2173.610 ;
        RECT 1415.060 2173.290 1415.320 2173.610 ;
        RECT 1415.120 2125.525 1415.260 2173.290 ;
        RECT 1413.210 2125.155 1413.490 2125.525 ;
        RECT 1415.050 2125.155 1415.330 2125.525 ;
        RECT 1413.280 2069.910 1413.420 2125.155 ;
        RECT 1413.220 2069.765 1413.480 2069.910 ;
        RECT 1413.210 2069.395 1413.490 2069.765 ;
        RECT 2063.200 2069.590 2063.460 2069.910 ;
        RECT 1413.280 2069.265 1413.420 2069.395 ;
        RECT 2063.260 2069.085 2063.400 2069.590 ;
        RECT 2063.190 2068.715 2063.470 2069.085 ;
        RECT 304.690 1600.450 304.970 1604.000 ;
        RECT 304.690 1600.310 307.120 1600.450 ;
        RECT 304.690 1600.000 304.970 1600.310 ;
        RECT 306.980 1586.965 307.120 1600.310 ;
        RECT 306.910 1586.595 307.190 1586.965 ;
        RECT 306.980 16.310 307.120 1586.595 ;
        RECT 2.860 15.990 3.120 16.310 ;
        RECT 306.920 15.990 307.180 16.310 ;
        RECT 2.920 2.400 3.060 15.990 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 1566.850 2794.320 1567.130 2794.600 ;
        RECT 972.070 2793.640 972.350 2793.920 ;
        RECT 1145.490 2788.880 1145.770 2789.160 ;
        RECT 1193.330 2788.880 1193.610 2789.160 ;
        RECT 1208.050 2787.520 1208.330 2787.800 ;
        RECT 1255.430 2787.520 1255.710 2787.800 ;
        RECT 1304.190 2787.520 1304.470 2787.800 ;
        RECT 1352.030 2787.520 1352.310 2787.800 ;
        RECT 1411.830 2463.160 1412.110 2463.440 ;
        RECT 1412.750 2463.160 1413.030 2463.440 ;
        RECT 1411.830 2366.600 1412.110 2366.880 ;
        RECT 1412.750 2366.600 1413.030 2366.880 ;
        RECT 1411.830 2270.040 1412.110 2270.320 ;
        RECT 1412.750 2270.040 1413.030 2270.320 ;
        RECT 1413.210 2125.200 1413.490 2125.480 ;
        RECT 1415.050 2125.200 1415.330 2125.480 ;
        RECT 1413.210 2069.440 1413.490 2069.720 ;
        RECT 2063.190 2068.760 2063.470 2069.040 ;
        RECT 306.910 1586.640 307.190 1586.920 ;
      LAYER met3 ;
        RECT 1566.825 2794.620 1567.155 2794.625 ;
        RECT 1566.825 2794.610 1567.410 2794.620 ;
        RECT 1566.825 2794.310 1567.610 2794.610 ;
        RECT 1566.825 2794.300 1567.410 2794.310 ;
        RECT 1566.825 2794.295 1567.155 2794.300 ;
        RECT 972.045 2793.940 972.375 2793.945 ;
        RECT 321.350 2793.930 321.730 2793.940 ;
        RECT 971.790 2793.930 972.375 2793.940 ;
        RECT 321.350 2793.630 972.375 2793.930 ;
        RECT 321.350 2793.620 321.730 2793.630 ;
        RECT 971.790 2793.620 972.375 2793.630 ;
        RECT 972.045 2793.615 972.375 2793.620 ;
        RECT 1145.465 2789.170 1145.795 2789.185 ;
        RECT 1193.305 2789.170 1193.635 2789.185 ;
        RECT 1145.465 2788.870 1193.635 2789.170 ;
        RECT 1145.465 2788.855 1145.795 2788.870 ;
        RECT 1193.305 2788.855 1193.635 2788.870 ;
        RECT 1208.025 2787.810 1208.355 2787.825 ;
        RECT 1255.405 2787.810 1255.735 2787.825 ;
        RECT 1208.025 2787.510 1255.735 2787.810 ;
        RECT 1208.025 2787.495 1208.355 2787.510 ;
        RECT 1255.405 2787.495 1255.735 2787.510 ;
        RECT 1304.165 2787.810 1304.495 2787.825 ;
        RECT 1352.005 2787.810 1352.335 2787.825 ;
        RECT 1304.165 2787.510 1352.335 2787.810 ;
        RECT 1304.165 2787.495 1304.495 2787.510 ;
        RECT 1352.005 2787.495 1352.335 2787.510 ;
        RECT 1411.805 2463.450 1412.135 2463.465 ;
        RECT 1412.725 2463.450 1413.055 2463.465 ;
        RECT 1411.805 2463.150 1413.055 2463.450 ;
        RECT 1411.805 2463.135 1412.135 2463.150 ;
        RECT 1412.725 2463.135 1413.055 2463.150 ;
        RECT 1411.805 2366.890 1412.135 2366.905 ;
        RECT 1412.725 2366.890 1413.055 2366.905 ;
        RECT 1411.805 2366.590 1413.055 2366.890 ;
        RECT 1411.805 2366.575 1412.135 2366.590 ;
        RECT 1412.725 2366.575 1413.055 2366.590 ;
        RECT 1411.805 2270.330 1412.135 2270.345 ;
        RECT 1412.725 2270.330 1413.055 2270.345 ;
        RECT 1411.805 2270.030 1413.055 2270.330 ;
        RECT 1411.805 2270.015 1412.135 2270.030 ;
        RECT 1412.725 2270.015 1413.055 2270.030 ;
        RECT 1413.185 2125.490 1413.515 2125.505 ;
        RECT 1415.025 2125.490 1415.355 2125.505 ;
        RECT 1413.185 2125.190 1415.355 2125.490 ;
        RECT 1413.185 2125.175 1413.515 2125.190 ;
        RECT 1415.025 2125.175 1415.355 2125.190 ;
        RECT 1407.870 2069.730 1408.250 2069.740 ;
        RECT 1413.185 2069.730 1413.515 2069.745 ;
        RECT 1407.870 2069.430 1413.515 2069.730 ;
        RECT 1407.870 2069.420 1408.250 2069.430 ;
        RECT 1413.185 2069.415 1413.515 2069.430 ;
        RECT 2063.165 2069.050 2063.495 2069.065 ;
        RECT 2063.830 2069.050 2064.210 2069.060 ;
        RECT 2063.165 2068.750 2064.210 2069.050 ;
        RECT 2063.165 2068.735 2063.495 2068.750 ;
        RECT 2063.830 2068.740 2064.210 2068.750 ;
        RECT 306.885 1586.930 307.215 1586.945 ;
        RECT 1407.870 1586.930 1408.250 1586.940 ;
        RECT 306.885 1586.630 1408.250 1586.930 ;
        RECT 306.885 1586.615 307.215 1586.630 ;
        RECT 1407.870 1586.620 1408.250 1586.630 ;
      LAYER via3 ;
        RECT 1567.060 2794.300 1567.380 2794.620 ;
        RECT 321.380 2793.620 321.700 2793.940 ;
        RECT 971.820 2793.620 972.140 2793.940 ;
        RECT 1407.900 2069.420 1408.220 2069.740 ;
        RECT 2063.860 2068.740 2064.180 2069.060 ;
        RECT 1407.900 1586.620 1408.220 1586.940 ;
      LAYER met4 ;
        RECT 319.015 2801.750 319.315 2804.600 ;
        RECT 969.015 2801.750 969.315 2804.600 ;
        RECT 1569.015 2801.750 1569.315 2804.600 ;
        RECT 319.015 2801.450 321.690 2801.750 ;
        RECT 319.015 2800.000 319.315 2801.450 ;
        RECT 321.390 2793.945 321.690 2801.450 ;
        RECT 969.015 2801.450 972.130 2801.750 ;
        RECT 969.015 2800.000 969.315 2801.450 ;
        RECT 971.830 2793.945 972.130 2801.450 ;
        RECT 1567.070 2801.450 1569.315 2801.750 ;
        RECT 1567.070 2794.625 1567.370 2801.450 ;
        RECT 1569.015 2800.000 1569.315 2801.450 ;
        RECT 1567.055 2794.295 1567.385 2794.625 ;
        RECT 321.375 2793.615 321.705 2793.945 ;
        RECT 971.815 2793.615 972.145 2793.945 ;
        RECT 1407.895 2069.415 1408.225 2069.745 ;
        RECT 1407.910 1586.945 1408.210 2069.415 ;
        RECT 2063.855 2068.735 2064.185 2069.065 ;
        RECT 2063.870 2055.450 2064.170 2068.735 ;
        RECT 2067.165 2055.450 2067.465 2056.235 ;
        RECT 2063.870 2055.150 2067.465 2055.450 ;
        RECT 2067.165 2051.635 2067.465 2055.150 ;
        RECT 1407.895 1586.615 1408.225 1586.945 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.410 1589.400 13.730 1589.460 ;
        RECT 314.250 1589.400 314.570 1589.460 ;
        RECT 13.410 1589.260 314.570 1589.400 ;
        RECT 13.410 1589.200 13.730 1589.260 ;
        RECT 314.250 1589.200 314.570 1589.260 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 1589.200 13.700 1589.460 ;
        RECT 314.280 1589.200 314.540 1589.460 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 314.350 1600.380 314.630 1604.000 ;
        RECT 314.340 1600.000 314.630 1600.380 ;
        RECT 314.340 1589.490 314.480 1600.000 ;
        RECT 13.440 1589.170 13.700 1589.490 ;
        RECT 314.280 1589.170 314.540 1589.490 ;
        RECT 13.500 17.670 13.640 1589.170 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 1593.820 20.630 1593.880 ;
        RECT 323.910 1593.820 324.230 1593.880 ;
        RECT 20.310 1593.680 324.230 1593.820 ;
        RECT 20.310 1593.620 20.630 1593.680 ;
        RECT 323.910 1593.620 324.230 1593.680 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 20.310 17.580 20.630 17.640 ;
        RECT 14.330 17.440 20.630 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 20.310 17.380 20.630 17.440 ;
      LAYER via ;
        RECT 20.340 1593.620 20.600 1593.880 ;
        RECT 323.940 1593.620 324.200 1593.880 ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 20.340 17.380 20.600 17.640 ;
      LAYER met2 ;
        RECT 324.010 1600.380 324.290 1604.000 ;
        RECT 324.000 1600.000 324.290 1600.380 ;
        RECT 324.000 1593.910 324.140 1600.000 ;
        RECT 20.340 1593.590 20.600 1593.910 ;
        RECT 323.940 1593.590 324.200 1593.910 ;
        RECT 20.400 17.670 20.540 1593.590 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 20.340 17.350 20.600 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 1593.140 41.330 1593.200 ;
        RECT 362.550 1593.140 362.870 1593.200 ;
        RECT 41.010 1593.000 362.870 1593.140 ;
        RECT 41.010 1592.940 41.330 1593.000 ;
        RECT 362.550 1592.940 362.870 1593.000 ;
        RECT 38.250 17.580 38.570 17.640 ;
        RECT 41.010 17.580 41.330 17.640 ;
        RECT 38.250 17.440 41.330 17.580 ;
        RECT 38.250 17.380 38.570 17.440 ;
        RECT 41.010 17.380 41.330 17.440 ;
      LAYER via ;
        RECT 41.040 1592.940 41.300 1593.200 ;
        RECT 362.580 1592.940 362.840 1593.200 ;
        RECT 38.280 17.380 38.540 17.640 ;
        RECT 41.040 17.380 41.300 17.640 ;
      LAYER met2 ;
        RECT 362.650 1600.380 362.930 1604.000 ;
        RECT 362.640 1600.000 362.930 1600.380 ;
        RECT 362.640 1593.230 362.780 1600.000 ;
        RECT 41.040 1592.910 41.300 1593.230 ;
        RECT 362.580 1592.910 362.840 1593.230 ;
        RECT 41.100 17.670 41.240 1592.910 ;
        RECT 38.280 17.350 38.540 17.670 ;
        RECT 41.040 17.350 41.300 17.670 ;
        RECT 38.340 2.400 38.480 17.350 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 20.980 241.430 21.040 ;
        RECT 690.070 20.980 690.390 21.040 ;
        RECT 241.110 20.840 690.390 20.980 ;
        RECT 241.110 20.780 241.430 20.840 ;
        RECT 690.070 20.780 690.390 20.840 ;
      LAYER via ;
        RECT 241.140 20.780 241.400 21.040 ;
        RECT 690.100 20.780 690.360 21.040 ;
      LAYER met2 ;
        RECT 693.850 1600.450 694.130 1604.000 ;
        RECT 690.160 1600.310 694.130 1600.450 ;
        RECT 690.160 21.070 690.300 1600.310 ;
        RECT 693.850 1600.000 694.130 1600.310 ;
        RECT 241.140 20.750 241.400 21.070 ;
        RECT 690.100 20.750 690.360 21.070 ;
        RECT 241.200 10.610 241.340 20.750 ;
        RECT 240.740 10.470 241.340 10.610 ;
        RECT 240.740 2.400 240.880 10.470 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 258.130 21.320 258.450 21.380 ;
        RECT 717.670 21.320 717.990 21.380 ;
        RECT 258.130 21.180 717.990 21.320 ;
        RECT 258.130 21.120 258.450 21.180 ;
        RECT 717.670 21.120 717.990 21.180 ;
      LAYER via ;
        RECT 258.160 21.120 258.420 21.380 ;
        RECT 717.700 21.120 717.960 21.380 ;
      LAYER met2 ;
        RECT 722.830 1600.450 723.110 1604.000 ;
        RECT 717.760 1600.310 723.110 1600.450 ;
        RECT 717.760 21.410 717.900 1600.310 ;
        RECT 722.830 1600.000 723.110 1600.310 ;
        RECT 258.160 21.090 258.420 21.410 ;
        RECT 717.700 21.090 717.960 21.410 ;
        RECT 258.220 2.400 258.360 21.090 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 276.070 21.660 276.390 21.720 ;
        RECT 752.170 21.660 752.490 21.720 ;
        RECT 276.070 21.520 752.490 21.660 ;
        RECT 276.070 21.460 276.390 21.520 ;
        RECT 752.170 21.460 752.490 21.520 ;
      LAYER via ;
        RECT 276.100 21.460 276.360 21.720 ;
        RECT 752.200 21.460 752.460 21.720 ;
      LAYER met2 ;
        RECT 752.270 1600.380 752.550 1604.000 ;
        RECT 752.260 1600.000 752.550 1600.380 ;
        RECT 752.260 21.750 752.400 1600.000 ;
        RECT 276.100 21.430 276.360 21.750 ;
        RECT 752.200 21.430 752.460 21.750 ;
        RECT 276.160 2.400 276.300 21.430 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 22.000 294.330 22.060 ;
        RECT 779.770 22.000 780.090 22.060 ;
        RECT 294.010 21.860 780.090 22.000 ;
        RECT 294.010 21.800 294.330 21.860 ;
        RECT 779.770 21.800 780.090 21.860 ;
      LAYER via ;
        RECT 294.040 21.800 294.300 22.060 ;
        RECT 779.800 21.800 780.060 22.060 ;
      LAYER met2 ;
        RECT 781.250 1600.450 781.530 1604.000 ;
        RECT 779.860 1600.310 781.530 1600.450 ;
        RECT 779.860 22.090 780.000 1600.310 ;
        RECT 781.250 1600.000 781.530 1600.310 ;
        RECT 294.040 21.770 294.300 22.090 ;
        RECT 779.800 21.770 780.060 22.090 ;
        RECT 294.100 2.400 294.240 21.770 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 22.340 312.270 22.400 ;
        RECT 807.370 22.340 807.690 22.400 ;
        RECT 311.950 22.200 807.690 22.340 ;
        RECT 311.950 22.140 312.270 22.200 ;
        RECT 807.370 22.140 807.690 22.200 ;
      LAYER via ;
        RECT 311.980 22.140 312.240 22.400 ;
        RECT 807.400 22.140 807.660 22.400 ;
      LAYER met2 ;
        RECT 810.690 1600.450 810.970 1604.000 ;
        RECT 807.460 1600.310 810.970 1600.450 ;
        RECT 807.460 22.430 807.600 1600.310 ;
        RECT 810.690 1600.000 810.970 1600.310 ;
        RECT 311.980 22.110 312.240 22.430 ;
        RECT 807.400 22.110 807.660 22.430 ;
        RECT 312.040 2.400 312.180 22.110 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 22.680 330.210 22.740 ;
        RECT 834.970 22.680 835.290 22.740 ;
        RECT 329.890 22.540 835.290 22.680 ;
        RECT 329.890 22.480 330.210 22.540 ;
        RECT 834.970 22.480 835.290 22.540 ;
      LAYER via ;
        RECT 329.920 22.480 330.180 22.740 ;
        RECT 835.000 22.480 835.260 22.740 ;
      LAYER met2 ;
        RECT 839.670 1600.450 839.950 1604.000 ;
        RECT 835.060 1600.310 839.950 1600.450 ;
        RECT 835.060 22.770 835.200 1600.310 ;
        RECT 839.670 1600.000 839.950 1600.310 ;
        RECT 329.920 22.450 330.180 22.770 ;
        RECT 835.000 22.450 835.260 22.770 ;
        RECT 329.980 2.400 330.120 22.450 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 23.020 347.690 23.080 ;
        RECT 862.570 23.020 862.890 23.080 ;
        RECT 347.370 22.880 862.890 23.020 ;
        RECT 347.370 22.820 347.690 22.880 ;
        RECT 862.570 22.820 862.890 22.880 ;
      LAYER via ;
        RECT 347.400 22.820 347.660 23.080 ;
        RECT 862.600 22.820 862.860 23.080 ;
      LAYER met2 ;
        RECT 869.110 1600.450 869.390 1604.000 ;
        RECT 862.660 1600.310 869.390 1600.450 ;
        RECT 862.660 23.110 862.800 1600.310 ;
        RECT 869.110 1600.000 869.390 1600.310 ;
        RECT 347.400 22.790 347.660 23.110 ;
        RECT 862.600 22.790 862.860 23.110 ;
        RECT 347.460 2.400 347.600 22.790 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 23.360 365.630 23.420 ;
        RECT 897.070 23.360 897.390 23.420 ;
        RECT 365.310 23.220 897.390 23.360 ;
        RECT 365.310 23.160 365.630 23.220 ;
        RECT 897.070 23.160 897.390 23.220 ;
      LAYER via ;
        RECT 365.340 23.160 365.600 23.420 ;
        RECT 897.100 23.160 897.360 23.420 ;
      LAYER met2 ;
        RECT 898.090 1600.450 898.370 1604.000 ;
        RECT 897.160 1600.310 898.370 1600.450 ;
        RECT 897.160 23.450 897.300 1600.310 ;
        RECT 898.090 1600.000 898.370 1600.310 ;
        RECT 365.340 23.130 365.600 23.450 ;
        RECT 897.100 23.130 897.360 23.450 ;
        RECT 365.400 21.490 365.540 23.130 ;
        RECT 365.400 21.350 366.000 21.490 ;
        RECT 365.860 20.130 366.000 21.350 ;
        RECT 365.400 19.990 366.000 20.130 ;
        RECT 365.400 2.400 365.540 19.990 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 23.700 383.570 23.760 ;
        RECT 924.670 23.700 924.990 23.760 ;
        RECT 383.250 23.560 924.990 23.700 ;
        RECT 383.250 23.500 383.570 23.560 ;
        RECT 924.670 23.500 924.990 23.560 ;
      LAYER via ;
        RECT 383.280 23.500 383.540 23.760 ;
        RECT 924.700 23.500 924.960 23.760 ;
      LAYER met2 ;
        RECT 927.530 1600.450 927.810 1604.000 ;
        RECT 924.760 1600.310 927.810 1600.450 ;
        RECT 924.760 23.790 924.900 1600.310 ;
        RECT 927.530 1600.000 927.810 1600.310 ;
        RECT 383.280 23.470 383.540 23.790 ;
        RECT 924.700 23.470 924.960 23.790 ;
        RECT 383.340 2.400 383.480 23.470 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 27.440 401.510 27.500 ;
        RECT 952.270 27.440 952.590 27.500 ;
        RECT 401.190 27.300 952.590 27.440 ;
        RECT 401.190 27.240 401.510 27.300 ;
        RECT 952.270 27.240 952.590 27.300 ;
      LAYER via ;
        RECT 401.220 27.240 401.480 27.500 ;
        RECT 952.300 27.240 952.560 27.500 ;
      LAYER met2 ;
        RECT 956.510 1600.450 956.790 1604.000 ;
        RECT 952.360 1600.310 956.790 1600.450 ;
        RECT 952.360 27.530 952.500 1600.310 ;
        RECT 956.510 1600.000 956.790 1600.310 ;
        RECT 401.220 27.210 401.480 27.530 ;
        RECT 952.300 27.210 952.560 27.530 ;
        RECT 401.280 2.400 401.420 27.210 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 400.270 27.440 400.590 27.500 ;
        RECT 393.460 27.300 400.590 27.440 ;
        RECT 62.170 26.760 62.490 26.820 ;
        RECT 393.460 26.760 393.600 27.300 ;
        RECT 400.270 27.240 400.590 27.300 ;
        RECT 62.170 26.620 393.600 26.760 ;
        RECT 62.170 26.560 62.490 26.620 ;
      LAYER via ;
        RECT 62.200 26.560 62.460 26.820 ;
        RECT 400.300 27.240 400.560 27.500 ;
      LAYER met2 ;
        RECT 401.750 1600.450 402.030 1604.000 ;
        RECT 400.360 1600.310 402.030 1600.450 ;
        RECT 400.360 27.530 400.500 1600.310 ;
        RECT 401.750 1600.000 402.030 1600.310 ;
        RECT 400.300 27.210 400.560 27.530 ;
        RECT 62.200 26.530 62.460 26.850 ;
        RECT 62.260 2.400 62.400 26.530 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 27.100 419.450 27.160 ;
        RECT 979.870 27.100 980.190 27.160 ;
        RECT 419.130 26.960 980.190 27.100 ;
        RECT 419.130 26.900 419.450 26.960 ;
        RECT 979.870 26.900 980.190 26.960 ;
      LAYER via ;
        RECT 419.160 26.900 419.420 27.160 ;
        RECT 979.900 26.900 980.160 27.160 ;
      LAYER met2 ;
        RECT 985.950 1600.450 986.230 1604.000 ;
        RECT 979.960 1600.310 986.230 1600.450 ;
        RECT 979.960 27.190 980.100 1600.310 ;
        RECT 985.950 1600.000 986.230 1600.310 ;
        RECT 419.160 26.870 419.420 27.190 ;
        RECT 979.900 26.870 980.160 27.190 ;
        RECT 419.220 2.400 419.360 26.870 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 26.760 436.930 26.820 ;
        RECT 1014.370 26.760 1014.690 26.820 ;
        RECT 436.610 26.620 1014.690 26.760 ;
        RECT 436.610 26.560 436.930 26.620 ;
        RECT 1014.370 26.560 1014.690 26.620 ;
      LAYER via ;
        RECT 436.640 26.560 436.900 26.820 ;
        RECT 1014.400 26.560 1014.660 26.820 ;
      LAYER met2 ;
        RECT 1014.930 1600.450 1015.210 1604.000 ;
        RECT 1014.460 1600.310 1015.210 1600.450 ;
        RECT 1014.460 26.850 1014.600 1600.310 ;
        RECT 1014.930 1600.000 1015.210 1600.310 ;
        RECT 436.640 26.530 436.900 26.850 ;
        RECT 1014.400 26.530 1014.660 26.850 ;
        RECT 436.700 2.400 436.840 26.530 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.370 1600.450 1044.650 1604.000 ;
        RECT 1042.060 1600.310 1044.650 1600.450 ;
        RECT 1042.060 26.365 1042.200 1600.310 ;
        RECT 1044.370 1600.000 1044.650 1600.310 ;
        RECT 454.570 25.995 454.850 26.365 ;
        RECT 1041.990 25.995 1042.270 26.365 ;
        RECT 454.640 2.400 454.780 25.995 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 454.570 26.040 454.850 26.320 ;
        RECT 1041.990 26.040 1042.270 26.320 ;
      LAYER met3 ;
        RECT 454.545 26.330 454.875 26.345 ;
        RECT 1041.965 26.330 1042.295 26.345 ;
        RECT 454.545 26.030 1042.295 26.330 ;
        RECT 454.545 26.015 454.875 26.030 ;
        RECT 1041.965 26.015 1042.295 26.030 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.350 1600.450 1073.630 1604.000 ;
        RECT 1069.660 1600.310 1073.630 1600.450 ;
        RECT 1069.660 25.685 1069.800 1600.310 ;
        RECT 1073.350 1600.000 1073.630 1600.310 ;
        RECT 472.510 25.315 472.790 25.685 ;
        RECT 1069.590 25.315 1069.870 25.685 ;
        RECT 472.580 2.400 472.720 25.315 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 472.510 25.360 472.790 25.640 ;
        RECT 1069.590 25.360 1069.870 25.640 ;
      LAYER met3 ;
        RECT 472.485 25.650 472.815 25.665 ;
        RECT 1069.565 25.650 1069.895 25.665 ;
        RECT 472.485 25.350 1069.895 25.650 ;
        RECT 472.485 25.335 472.815 25.350 ;
        RECT 1069.565 25.335 1069.895 25.350 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.390 27.780 525.710 27.840 ;
        RECT 545.170 27.780 545.490 27.840 ;
        RECT 525.390 27.640 545.490 27.780 ;
        RECT 525.390 27.580 525.710 27.640 ;
        RECT 545.170 27.580 545.490 27.640 ;
        RECT 545.170 26.420 545.490 26.480 ;
        RECT 1097.170 26.420 1097.490 26.480 ;
        RECT 545.170 26.280 1097.490 26.420 ;
        RECT 545.170 26.220 545.490 26.280 ;
        RECT 1097.170 26.220 1097.490 26.280 ;
        RECT 490.430 26.080 490.750 26.140 ;
        RECT 525.390 26.080 525.710 26.140 ;
        RECT 490.430 25.940 525.710 26.080 ;
        RECT 490.430 25.880 490.750 25.940 ;
        RECT 525.390 25.880 525.710 25.940 ;
      LAYER via ;
        RECT 525.420 27.580 525.680 27.840 ;
        RECT 545.200 27.580 545.460 27.840 ;
        RECT 545.200 26.220 545.460 26.480 ;
        RECT 1097.200 26.220 1097.460 26.480 ;
        RECT 490.460 25.880 490.720 26.140 ;
        RECT 525.420 25.880 525.680 26.140 ;
      LAYER met2 ;
        RECT 1102.790 1600.450 1103.070 1604.000 ;
        RECT 1097.260 1600.310 1103.070 1600.450 ;
        RECT 525.420 27.550 525.680 27.870 ;
        RECT 545.200 27.550 545.460 27.870 ;
        RECT 525.480 26.170 525.620 27.550 ;
        RECT 545.260 26.510 545.400 27.550 ;
        RECT 1097.260 26.510 1097.400 1600.310 ;
        RECT 1102.790 1600.000 1103.070 1600.310 ;
        RECT 545.200 26.190 545.460 26.510 ;
        RECT 1097.200 26.190 1097.460 26.510 ;
        RECT 490.460 25.850 490.720 26.170 ;
        RECT 525.420 25.850 525.680 26.170 ;
        RECT 490.520 2.400 490.660 25.850 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.770 1600.380 1132.050 1604.000 ;
        RECT 1131.760 1600.000 1132.050 1600.380 ;
        RECT 1131.760 25.005 1131.900 1600.000 ;
        RECT 507.930 24.635 508.210 25.005 ;
        RECT 1131.690 24.635 1131.970 25.005 ;
        RECT 508.000 2.400 508.140 24.635 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 507.930 24.680 508.210 24.960 ;
        RECT 1131.690 24.680 1131.970 24.960 ;
      LAYER met3 ;
        RECT 507.905 24.970 508.235 24.985 ;
        RECT 1131.665 24.970 1131.995 24.985 ;
        RECT 507.905 24.670 1131.995 24.970 ;
        RECT 507.905 24.655 508.235 24.670 ;
        RECT 1131.665 24.655 1131.995 24.670 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 525.850 26.080 526.170 26.140 ;
        RECT 1159.270 26.080 1159.590 26.140 ;
        RECT 525.850 25.940 1159.590 26.080 ;
        RECT 525.850 25.880 526.170 25.940 ;
        RECT 1159.270 25.880 1159.590 25.940 ;
      LAYER via ;
        RECT 525.880 25.880 526.140 26.140 ;
        RECT 1159.300 25.880 1159.560 26.140 ;
      LAYER met2 ;
        RECT 1161.210 1600.450 1161.490 1604.000 ;
        RECT 1159.360 1600.310 1161.490 1600.450 ;
        RECT 1159.360 26.170 1159.500 1600.310 ;
        RECT 1161.210 1600.000 1161.490 1600.310 ;
        RECT 525.880 25.850 526.140 26.170 ;
        RECT 1159.300 25.850 1159.560 26.170 ;
        RECT 525.940 2.400 526.080 25.850 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 543.790 31.860 544.110 31.920 ;
        RECT 1186.870 31.860 1187.190 31.920 ;
        RECT 543.790 31.720 1187.190 31.860 ;
        RECT 543.790 31.660 544.110 31.720 ;
        RECT 1186.870 31.660 1187.190 31.720 ;
      LAYER via ;
        RECT 543.820 31.660 544.080 31.920 ;
        RECT 1186.900 31.660 1187.160 31.920 ;
      LAYER met2 ;
        RECT 1190.190 1600.450 1190.470 1604.000 ;
        RECT 1186.960 1600.310 1190.470 1600.450 ;
        RECT 1186.960 31.950 1187.100 1600.310 ;
        RECT 1190.190 1600.000 1190.470 1600.310 ;
        RECT 543.820 31.630 544.080 31.950 ;
        RECT 1186.900 31.630 1187.160 31.950 ;
        RECT 543.880 2.400 544.020 31.630 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 561.730 31.520 562.050 31.580 ;
        RECT 1214.470 31.520 1214.790 31.580 ;
        RECT 561.730 31.380 1214.790 31.520 ;
        RECT 561.730 31.320 562.050 31.380 ;
        RECT 1214.470 31.320 1214.790 31.380 ;
      LAYER via ;
        RECT 561.760 31.320 562.020 31.580 ;
        RECT 1214.500 31.320 1214.760 31.580 ;
      LAYER met2 ;
        RECT 1219.170 1600.450 1219.450 1604.000 ;
        RECT 1214.560 1600.310 1219.450 1600.450 ;
        RECT 1214.560 31.610 1214.700 1600.310 ;
        RECT 1219.170 1600.000 1219.450 1600.310 ;
        RECT 561.760 31.290 562.020 31.610 ;
        RECT 1214.500 31.290 1214.760 31.610 ;
        RECT 561.820 2.400 561.960 31.290 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 31.180 579.990 31.240 ;
        RECT 1242.070 31.180 1242.390 31.240 ;
        RECT 579.670 31.040 1242.390 31.180 ;
        RECT 579.670 30.980 579.990 31.040 ;
        RECT 1242.070 30.980 1242.390 31.040 ;
      LAYER via ;
        RECT 579.700 30.980 579.960 31.240 ;
        RECT 1242.100 30.980 1242.360 31.240 ;
      LAYER met2 ;
        RECT 1248.610 1600.450 1248.890 1604.000 ;
        RECT 1242.160 1600.310 1248.890 1600.450 ;
        RECT 1242.160 31.270 1242.300 1600.310 ;
        RECT 1248.610 1600.000 1248.890 1600.310 ;
        RECT 579.700 30.950 579.960 31.270 ;
        RECT 1242.100 30.950 1242.360 31.270 ;
        RECT 579.760 2.400 579.900 30.950 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 252.150 1593.480 252.470 1593.540 ;
        RECT 440.750 1593.480 441.070 1593.540 ;
        RECT 252.150 1593.340 441.070 1593.480 ;
        RECT 252.150 1593.280 252.470 1593.340 ;
        RECT 440.750 1593.280 441.070 1593.340 ;
        RECT 86.090 15.540 86.410 15.600 ;
        RECT 252.150 15.540 252.470 15.600 ;
        RECT 86.090 15.400 187.980 15.540 ;
        RECT 86.090 15.340 86.410 15.400 ;
        RECT 187.840 14.860 187.980 15.400 ;
        RECT 239.820 15.400 252.470 15.540 ;
        RECT 239.820 14.860 239.960 15.400 ;
        RECT 252.150 15.340 252.470 15.400 ;
        RECT 187.840 14.720 239.960 14.860 ;
      LAYER via ;
        RECT 252.180 1593.280 252.440 1593.540 ;
        RECT 440.780 1593.280 441.040 1593.540 ;
        RECT 86.120 15.340 86.380 15.600 ;
        RECT 252.180 15.340 252.440 15.600 ;
      LAYER met2 ;
        RECT 440.850 1600.380 441.130 1604.000 ;
        RECT 440.840 1600.000 441.130 1600.380 ;
        RECT 440.840 1593.570 440.980 1600.000 ;
        RECT 252.180 1593.250 252.440 1593.570 ;
        RECT 440.780 1593.250 441.040 1593.570 ;
        RECT 252.240 15.630 252.380 1593.250 ;
        RECT 86.120 15.310 86.380 15.630 ;
        RECT 252.180 15.310 252.440 15.630 ;
        RECT 86.180 2.400 86.320 15.310 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 672.590 1592.120 672.910 1592.180 ;
        RECT 1277.490 1592.120 1277.810 1592.180 ;
        RECT 672.590 1591.980 1277.810 1592.120 ;
        RECT 672.590 1591.920 672.910 1591.980 ;
        RECT 1277.490 1591.920 1277.810 1591.980 ;
        RECT 597.150 25.060 597.470 25.120 ;
        RECT 672.590 25.060 672.910 25.120 ;
        RECT 597.150 24.920 672.910 25.060 ;
        RECT 597.150 24.860 597.470 24.920 ;
        RECT 672.590 24.860 672.910 24.920 ;
      LAYER via ;
        RECT 672.620 1591.920 672.880 1592.180 ;
        RECT 1277.520 1591.920 1277.780 1592.180 ;
        RECT 597.180 24.860 597.440 25.120 ;
        RECT 672.620 24.860 672.880 25.120 ;
      LAYER met2 ;
        RECT 1277.590 1600.380 1277.870 1604.000 ;
        RECT 1277.580 1600.000 1277.870 1600.380 ;
        RECT 1277.580 1592.210 1277.720 1600.000 ;
        RECT 672.620 1591.890 672.880 1592.210 ;
        RECT 1277.520 1591.890 1277.780 1592.210 ;
        RECT 672.680 25.150 672.820 1591.890 ;
        RECT 597.180 24.830 597.440 25.150 ;
        RECT 672.620 24.830 672.880 25.150 ;
        RECT 597.240 2.400 597.380 24.830 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 30.840 615.410 30.900 ;
        RECT 1304.170 30.840 1304.490 30.900 ;
        RECT 615.090 30.700 1304.490 30.840 ;
        RECT 615.090 30.640 615.410 30.700 ;
        RECT 1304.170 30.640 1304.490 30.700 ;
      LAYER via ;
        RECT 615.120 30.640 615.380 30.900 ;
        RECT 1304.200 30.640 1304.460 30.900 ;
      LAYER met2 ;
        RECT 1307.030 1600.450 1307.310 1604.000 ;
        RECT 1304.260 1600.310 1307.310 1600.450 ;
        RECT 1304.260 30.930 1304.400 1600.310 ;
        RECT 1307.030 1600.000 1307.310 1600.310 ;
        RECT 615.120 30.610 615.380 30.930 ;
        RECT 1304.200 30.610 1304.460 30.930 ;
        RECT 615.180 2.400 615.320 30.610 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 26.080 110.330 26.140 ;
        RECT 476.170 26.080 476.490 26.140 ;
        RECT 110.010 25.940 476.490 26.080 ;
        RECT 110.010 25.880 110.330 25.940 ;
        RECT 476.170 25.880 476.490 25.940 ;
      LAYER via ;
        RECT 110.040 25.880 110.300 26.140 ;
        RECT 476.200 25.880 476.460 26.140 ;
      LAYER met2 ;
        RECT 479.490 1600.450 479.770 1604.000 ;
        RECT 476.260 1600.310 479.770 1600.450 ;
        RECT 476.260 26.170 476.400 1600.310 ;
        RECT 479.490 1600.000 479.770 1600.310 ;
        RECT 110.040 25.850 110.300 26.170 ;
        RECT 476.200 25.850 476.460 26.170 ;
        RECT 110.100 13.330 110.240 25.850 ;
        RECT 109.640 13.190 110.240 13.330 ;
        RECT 109.640 2.400 109.780 13.190 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 25.740 133.790 25.800 ;
        RECT 409.470 25.740 409.790 25.800 ;
        RECT 133.470 25.600 409.790 25.740 ;
        RECT 133.470 25.540 133.790 25.600 ;
        RECT 409.470 25.540 409.790 25.600 ;
        RECT 410.390 25.740 410.710 25.800 ;
        RECT 517.570 25.740 517.890 25.800 ;
        RECT 410.390 25.600 517.890 25.740 ;
        RECT 410.390 25.540 410.710 25.600 ;
        RECT 517.570 25.540 517.890 25.600 ;
      LAYER via ;
        RECT 133.500 25.540 133.760 25.800 ;
        RECT 409.500 25.540 409.760 25.800 ;
        RECT 410.420 25.540 410.680 25.800 ;
        RECT 517.600 25.540 517.860 25.800 ;
      LAYER met2 ;
        RECT 518.590 1600.450 518.870 1604.000 ;
        RECT 517.660 1600.310 518.870 1600.450 ;
        RECT 409.560 26.110 410.620 26.250 ;
        RECT 409.560 25.830 409.700 26.110 ;
        RECT 410.480 25.830 410.620 26.110 ;
        RECT 517.660 25.830 517.800 1600.310 ;
        RECT 518.590 1600.000 518.870 1600.310 ;
        RECT 133.500 25.510 133.760 25.830 ;
        RECT 409.500 25.510 409.760 25.830 ;
        RECT 410.420 25.510 410.680 25.830 ;
        RECT 517.600 25.510 517.860 25.830 ;
        RECT 133.560 2.400 133.700 25.510 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 25.400 151.730 25.460 ;
        RECT 409.930 25.400 410.250 25.460 ;
        RECT 151.410 25.260 410.250 25.400 ;
        RECT 151.410 25.200 151.730 25.260 ;
        RECT 409.930 25.200 410.250 25.260 ;
        RECT 434.310 25.400 434.630 25.460 ;
        RECT 545.630 25.400 545.950 25.460 ;
        RECT 434.310 25.260 545.950 25.400 ;
        RECT 434.310 25.200 434.630 25.260 ;
        RECT 545.630 25.200 545.950 25.260 ;
      LAYER via ;
        RECT 151.440 25.200 151.700 25.460 ;
        RECT 409.960 25.200 410.220 25.460 ;
        RECT 434.340 25.200 434.600 25.460 ;
        RECT 545.660 25.200 545.920 25.460 ;
      LAYER met2 ;
        RECT 547.570 1600.450 547.850 1604.000 ;
        RECT 545.260 1600.310 547.850 1600.450 ;
        RECT 545.260 28.290 545.400 1600.310 ;
        RECT 547.570 1600.000 547.850 1600.310 ;
        RECT 545.260 28.150 545.860 28.290 ;
        RECT 151.440 25.170 151.700 25.490 ;
        RECT 409.950 25.315 410.230 25.685 ;
        RECT 434.330 25.315 434.610 25.685 ;
        RECT 545.720 25.490 545.860 28.150 ;
        RECT 409.960 25.170 410.220 25.315 ;
        RECT 434.340 25.170 434.600 25.315 ;
        RECT 545.660 25.170 545.920 25.490 ;
        RECT 151.500 2.400 151.640 25.170 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 409.950 25.360 410.230 25.640 ;
        RECT 434.330 25.360 434.610 25.640 ;
      LAYER met3 ;
        RECT 409.925 25.650 410.255 25.665 ;
        RECT 434.305 25.650 434.635 25.665 ;
        RECT 409.925 25.350 434.635 25.650 ;
        RECT 409.925 25.335 410.255 25.350 ;
        RECT 434.305 25.335 434.635 25.350 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 410.480 25.260 433.160 25.400 ;
        RECT 169.350 25.060 169.670 25.120 ;
        RECT 410.480 25.060 410.620 25.260 ;
        RECT 169.350 24.920 410.620 25.060 ;
        RECT 433.020 25.060 433.160 25.260 ;
        RECT 572.770 25.060 573.090 25.120 ;
        RECT 433.020 24.920 573.090 25.060 ;
        RECT 169.350 24.860 169.670 24.920 ;
        RECT 572.770 24.860 573.090 24.920 ;
      LAYER via ;
        RECT 169.380 24.860 169.640 25.120 ;
        RECT 572.800 24.860 573.060 25.120 ;
      LAYER met2 ;
        RECT 577.010 1600.450 577.290 1604.000 ;
        RECT 572.860 1600.310 577.290 1600.450 ;
        RECT 572.860 25.150 573.000 1600.310 ;
        RECT 577.010 1600.000 577.290 1600.310 ;
        RECT 169.380 24.830 169.640 25.150 ;
        RECT 572.800 24.830 573.060 25.150 ;
        RECT 169.440 2.400 169.580 24.830 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 186.830 24.720 187.150 24.780 ;
        RECT 409.930 24.720 410.250 24.780 ;
        RECT 186.830 24.580 410.250 24.720 ;
        RECT 186.830 24.520 187.150 24.580 ;
        RECT 409.930 24.520 410.250 24.580 ;
        RECT 433.850 24.720 434.170 24.780 ;
        RECT 600.370 24.720 600.690 24.780 ;
        RECT 433.850 24.580 600.690 24.720 ;
        RECT 433.850 24.520 434.170 24.580 ;
        RECT 600.370 24.520 600.690 24.580 ;
      LAYER via ;
        RECT 186.860 24.520 187.120 24.780 ;
        RECT 409.960 24.520 410.220 24.780 ;
        RECT 433.880 24.520 434.140 24.780 ;
        RECT 600.400 24.520 600.660 24.780 ;
      LAYER met2 ;
        RECT 605.990 1600.450 606.270 1604.000 ;
        RECT 600.460 1600.310 606.270 1600.450 ;
        RECT 186.860 24.490 187.120 24.810 ;
        RECT 409.950 24.635 410.230 25.005 ;
        RECT 433.870 24.635 434.150 25.005 ;
        RECT 600.460 24.810 600.600 1600.310 ;
        RECT 605.990 1600.000 606.270 1600.310 ;
        RECT 409.960 24.490 410.220 24.635 ;
        RECT 433.880 24.490 434.140 24.635 ;
        RECT 600.400 24.490 600.660 24.810 ;
        RECT 186.920 2.400 187.060 24.490 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 409.950 24.680 410.230 24.960 ;
        RECT 433.870 24.680 434.150 24.960 ;
      LAYER met3 ;
        RECT 409.925 24.970 410.255 24.985 ;
        RECT 433.845 24.970 434.175 24.985 ;
        RECT 409.925 24.670 434.175 24.970 ;
        RECT 409.925 24.655 410.255 24.670 ;
        RECT 433.845 24.655 434.175 24.670 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 204.770 24.380 205.090 24.440 ;
        RECT 394.290 24.380 394.610 24.440 ;
        RECT 204.770 24.240 394.610 24.380 ;
        RECT 204.770 24.180 205.090 24.240 ;
        RECT 394.290 24.180 394.610 24.240 ;
        RECT 434.310 24.380 434.630 24.440 ;
        RECT 634.870 24.380 635.190 24.440 ;
        RECT 434.310 24.240 635.190 24.380 ;
        RECT 434.310 24.180 434.630 24.240 ;
        RECT 634.870 24.180 635.190 24.240 ;
      LAYER via ;
        RECT 204.800 24.180 205.060 24.440 ;
        RECT 394.320 24.180 394.580 24.440 ;
        RECT 434.340 24.180 434.600 24.440 ;
        RECT 634.900 24.180 635.160 24.440 ;
      LAYER met2 ;
        RECT 635.430 1600.450 635.710 1604.000 ;
        RECT 634.960 1600.310 635.710 1600.450 ;
        RECT 634.960 24.470 635.100 1600.310 ;
        RECT 635.430 1600.000 635.710 1600.310 ;
        RECT 204.800 24.150 205.060 24.470 ;
        RECT 394.320 24.325 394.580 24.470 ;
        RECT 434.340 24.325 434.600 24.470 ;
        RECT 204.860 2.400 205.000 24.150 ;
        RECT 394.310 23.955 394.590 24.325 ;
        RECT 434.330 23.955 434.610 24.325 ;
        RECT 634.900 24.150 635.160 24.470 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 394.310 24.000 394.590 24.280 ;
        RECT 434.330 24.000 434.610 24.280 ;
      LAYER met3 ;
        RECT 394.285 24.290 394.615 24.305 ;
        RECT 434.305 24.290 434.635 24.305 ;
        RECT 394.285 23.990 434.635 24.290 ;
        RECT 394.285 23.975 394.615 23.990 ;
        RECT 434.305 23.975 434.635 23.990 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 222.710 24.040 223.030 24.100 ;
        RECT 662.470 24.040 662.790 24.100 ;
        RECT 222.710 23.900 662.790 24.040 ;
        RECT 222.710 23.840 223.030 23.900 ;
        RECT 662.470 23.840 662.790 23.900 ;
      LAYER via ;
        RECT 222.740 23.840 223.000 24.100 ;
        RECT 662.500 23.840 662.760 24.100 ;
      LAYER met2 ;
        RECT 664.410 1600.450 664.690 1604.000 ;
        RECT 662.560 1600.310 664.690 1600.450 ;
        RECT 662.560 24.130 662.700 1600.310 ;
        RECT 664.410 1600.000 664.690 1600.310 ;
        RECT 222.740 23.810 223.000 24.130 ;
        RECT 662.500 23.810 662.760 24.130 ;
        RECT 222.800 2.400 222.940 23.810 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 310.570 16.900 310.890 16.960 ;
        RECT 331.730 16.900 332.050 16.960 ;
        RECT 310.570 16.760 332.050 16.900 ;
        RECT 310.570 16.700 310.890 16.760 ;
        RECT 331.730 16.700 332.050 16.760 ;
        RECT 20.310 16.560 20.630 16.620 ;
        RECT 305.050 16.560 305.370 16.620 ;
        RECT 20.310 16.420 305.370 16.560 ;
        RECT 20.310 16.360 20.630 16.420 ;
        RECT 305.050 16.360 305.370 16.420 ;
      LAYER via ;
        RECT 310.600 16.700 310.860 16.960 ;
        RECT 331.760 16.700 332.020 16.960 ;
        RECT 20.340 16.360 20.600 16.620 ;
        RECT 305.080 16.360 305.340 16.620 ;
      LAYER met2 ;
        RECT 333.670 1600.450 333.950 1604.000 ;
        RECT 331.820 1600.310 333.950 1600.450 ;
        RECT 331.820 16.990 331.960 1600.310 ;
        RECT 333.670 1600.000 333.950 1600.310 ;
        RECT 310.600 16.845 310.860 16.990 ;
        RECT 20.340 16.330 20.600 16.650 ;
        RECT 305.070 16.475 305.350 16.845 ;
        RECT 310.590 16.475 310.870 16.845 ;
        RECT 331.760 16.670 332.020 16.990 ;
        RECT 305.080 16.330 305.340 16.475 ;
        RECT 20.400 2.400 20.540 16.330 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 305.070 16.520 305.350 16.800 ;
        RECT 310.590 16.520 310.870 16.800 ;
      LAYER met3 ;
        RECT 305.045 16.810 305.375 16.825 ;
        RECT 310.565 16.810 310.895 16.825 ;
        RECT 305.045 16.510 310.895 16.810 ;
        RECT 305.045 16.495 305.375 16.510 ;
        RECT 310.565 16.495 310.895 16.510 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 44.230 20.640 44.550 20.700 ;
        RECT 358.870 20.640 359.190 20.700 ;
        RECT 44.230 20.500 359.190 20.640 ;
        RECT 44.230 20.440 44.550 20.500 ;
        RECT 358.870 20.440 359.190 20.500 ;
        RECT 365.310 20.640 365.630 20.700 ;
        RECT 372.670 20.640 372.990 20.700 ;
        RECT 365.310 20.500 372.990 20.640 ;
        RECT 365.310 20.440 365.630 20.500 ;
        RECT 372.670 20.440 372.990 20.500 ;
      LAYER via ;
        RECT 44.260 20.440 44.520 20.700 ;
        RECT 358.900 20.440 359.160 20.700 ;
        RECT 365.340 20.440 365.600 20.700 ;
        RECT 372.700 20.440 372.960 20.700 ;
      LAYER met2 ;
        RECT 372.770 1600.380 373.050 1604.000 ;
        RECT 372.760 1600.000 373.050 1600.380 ;
        RECT 44.260 20.410 44.520 20.730 ;
        RECT 358.890 20.555 359.170 20.925 ;
        RECT 365.330 20.555 365.610 20.925 ;
        RECT 372.760 20.730 372.900 1600.000 ;
        RECT 358.900 20.410 359.160 20.555 ;
        RECT 365.340 20.410 365.600 20.555 ;
        RECT 372.700 20.410 372.960 20.730 ;
        RECT 44.320 2.400 44.460 20.410 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 358.890 20.600 359.170 20.880 ;
        RECT 365.330 20.600 365.610 20.880 ;
      LAYER met3 ;
        RECT 358.865 20.890 359.195 20.905 ;
        RECT 365.305 20.890 365.635 20.905 ;
        RECT 358.865 20.590 365.635 20.890 ;
        RECT 358.865 20.575 359.195 20.590 ;
        RECT 365.305 20.575 365.635 20.590 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 14.860 246.950 14.920 ;
        RECT 696.970 14.860 697.290 14.920 ;
        RECT 246.630 14.720 697.290 14.860 ;
        RECT 246.630 14.660 246.950 14.720 ;
        RECT 696.970 14.660 697.290 14.720 ;
      LAYER via ;
        RECT 246.660 14.660 246.920 14.920 ;
        RECT 697.000 14.660 697.260 14.920 ;
      LAYER met2 ;
        RECT 703.510 1600.450 703.790 1604.000 ;
        RECT 697.060 1600.310 703.790 1600.450 ;
        RECT 697.060 14.950 697.200 1600.310 ;
        RECT 703.510 1600.000 703.790 1600.310 ;
        RECT 246.660 14.630 246.920 14.950 ;
        RECT 697.000 14.630 697.260 14.950 ;
        RECT 246.720 2.400 246.860 14.630 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 624.290 1587.360 624.610 1587.420 ;
        RECT 732.850 1587.360 733.170 1587.420 ;
        RECT 624.290 1587.220 733.170 1587.360 ;
        RECT 624.290 1587.160 624.610 1587.220 ;
        RECT 732.850 1587.160 733.170 1587.220 ;
        RECT 469.270 27.780 469.590 27.840 ;
        RECT 518.030 27.780 518.350 27.840 ;
        RECT 469.270 27.640 518.350 27.780 ;
        RECT 469.270 27.580 469.590 27.640 ;
        RECT 518.030 27.580 518.350 27.640 ;
        RECT 303.670 27.100 303.990 27.160 ;
        RECT 392.910 27.100 393.230 27.160 ;
        RECT 303.670 26.960 393.230 27.100 ;
        RECT 303.670 26.900 303.990 26.960 ;
        RECT 392.910 26.900 393.230 26.960 ;
        RECT 264.110 26.420 264.430 26.480 ;
        RECT 303.670 26.420 303.990 26.480 ;
        RECT 264.110 26.280 303.990 26.420 ;
        RECT 264.110 26.220 264.430 26.280 ;
        RECT 303.670 26.220 303.990 26.280 ;
        RECT 392.910 26.420 393.230 26.480 ;
        RECT 469.270 26.420 469.590 26.480 ;
        RECT 392.910 26.280 469.590 26.420 ;
        RECT 392.910 26.220 393.230 26.280 ;
        RECT 469.270 26.220 469.590 26.280 ;
        RECT 518.030 25.740 518.350 25.800 ;
        RECT 518.030 25.600 546.320 25.740 ;
        RECT 518.030 25.540 518.350 25.600 ;
        RECT 546.180 25.400 546.320 25.600 ;
        RECT 624.290 25.400 624.610 25.460 ;
        RECT 546.180 25.260 624.610 25.400 ;
        RECT 624.290 25.200 624.610 25.260 ;
      LAYER via ;
        RECT 624.320 1587.160 624.580 1587.420 ;
        RECT 732.880 1587.160 733.140 1587.420 ;
        RECT 469.300 27.580 469.560 27.840 ;
        RECT 518.060 27.580 518.320 27.840 ;
        RECT 303.700 26.900 303.960 27.160 ;
        RECT 392.940 26.900 393.200 27.160 ;
        RECT 264.140 26.220 264.400 26.480 ;
        RECT 303.700 26.220 303.960 26.480 ;
        RECT 392.940 26.220 393.200 26.480 ;
        RECT 469.300 26.220 469.560 26.480 ;
        RECT 518.060 25.540 518.320 25.800 ;
        RECT 624.320 25.200 624.580 25.460 ;
      LAYER met2 ;
        RECT 732.950 1600.380 733.230 1604.000 ;
        RECT 732.940 1600.000 733.230 1600.380 ;
        RECT 732.940 1587.450 733.080 1600.000 ;
        RECT 624.320 1587.130 624.580 1587.450 ;
        RECT 732.880 1587.130 733.140 1587.450 ;
        RECT 469.300 27.550 469.560 27.870 ;
        RECT 518.060 27.550 518.320 27.870 ;
        RECT 303.700 26.870 303.960 27.190 ;
        RECT 392.940 26.870 393.200 27.190 ;
        RECT 303.760 26.510 303.900 26.870 ;
        RECT 393.000 26.510 393.140 26.870 ;
        RECT 469.360 26.510 469.500 27.550 ;
        RECT 264.140 26.190 264.400 26.510 ;
        RECT 303.700 26.190 303.960 26.510 ;
        RECT 392.940 26.190 393.200 26.510 ;
        RECT 469.300 26.190 469.560 26.510 ;
        RECT 264.200 2.400 264.340 26.190 ;
        RECT 518.120 25.830 518.260 27.550 ;
        RECT 518.060 25.510 518.320 25.830 ;
        RECT 624.380 25.490 624.520 1587.130 ;
        RECT 624.320 25.170 624.580 25.490 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 15.880 282.370 15.940 ;
        RECT 759.070 15.880 759.390 15.940 ;
        RECT 282.050 15.740 759.390 15.880 ;
        RECT 282.050 15.680 282.370 15.740 ;
        RECT 759.070 15.680 759.390 15.740 ;
      LAYER via ;
        RECT 282.080 15.680 282.340 15.940 ;
        RECT 759.100 15.680 759.360 15.940 ;
      LAYER met2 ;
        RECT 761.930 1600.450 762.210 1604.000 ;
        RECT 759.160 1600.310 762.210 1600.450 ;
        RECT 759.160 15.970 759.300 1600.310 ;
        RECT 761.930 1600.000 762.210 1600.310 ;
        RECT 282.080 15.650 282.340 15.970 ;
        RECT 759.100 15.650 759.360 15.970 ;
        RECT 282.140 2.400 282.280 15.650 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 299.990 32.200 300.310 32.260 ;
        RECT 786.670 32.200 786.990 32.260 ;
        RECT 299.990 32.060 786.990 32.200 ;
        RECT 299.990 32.000 300.310 32.060 ;
        RECT 786.670 32.000 786.990 32.060 ;
      LAYER via ;
        RECT 300.020 32.000 300.280 32.260 ;
        RECT 786.700 32.000 786.960 32.260 ;
      LAYER met2 ;
        RECT 790.910 1600.450 791.190 1604.000 ;
        RECT 786.760 1600.310 791.190 1600.450 ;
        RECT 786.760 32.290 786.900 1600.310 ;
        RECT 790.910 1600.000 791.190 1600.310 ;
        RECT 300.020 31.970 300.280 32.290 ;
        RECT 786.700 31.970 786.960 32.290 ;
        RECT 300.080 2.400 300.220 31.970 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.930 16.220 318.250 16.280 ;
        RECT 814.270 16.220 814.590 16.280 ;
        RECT 317.930 16.080 814.590 16.220 ;
        RECT 317.930 16.020 318.250 16.080 ;
        RECT 814.270 16.020 814.590 16.080 ;
      LAYER via ;
        RECT 317.960 16.020 318.220 16.280 ;
        RECT 814.300 16.020 814.560 16.280 ;
      LAYER met2 ;
        RECT 820.350 1600.450 820.630 1604.000 ;
        RECT 814.360 1600.310 820.630 1600.450 ;
        RECT 814.360 16.310 814.500 1600.310 ;
        RECT 820.350 1600.000 820.630 1600.310 ;
        RECT 317.960 15.990 318.220 16.310 ;
        RECT 814.300 15.990 814.560 16.310 ;
        RECT 318.020 2.400 318.160 15.990 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 337.710 1589.060 338.030 1589.120 ;
        RECT 849.230 1589.060 849.550 1589.120 ;
        RECT 337.710 1588.920 849.550 1589.060 ;
        RECT 337.710 1588.860 338.030 1588.920 ;
        RECT 849.230 1588.860 849.550 1588.920 ;
        RECT 335.410 23.700 335.730 23.760 ;
        RECT 337.710 23.700 338.030 23.760 ;
        RECT 335.410 23.560 338.030 23.700 ;
        RECT 335.410 23.500 335.730 23.560 ;
        RECT 337.710 23.500 338.030 23.560 ;
        RECT 335.410 2.960 335.730 3.020 ;
        RECT 335.870 2.960 336.190 3.020 ;
        RECT 335.410 2.820 336.190 2.960 ;
        RECT 335.410 2.760 335.730 2.820 ;
        RECT 335.870 2.760 336.190 2.820 ;
      LAYER via ;
        RECT 337.740 1588.860 338.000 1589.120 ;
        RECT 849.260 1588.860 849.520 1589.120 ;
        RECT 335.440 23.500 335.700 23.760 ;
        RECT 337.740 23.500 338.000 23.760 ;
        RECT 335.440 2.760 335.700 3.020 ;
        RECT 335.900 2.760 336.160 3.020 ;
      LAYER met2 ;
        RECT 849.330 1600.380 849.610 1604.000 ;
        RECT 849.320 1600.000 849.610 1600.380 ;
        RECT 849.320 1589.150 849.460 1600.000 ;
        RECT 337.740 1588.830 338.000 1589.150 ;
        RECT 849.260 1588.830 849.520 1589.150 ;
        RECT 337.800 23.790 337.940 1588.830 ;
        RECT 335.440 23.470 335.700 23.790 ;
        RECT 337.740 23.470 338.000 23.790 ;
        RECT 335.500 3.050 335.640 23.470 ;
        RECT 335.440 2.730 335.700 3.050 ;
        RECT 335.900 2.730 336.160 3.050 ;
        RECT 335.960 2.400 336.100 2.730 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 376.350 16.900 376.670 16.960 ;
        RECT 876.370 16.900 876.690 16.960 ;
        RECT 376.350 16.760 876.690 16.900 ;
        RECT 376.350 16.700 376.670 16.760 ;
        RECT 876.370 16.700 876.690 16.760 ;
        RECT 353.350 16.560 353.670 16.620 ;
        RECT 375.430 16.560 375.750 16.620 ;
        RECT 353.350 16.420 375.750 16.560 ;
        RECT 353.350 16.360 353.670 16.420 ;
        RECT 375.430 16.360 375.750 16.420 ;
      LAYER via ;
        RECT 376.380 16.700 376.640 16.960 ;
        RECT 876.400 16.700 876.660 16.960 ;
        RECT 353.380 16.360 353.640 16.620 ;
        RECT 375.460 16.360 375.720 16.620 ;
      LAYER met2 ;
        RECT 878.770 1600.450 879.050 1604.000 ;
        RECT 876.460 1600.310 879.050 1600.450 ;
        RECT 876.460 16.990 876.600 1600.310 ;
        RECT 878.770 1600.000 879.050 1600.310 ;
        RECT 376.380 16.730 376.640 16.990 ;
        RECT 375.520 16.670 376.640 16.730 ;
        RECT 876.400 16.670 876.660 16.990 ;
        RECT 375.520 16.650 376.580 16.670 ;
        RECT 353.380 16.330 353.640 16.650 ;
        RECT 375.460 16.590 376.580 16.650 ;
        RECT 375.460 16.330 375.720 16.590 ;
        RECT 353.440 2.400 353.580 16.330 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1589.740 372.530 1589.800 ;
        RECT 907.650 1589.740 907.970 1589.800 ;
        RECT 372.210 1589.600 907.970 1589.740 ;
        RECT 372.210 1589.540 372.530 1589.600 ;
        RECT 907.650 1589.540 907.970 1589.600 ;
        RECT 372.210 1498.080 372.530 1498.340 ;
        RECT 372.300 1497.660 372.440 1498.080 ;
        RECT 372.210 1497.400 372.530 1497.660 ;
        RECT 371.290 1490.460 371.610 1490.520 ;
        RECT 372.210 1490.460 372.530 1490.520 ;
        RECT 371.290 1490.320 372.530 1490.460 ;
        RECT 371.290 1490.260 371.610 1490.320 ;
        RECT 372.210 1490.260 372.530 1490.320 ;
        RECT 371.290 1442.180 371.610 1442.240 ;
        RECT 371.750 1442.180 372.070 1442.240 ;
        RECT 371.290 1442.040 372.070 1442.180 ;
        RECT 371.290 1441.980 371.610 1442.040 ;
        RECT 371.750 1441.980 372.070 1442.040 ;
        RECT 371.290 1345.620 371.610 1345.680 ;
        RECT 371.750 1345.620 372.070 1345.680 ;
        RECT 371.290 1345.480 372.070 1345.620 ;
        RECT 371.290 1345.420 371.610 1345.480 ;
        RECT 371.750 1345.420 372.070 1345.480 ;
        RECT 371.290 1249.060 371.610 1249.120 ;
        RECT 372.210 1249.060 372.530 1249.120 ;
        RECT 371.290 1248.920 372.530 1249.060 ;
        RECT 371.290 1248.860 371.610 1248.920 ;
        RECT 372.210 1248.860 372.530 1248.920 ;
        RECT 371.750 1207.580 372.070 1207.640 ;
        RECT 372.210 1207.580 372.530 1207.640 ;
        RECT 371.750 1207.440 372.530 1207.580 ;
        RECT 371.750 1207.380 372.070 1207.440 ;
        RECT 372.210 1207.380 372.530 1207.440 ;
        RECT 371.290 1152.500 371.610 1152.560 ;
        RECT 372.210 1152.500 372.530 1152.560 ;
        RECT 371.290 1152.360 372.530 1152.500 ;
        RECT 371.290 1152.300 371.610 1152.360 ;
        RECT 372.210 1152.300 372.530 1152.360 ;
        RECT 371.290 1007.320 371.610 1007.380 ;
        RECT 372.210 1007.320 372.530 1007.380 ;
        RECT 371.290 1007.180 372.530 1007.320 ;
        RECT 371.290 1007.120 371.610 1007.180 ;
        RECT 372.210 1007.120 372.530 1007.180 ;
        RECT 371.290 959.380 371.610 959.440 ;
        RECT 371.750 959.380 372.070 959.440 ;
        RECT 371.290 959.240 372.070 959.380 ;
        RECT 371.290 959.180 371.610 959.240 ;
        RECT 371.750 959.180 372.070 959.240 ;
        RECT 371.750 917.900 372.070 917.960 ;
        RECT 372.210 917.900 372.530 917.960 ;
        RECT 371.750 917.760 372.530 917.900 ;
        RECT 371.750 917.700 372.070 917.760 ;
        RECT 372.210 917.700 372.530 917.760 ;
        RECT 371.290 910.760 371.610 910.820 ;
        RECT 372.210 910.760 372.530 910.820 ;
        RECT 371.290 910.620 372.530 910.760 ;
        RECT 371.290 910.560 371.610 910.620 ;
        RECT 372.210 910.560 372.530 910.620 ;
        RECT 371.290 814.200 371.610 814.260 ;
        RECT 372.210 814.200 372.530 814.260 ;
        RECT 371.290 814.060 372.530 814.200 ;
        RECT 371.290 814.000 371.610 814.060 ;
        RECT 372.210 814.000 372.530 814.060 ;
        RECT 372.210 717.640 372.530 717.700 ;
        RECT 373.130 717.640 373.450 717.700 ;
        RECT 372.210 717.500 373.450 717.640 ;
        RECT 372.210 717.440 372.530 717.500 ;
        RECT 373.130 717.440 373.450 717.500 ;
        RECT 371.750 572.800 372.070 572.860 ;
        RECT 373.590 572.800 373.910 572.860 ;
        RECT 371.750 572.660 373.910 572.800 ;
        RECT 371.750 572.600 372.070 572.660 ;
        RECT 373.590 572.600 373.910 572.660 ;
        RECT 371.750 532.000 372.070 532.060 ;
        RECT 372.210 532.000 372.530 532.060 ;
        RECT 371.750 531.860 372.530 532.000 ;
        RECT 371.750 531.800 372.070 531.860 ;
        RECT 372.210 531.800 372.530 531.860 ;
        RECT 371.290 524.180 371.610 524.240 ;
        RECT 372.210 524.180 372.530 524.240 ;
        RECT 371.290 524.040 372.530 524.180 ;
        RECT 371.290 523.980 371.610 524.040 ;
        RECT 372.210 523.980 372.530 524.040 ;
        RECT 371.290 476.240 371.610 476.300 ;
        RECT 371.750 476.240 372.070 476.300 ;
        RECT 371.290 476.100 372.070 476.240 ;
        RECT 371.290 476.040 371.610 476.100 ;
        RECT 371.750 476.040 372.070 476.100 ;
        RECT 371.750 435.440 372.070 435.500 ;
        RECT 372.210 435.440 372.530 435.500 ;
        RECT 371.750 435.300 372.530 435.440 ;
        RECT 371.750 435.240 372.070 435.300 ;
        RECT 372.210 435.240 372.530 435.300 ;
        RECT 371.290 427.620 371.610 427.680 ;
        RECT 372.210 427.620 372.530 427.680 ;
        RECT 371.290 427.480 372.530 427.620 ;
        RECT 371.290 427.420 371.610 427.480 ;
        RECT 372.210 427.420 372.530 427.480 ;
        RECT 371.290 379.680 371.610 379.740 ;
        RECT 371.750 379.680 372.070 379.740 ;
        RECT 371.290 379.540 372.070 379.680 ;
        RECT 371.290 379.480 371.610 379.540 ;
        RECT 371.750 379.480 372.070 379.540 ;
        RECT 371.750 338.540 372.070 338.600 ;
        RECT 372.210 338.540 372.530 338.600 ;
        RECT 371.750 338.400 372.530 338.540 ;
        RECT 371.750 338.340 372.070 338.400 ;
        RECT 372.210 338.340 372.530 338.400 ;
        RECT 371.290 331.060 371.610 331.120 ;
        RECT 372.210 331.060 372.530 331.120 ;
        RECT 371.290 330.920 372.530 331.060 ;
        RECT 371.290 330.860 371.610 330.920 ;
        RECT 372.210 330.860 372.530 330.920 ;
        RECT 371.290 283.120 371.610 283.180 ;
        RECT 372.210 283.120 372.530 283.180 ;
        RECT 371.290 282.980 372.530 283.120 ;
        RECT 371.290 282.920 371.610 282.980 ;
        RECT 372.210 282.920 372.530 282.980 ;
        RECT 371.290 234.500 371.610 234.560 ;
        RECT 372.210 234.500 372.530 234.560 ;
        RECT 371.290 234.360 372.530 234.500 ;
        RECT 371.290 234.300 371.610 234.360 ;
        RECT 372.210 234.300 372.530 234.360 ;
        RECT 371.290 186.560 371.610 186.620 ;
        RECT 371.750 186.560 372.070 186.620 ;
        RECT 371.290 186.420 372.070 186.560 ;
        RECT 371.290 186.360 371.610 186.420 ;
        RECT 371.750 186.360 372.070 186.420 ;
        RECT 371.290 137.940 371.610 138.000 ;
        RECT 372.210 137.940 372.530 138.000 ;
        RECT 371.290 137.800 372.530 137.940 ;
        RECT 371.290 137.740 371.610 137.800 ;
        RECT 372.210 137.740 372.530 137.800 ;
        RECT 370.370 90.000 370.690 90.060 ;
        RECT 371.290 90.000 371.610 90.060 ;
        RECT 370.370 89.860 371.610 90.000 ;
        RECT 370.370 89.800 370.690 89.860 ;
        RECT 371.290 89.800 371.610 89.860 ;
        RECT 370.370 48.520 370.690 48.580 ;
        RECT 371.290 48.520 371.610 48.580 ;
        RECT 370.370 48.380 371.610 48.520 ;
        RECT 370.370 48.320 370.690 48.380 ;
        RECT 371.290 48.320 371.610 48.380 ;
      LAYER via ;
        RECT 372.240 1589.540 372.500 1589.800 ;
        RECT 907.680 1589.540 907.940 1589.800 ;
        RECT 372.240 1498.080 372.500 1498.340 ;
        RECT 372.240 1497.400 372.500 1497.660 ;
        RECT 371.320 1490.260 371.580 1490.520 ;
        RECT 372.240 1490.260 372.500 1490.520 ;
        RECT 371.320 1441.980 371.580 1442.240 ;
        RECT 371.780 1441.980 372.040 1442.240 ;
        RECT 371.320 1345.420 371.580 1345.680 ;
        RECT 371.780 1345.420 372.040 1345.680 ;
        RECT 371.320 1248.860 371.580 1249.120 ;
        RECT 372.240 1248.860 372.500 1249.120 ;
        RECT 371.780 1207.380 372.040 1207.640 ;
        RECT 372.240 1207.380 372.500 1207.640 ;
        RECT 371.320 1152.300 371.580 1152.560 ;
        RECT 372.240 1152.300 372.500 1152.560 ;
        RECT 371.320 1007.120 371.580 1007.380 ;
        RECT 372.240 1007.120 372.500 1007.380 ;
        RECT 371.320 959.180 371.580 959.440 ;
        RECT 371.780 959.180 372.040 959.440 ;
        RECT 371.780 917.700 372.040 917.960 ;
        RECT 372.240 917.700 372.500 917.960 ;
        RECT 371.320 910.560 371.580 910.820 ;
        RECT 372.240 910.560 372.500 910.820 ;
        RECT 371.320 814.000 371.580 814.260 ;
        RECT 372.240 814.000 372.500 814.260 ;
        RECT 372.240 717.440 372.500 717.700 ;
        RECT 373.160 717.440 373.420 717.700 ;
        RECT 371.780 572.600 372.040 572.860 ;
        RECT 373.620 572.600 373.880 572.860 ;
        RECT 371.780 531.800 372.040 532.060 ;
        RECT 372.240 531.800 372.500 532.060 ;
        RECT 371.320 523.980 371.580 524.240 ;
        RECT 372.240 523.980 372.500 524.240 ;
        RECT 371.320 476.040 371.580 476.300 ;
        RECT 371.780 476.040 372.040 476.300 ;
        RECT 371.780 435.240 372.040 435.500 ;
        RECT 372.240 435.240 372.500 435.500 ;
        RECT 371.320 427.420 371.580 427.680 ;
        RECT 372.240 427.420 372.500 427.680 ;
        RECT 371.320 379.480 371.580 379.740 ;
        RECT 371.780 379.480 372.040 379.740 ;
        RECT 371.780 338.340 372.040 338.600 ;
        RECT 372.240 338.340 372.500 338.600 ;
        RECT 371.320 330.860 371.580 331.120 ;
        RECT 372.240 330.860 372.500 331.120 ;
        RECT 371.320 282.920 371.580 283.180 ;
        RECT 372.240 282.920 372.500 283.180 ;
        RECT 371.320 234.300 371.580 234.560 ;
        RECT 372.240 234.300 372.500 234.560 ;
        RECT 371.320 186.360 371.580 186.620 ;
        RECT 371.780 186.360 372.040 186.620 ;
        RECT 371.320 137.740 371.580 138.000 ;
        RECT 372.240 137.740 372.500 138.000 ;
        RECT 370.400 89.800 370.660 90.060 ;
        RECT 371.320 89.800 371.580 90.060 ;
        RECT 370.400 48.320 370.660 48.580 ;
        RECT 371.320 48.320 371.580 48.580 ;
      LAYER met2 ;
        RECT 907.750 1600.380 908.030 1604.000 ;
        RECT 907.740 1600.000 908.030 1600.380 ;
        RECT 907.740 1589.830 907.880 1600.000 ;
        RECT 372.240 1589.510 372.500 1589.830 ;
        RECT 907.680 1589.510 907.940 1589.830 ;
        RECT 372.300 1498.370 372.440 1589.510 ;
        RECT 372.240 1498.050 372.500 1498.370 ;
        RECT 372.240 1497.370 372.500 1497.690 ;
        RECT 372.300 1490.550 372.440 1497.370 ;
        RECT 371.320 1490.230 371.580 1490.550 ;
        RECT 372.240 1490.230 372.500 1490.550 ;
        RECT 371.380 1442.270 371.520 1490.230 ;
        RECT 371.320 1441.950 371.580 1442.270 ;
        RECT 371.780 1441.950 372.040 1442.270 ;
        RECT 371.840 1401.210 371.980 1441.950 ;
        RECT 371.840 1401.070 372.440 1401.210 ;
        RECT 372.300 1393.845 372.440 1401.070 ;
        RECT 371.310 1393.475 371.590 1393.845 ;
        RECT 372.230 1393.475 372.510 1393.845 ;
        RECT 371.380 1345.710 371.520 1393.475 ;
        RECT 371.320 1345.390 371.580 1345.710 ;
        RECT 371.780 1345.390 372.040 1345.710 ;
        RECT 371.840 1304.650 371.980 1345.390 ;
        RECT 371.840 1304.510 372.440 1304.650 ;
        RECT 372.300 1297.285 372.440 1304.510 ;
        RECT 371.310 1296.915 371.590 1297.285 ;
        RECT 372.230 1296.915 372.510 1297.285 ;
        RECT 371.380 1249.150 371.520 1296.915 ;
        RECT 371.320 1248.830 371.580 1249.150 ;
        RECT 372.240 1248.830 372.500 1249.150 ;
        RECT 372.300 1208.770 372.440 1248.830 ;
        RECT 371.840 1208.630 372.440 1208.770 ;
        RECT 371.840 1207.670 371.980 1208.630 ;
        RECT 371.780 1207.350 372.040 1207.670 ;
        RECT 372.240 1207.350 372.500 1207.670 ;
        RECT 372.300 1200.725 372.440 1207.350 ;
        RECT 371.310 1200.355 371.590 1200.725 ;
        RECT 372.230 1200.355 372.510 1200.725 ;
        RECT 371.380 1152.590 371.520 1200.355 ;
        RECT 371.320 1152.270 371.580 1152.590 ;
        RECT 372.240 1152.270 372.500 1152.590 ;
        RECT 372.300 1104.165 372.440 1152.270 ;
        RECT 371.310 1103.795 371.590 1104.165 ;
        RECT 372.230 1103.795 372.510 1104.165 ;
        RECT 371.380 1055.885 371.520 1103.795 ;
        RECT 371.310 1055.515 371.590 1055.885 ;
        RECT 372.230 1055.515 372.510 1055.885 ;
        RECT 372.300 1007.410 372.440 1055.515 ;
        RECT 371.320 1007.090 371.580 1007.410 ;
        RECT 372.240 1007.090 372.500 1007.410 ;
        RECT 371.380 959.470 371.520 1007.090 ;
        RECT 371.320 959.150 371.580 959.470 ;
        RECT 371.780 959.150 372.040 959.470 ;
        RECT 371.840 917.990 371.980 959.150 ;
        RECT 371.780 917.670 372.040 917.990 ;
        RECT 372.240 917.670 372.500 917.990 ;
        RECT 372.300 910.850 372.440 917.670 ;
        RECT 371.320 910.530 371.580 910.850 ;
        RECT 372.240 910.530 372.500 910.850 ;
        RECT 371.380 862.765 371.520 910.530 ;
        RECT 371.310 862.395 371.590 862.765 ;
        RECT 372.230 862.395 372.510 862.765 ;
        RECT 372.300 814.290 372.440 862.395 ;
        RECT 371.320 813.970 371.580 814.290 ;
        RECT 372.240 813.970 372.500 814.290 ;
        RECT 371.380 766.205 371.520 813.970 ;
        RECT 371.310 765.835 371.590 766.205 ;
        RECT 372.230 765.835 372.510 766.205 ;
        RECT 372.300 717.730 372.440 765.835 ;
        RECT 372.240 717.410 372.500 717.730 ;
        RECT 373.160 717.410 373.420 717.730 ;
        RECT 373.220 628.165 373.360 717.410 ;
        RECT 372.230 627.795 372.510 628.165 ;
        RECT 373.150 627.795 373.430 628.165 ;
        RECT 372.300 620.685 372.440 627.795 ;
        RECT 372.230 620.315 372.510 620.685 ;
        RECT 373.610 620.315 373.890 620.685 ;
        RECT 373.680 572.890 373.820 620.315 ;
        RECT 371.780 572.570 372.040 572.890 ;
        RECT 373.620 572.570 373.880 572.890 ;
        RECT 371.840 532.090 371.980 572.570 ;
        RECT 371.780 531.770 372.040 532.090 ;
        RECT 372.240 531.770 372.500 532.090 ;
        RECT 372.300 524.270 372.440 531.770 ;
        RECT 371.320 523.950 371.580 524.270 ;
        RECT 372.240 523.950 372.500 524.270 ;
        RECT 371.380 476.330 371.520 523.950 ;
        RECT 371.320 476.010 371.580 476.330 ;
        RECT 371.780 476.010 372.040 476.330 ;
        RECT 371.840 435.530 371.980 476.010 ;
        RECT 371.780 435.210 372.040 435.530 ;
        RECT 372.240 435.210 372.500 435.530 ;
        RECT 372.300 427.710 372.440 435.210 ;
        RECT 371.320 427.390 371.580 427.710 ;
        RECT 372.240 427.390 372.500 427.710 ;
        RECT 371.380 379.770 371.520 427.390 ;
        RECT 371.320 379.450 371.580 379.770 ;
        RECT 371.780 379.450 372.040 379.770 ;
        RECT 371.840 338.630 371.980 379.450 ;
        RECT 371.780 338.310 372.040 338.630 ;
        RECT 372.240 338.310 372.500 338.630 ;
        RECT 372.300 331.150 372.440 338.310 ;
        RECT 371.320 330.830 371.580 331.150 ;
        RECT 372.240 330.830 372.500 331.150 ;
        RECT 371.380 283.210 371.520 330.830 ;
        RECT 371.320 282.890 371.580 283.210 ;
        RECT 372.240 282.890 372.500 283.210 ;
        RECT 372.300 242.490 372.440 282.890 ;
        RECT 371.840 242.350 372.440 242.490 ;
        RECT 371.840 241.810 371.980 242.350 ;
        RECT 371.840 241.670 372.440 241.810 ;
        RECT 372.300 234.590 372.440 241.670 ;
        RECT 371.320 234.270 371.580 234.590 ;
        RECT 372.240 234.270 372.500 234.590 ;
        RECT 371.380 186.650 371.520 234.270 ;
        RECT 371.320 186.330 371.580 186.650 ;
        RECT 371.780 186.330 372.040 186.650 ;
        RECT 371.840 145.250 371.980 186.330 ;
        RECT 371.840 145.110 372.440 145.250 ;
        RECT 372.300 138.030 372.440 145.110 ;
        RECT 371.320 137.710 371.580 138.030 ;
        RECT 372.240 137.710 372.500 138.030 ;
        RECT 371.380 90.090 371.520 137.710 ;
        RECT 370.400 89.770 370.660 90.090 ;
        RECT 371.320 89.770 371.580 90.090 ;
        RECT 370.460 48.610 370.600 89.770 ;
        RECT 370.400 48.290 370.660 48.610 ;
        RECT 371.320 48.290 371.580 48.610 ;
        RECT 371.380 2.400 371.520 48.290 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 371.310 1393.520 371.590 1393.800 ;
        RECT 372.230 1393.520 372.510 1393.800 ;
        RECT 371.310 1296.960 371.590 1297.240 ;
        RECT 372.230 1296.960 372.510 1297.240 ;
        RECT 371.310 1200.400 371.590 1200.680 ;
        RECT 372.230 1200.400 372.510 1200.680 ;
        RECT 371.310 1103.840 371.590 1104.120 ;
        RECT 372.230 1103.840 372.510 1104.120 ;
        RECT 371.310 1055.560 371.590 1055.840 ;
        RECT 372.230 1055.560 372.510 1055.840 ;
        RECT 371.310 862.440 371.590 862.720 ;
        RECT 372.230 862.440 372.510 862.720 ;
        RECT 371.310 765.880 371.590 766.160 ;
        RECT 372.230 765.880 372.510 766.160 ;
        RECT 372.230 627.840 372.510 628.120 ;
        RECT 373.150 627.840 373.430 628.120 ;
        RECT 372.230 620.360 372.510 620.640 ;
        RECT 373.610 620.360 373.890 620.640 ;
      LAYER met3 ;
        RECT 371.285 1393.810 371.615 1393.825 ;
        RECT 372.205 1393.810 372.535 1393.825 ;
        RECT 371.285 1393.510 372.535 1393.810 ;
        RECT 371.285 1393.495 371.615 1393.510 ;
        RECT 372.205 1393.495 372.535 1393.510 ;
        RECT 371.285 1297.250 371.615 1297.265 ;
        RECT 372.205 1297.250 372.535 1297.265 ;
        RECT 371.285 1296.950 372.535 1297.250 ;
        RECT 371.285 1296.935 371.615 1296.950 ;
        RECT 372.205 1296.935 372.535 1296.950 ;
        RECT 371.285 1200.690 371.615 1200.705 ;
        RECT 372.205 1200.690 372.535 1200.705 ;
        RECT 371.285 1200.390 372.535 1200.690 ;
        RECT 371.285 1200.375 371.615 1200.390 ;
        RECT 372.205 1200.375 372.535 1200.390 ;
        RECT 371.285 1104.130 371.615 1104.145 ;
        RECT 372.205 1104.130 372.535 1104.145 ;
        RECT 371.285 1103.830 372.535 1104.130 ;
        RECT 371.285 1103.815 371.615 1103.830 ;
        RECT 372.205 1103.815 372.535 1103.830 ;
        RECT 371.285 1055.850 371.615 1055.865 ;
        RECT 372.205 1055.850 372.535 1055.865 ;
        RECT 371.285 1055.550 372.535 1055.850 ;
        RECT 371.285 1055.535 371.615 1055.550 ;
        RECT 372.205 1055.535 372.535 1055.550 ;
        RECT 371.285 862.730 371.615 862.745 ;
        RECT 372.205 862.730 372.535 862.745 ;
        RECT 371.285 862.430 372.535 862.730 ;
        RECT 371.285 862.415 371.615 862.430 ;
        RECT 372.205 862.415 372.535 862.430 ;
        RECT 371.285 766.170 371.615 766.185 ;
        RECT 372.205 766.170 372.535 766.185 ;
        RECT 371.285 765.870 372.535 766.170 ;
        RECT 371.285 765.855 371.615 765.870 ;
        RECT 372.205 765.855 372.535 765.870 ;
        RECT 372.205 628.130 372.535 628.145 ;
        RECT 373.125 628.130 373.455 628.145 ;
        RECT 372.205 627.830 373.455 628.130 ;
        RECT 372.205 627.815 372.535 627.830 ;
        RECT 373.125 627.815 373.455 627.830 ;
        RECT 372.205 620.650 372.535 620.665 ;
        RECT 373.585 620.650 373.915 620.665 ;
        RECT 372.205 620.350 373.915 620.650 ;
        RECT 372.205 620.335 372.535 620.350 ;
        RECT 373.585 620.335 373.915 620.350 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.570 20.640 931.890 20.700 ;
        RECT 447.280 20.500 931.890 20.640 ;
        RECT 400.270 20.300 400.590 20.360 ;
        RECT 447.280 20.300 447.420 20.500 ;
        RECT 931.570 20.440 931.890 20.500 ;
        RECT 400.270 20.160 447.420 20.300 ;
        RECT 400.270 20.100 400.590 20.160 ;
      LAYER via ;
        RECT 400.300 20.100 400.560 20.360 ;
        RECT 931.600 20.440 931.860 20.700 ;
      LAYER met2 ;
        RECT 937.190 1600.450 937.470 1604.000 ;
        RECT 931.660 1600.310 937.470 1600.450 ;
        RECT 931.660 20.730 931.800 1600.310 ;
        RECT 937.190 1600.000 937.470 1600.310 ;
        RECT 931.600 20.410 931.860 20.730 ;
        RECT 400.300 20.245 400.560 20.390 ;
        RECT 389.250 19.875 389.530 20.245 ;
        RECT 400.290 19.875 400.570 20.245 ;
        RECT 389.320 2.400 389.460 19.875 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 389.250 19.920 389.530 20.200 ;
        RECT 400.290 19.920 400.570 20.200 ;
      LAYER met3 ;
        RECT 389.225 20.210 389.555 20.225 ;
        RECT 400.265 20.210 400.595 20.225 ;
        RECT 389.225 19.910 400.595 20.210 ;
        RECT 389.225 19.895 389.555 19.910 ;
        RECT 400.265 19.895 400.595 19.910 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 1593.820 413.930 1593.880 ;
        RECT 966.070 1593.820 966.390 1593.880 ;
        RECT 413.610 1593.680 966.390 1593.820 ;
        RECT 413.610 1593.620 413.930 1593.680 ;
        RECT 966.070 1593.620 966.390 1593.680 ;
        RECT 407.170 20.640 407.490 20.700 ;
        RECT 413.610 20.640 413.930 20.700 ;
        RECT 407.170 20.500 413.930 20.640 ;
        RECT 407.170 20.440 407.490 20.500 ;
        RECT 413.610 20.440 413.930 20.500 ;
      LAYER via ;
        RECT 413.640 1593.620 413.900 1593.880 ;
        RECT 966.100 1593.620 966.360 1593.880 ;
        RECT 407.200 20.440 407.460 20.700 ;
        RECT 413.640 20.440 413.900 20.700 ;
      LAYER met2 ;
        RECT 966.170 1600.380 966.450 1604.000 ;
        RECT 966.160 1600.000 966.450 1600.380 ;
        RECT 966.160 1593.910 966.300 1600.000 ;
        RECT 413.640 1593.590 413.900 1593.910 ;
        RECT 966.100 1593.590 966.360 1593.910 ;
        RECT 413.700 20.730 413.840 1593.590 ;
        RECT 407.200 20.410 407.460 20.730 ;
        RECT 413.640 20.410 413.900 20.730 ;
        RECT 407.260 2.400 407.400 20.410 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 406.710 20.640 407.030 20.700 ;
        RECT 375.980 20.500 407.030 20.640 ;
        RECT 68.150 20.300 68.470 20.360 ;
        RECT 375.980 20.300 376.120 20.500 ;
        RECT 406.710 20.440 407.030 20.500 ;
        RECT 68.150 20.160 376.120 20.300 ;
        RECT 68.150 20.100 68.470 20.160 ;
      LAYER via ;
        RECT 68.180 20.100 68.440 20.360 ;
        RECT 406.740 20.440 407.000 20.700 ;
      LAYER met2 ;
        RECT 411.410 1600.450 411.690 1604.000 ;
        RECT 407.260 1600.310 411.690 1600.450 ;
        RECT 407.260 21.490 407.400 1600.310 ;
        RECT 411.410 1600.000 411.690 1600.310 ;
        RECT 406.800 21.350 407.400 21.490 ;
        RECT 406.800 20.730 406.940 21.350 ;
        RECT 406.740 20.410 407.000 20.730 ;
        RECT 68.180 20.070 68.440 20.390 ;
        RECT 68.240 2.400 68.380 20.070 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 424.650 19.960 424.970 20.020 ;
        RECT 447.190 19.960 447.510 20.020 ;
        RECT 993.670 19.960 993.990 20.020 ;
        RECT 424.650 19.820 447.510 19.960 ;
        RECT 424.650 19.760 424.970 19.820 ;
        RECT 447.190 19.760 447.510 19.820 ;
        RECT 466.600 19.820 993.990 19.960 ;
        RECT 449.490 19.620 449.810 19.680 ;
        RECT 466.600 19.620 466.740 19.820 ;
        RECT 993.670 19.760 993.990 19.820 ;
        RECT 449.490 19.480 466.740 19.620 ;
        RECT 449.490 19.420 449.810 19.480 ;
      LAYER via ;
        RECT 424.680 19.760 424.940 20.020 ;
        RECT 447.220 19.760 447.480 20.020 ;
        RECT 449.520 19.420 449.780 19.680 ;
        RECT 993.700 19.760 993.960 20.020 ;
      LAYER met2 ;
        RECT 995.610 1600.450 995.890 1604.000 ;
        RECT 993.760 1600.310 995.890 1600.450 ;
        RECT 993.760 20.050 993.900 1600.310 ;
        RECT 995.610 1600.000 995.890 1600.310 ;
        RECT 424.680 19.730 424.940 20.050 ;
        RECT 447.220 19.730 447.480 20.050 ;
        RECT 993.700 19.730 993.960 20.050 ;
        RECT 424.740 2.400 424.880 19.730 ;
        RECT 447.280 19.565 447.420 19.730 ;
        RECT 449.520 19.565 449.780 19.710 ;
        RECT 447.210 19.195 447.490 19.565 ;
        RECT 449.510 19.195 449.790 19.565 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 447.210 19.240 447.490 19.520 ;
        RECT 449.510 19.240 449.790 19.520 ;
      LAYER met3 ;
        RECT 447.185 19.530 447.515 19.545 ;
        RECT 449.485 19.530 449.815 19.545 ;
        RECT 447.185 19.230 449.815 19.530 ;
        RECT 447.185 19.215 447.515 19.230 ;
        RECT 449.485 19.215 449.815 19.230 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1024.490 1593.140 1024.810 1593.200 ;
        RECT 472.580 1593.000 1024.810 1593.140 ;
        RECT 447.650 1592.460 447.970 1592.520 ;
        RECT 472.580 1592.460 472.720 1593.000 ;
        RECT 1024.490 1592.940 1024.810 1593.000 ;
        RECT 447.650 1592.320 472.720 1592.460 ;
        RECT 447.650 1592.260 447.970 1592.320 ;
        RECT 446.730 1014.460 447.050 1014.520 ;
        RECT 447.650 1014.460 447.970 1014.520 ;
        RECT 446.730 1014.320 447.970 1014.460 ;
        RECT 446.730 1014.260 447.050 1014.320 ;
        RECT 447.650 1014.260 447.970 1014.320 ;
        RECT 446.730 979.920 447.050 980.180 ;
        RECT 446.820 979.440 446.960 979.920 ;
        RECT 447.190 979.440 447.510 979.500 ;
        RECT 446.820 979.300 447.510 979.440 ;
        RECT 447.190 979.240 447.510 979.300 ;
        RECT 447.190 869.620 447.510 869.680 ;
        RECT 448.110 869.620 448.430 869.680 ;
        RECT 447.190 869.480 448.430 869.620 ;
        RECT 447.190 869.420 447.510 869.480 ;
        RECT 448.110 869.420 448.430 869.480 ;
        RECT 447.190 787.140 447.510 787.400 ;
        RECT 447.280 786.720 447.420 787.140 ;
        RECT 447.190 786.460 447.510 786.720 ;
        RECT 446.270 772.720 446.590 772.780 ;
        RECT 447.650 772.720 447.970 772.780 ;
        RECT 446.270 772.580 447.970 772.720 ;
        RECT 446.270 772.520 446.590 772.580 ;
        RECT 447.650 772.520 447.970 772.580 ;
        RECT 447.190 689.900 447.510 690.160 ;
        RECT 447.280 689.420 447.420 689.900 ;
        RECT 447.650 689.420 447.970 689.480 ;
        RECT 447.280 689.280 447.970 689.420 ;
        RECT 447.650 689.220 447.970 689.280 ;
        RECT 447.650 642.160 447.970 642.220 ;
        RECT 447.280 642.020 447.970 642.160 ;
        RECT 447.280 641.540 447.420 642.020 ;
        RECT 447.650 641.960 447.970 642.020 ;
        RECT 447.190 641.280 447.510 641.540 ;
        RECT 447.190 620.400 447.510 620.460 ;
        RECT 448.110 620.400 448.430 620.460 ;
        RECT 447.190 620.260 448.430 620.400 ;
        RECT 447.190 620.200 447.510 620.260 ;
        RECT 448.110 620.200 448.430 620.260 ;
        RECT 448.110 593.340 448.430 593.600 ;
        RECT 447.650 592.860 447.970 592.920 ;
        RECT 448.200 592.860 448.340 593.340 ;
        RECT 447.650 592.720 448.340 592.860 ;
        RECT 447.650 592.660 447.970 592.720 ;
        RECT 447.650 545.600 447.970 545.660 ;
        RECT 447.280 545.460 447.970 545.600 ;
        RECT 447.280 544.980 447.420 545.460 ;
        RECT 447.650 545.400 447.970 545.460 ;
        RECT 447.190 544.720 447.510 544.980 ;
        RECT 446.270 524.180 446.590 524.240 ;
        RECT 447.190 524.180 447.510 524.240 ;
        RECT 446.270 524.040 447.510 524.180 ;
        RECT 446.270 523.980 446.590 524.040 ;
        RECT 447.190 523.980 447.510 524.040 ;
        RECT 446.270 476.240 446.590 476.300 ;
        RECT 446.730 476.240 447.050 476.300 ;
        RECT 446.270 476.100 447.050 476.240 ;
        RECT 446.270 476.040 446.590 476.100 ;
        RECT 446.730 476.040 447.050 476.100 ;
        RECT 447.650 400.560 447.970 400.820 ;
        RECT 447.740 400.140 447.880 400.560 ;
        RECT 447.650 399.880 447.970 400.140 ;
        RECT 447.190 255.240 447.510 255.300 ;
        RECT 448.110 255.240 448.430 255.300 ;
        RECT 447.190 255.100 448.430 255.240 ;
        RECT 447.190 255.040 447.510 255.100 ;
        RECT 448.110 255.040 448.430 255.100 ;
        RECT 446.730 241.300 447.050 241.360 ;
        RECT 448.110 241.300 448.430 241.360 ;
        RECT 446.730 241.160 448.430 241.300 ;
        RECT 446.730 241.100 447.050 241.160 ;
        RECT 448.110 241.100 448.430 241.160 ;
        RECT 446.730 193.360 447.050 193.420 ;
        RECT 447.650 193.360 447.970 193.420 ;
        RECT 446.730 193.220 447.970 193.360 ;
        RECT 446.730 193.160 447.050 193.220 ;
        RECT 447.650 193.160 447.970 193.220 ;
        RECT 445.810 131.140 446.130 131.200 ;
        RECT 446.270 131.140 446.590 131.200 ;
        RECT 445.810 131.000 446.590 131.140 ;
        RECT 445.810 130.940 446.130 131.000 ;
        RECT 446.270 130.940 446.590 131.000 ;
        RECT 445.810 107.000 446.130 107.060 ;
        RECT 447.190 107.000 447.510 107.060 ;
        RECT 445.810 106.860 447.510 107.000 ;
        RECT 445.810 106.800 446.130 106.860 ;
        RECT 447.190 106.800 447.510 106.860 ;
        RECT 446.730 41.720 447.050 41.780 ;
        RECT 447.190 41.720 447.510 41.780 ;
        RECT 446.730 41.580 447.510 41.720 ;
        RECT 446.730 41.520 447.050 41.580 ;
        RECT 447.190 41.520 447.510 41.580 ;
        RECT 442.590 5.680 442.910 5.740 ;
        RECT 446.730 5.680 447.050 5.740 ;
        RECT 442.590 5.540 447.050 5.680 ;
        RECT 442.590 5.480 442.910 5.540 ;
        RECT 446.730 5.480 447.050 5.540 ;
      LAYER via ;
        RECT 447.680 1592.260 447.940 1592.520 ;
        RECT 1024.520 1592.940 1024.780 1593.200 ;
        RECT 446.760 1014.260 447.020 1014.520 ;
        RECT 447.680 1014.260 447.940 1014.520 ;
        RECT 446.760 979.920 447.020 980.180 ;
        RECT 447.220 979.240 447.480 979.500 ;
        RECT 447.220 869.420 447.480 869.680 ;
        RECT 448.140 869.420 448.400 869.680 ;
        RECT 447.220 787.140 447.480 787.400 ;
        RECT 447.220 786.460 447.480 786.720 ;
        RECT 446.300 772.520 446.560 772.780 ;
        RECT 447.680 772.520 447.940 772.780 ;
        RECT 447.220 689.900 447.480 690.160 ;
        RECT 447.680 689.220 447.940 689.480 ;
        RECT 447.680 641.960 447.940 642.220 ;
        RECT 447.220 641.280 447.480 641.540 ;
        RECT 447.220 620.200 447.480 620.460 ;
        RECT 448.140 620.200 448.400 620.460 ;
        RECT 448.140 593.340 448.400 593.600 ;
        RECT 447.680 592.660 447.940 592.920 ;
        RECT 447.680 545.400 447.940 545.660 ;
        RECT 447.220 544.720 447.480 544.980 ;
        RECT 446.300 523.980 446.560 524.240 ;
        RECT 447.220 523.980 447.480 524.240 ;
        RECT 446.300 476.040 446.560 476.300 ;
        RECT 446.760 476.040 447.020 476.300 ;
        RECT 447.680 400.560 447.940 400.820 ;
        RECT 447.680 399.880 447.940 400.140 ;
        RECT 447.220 255.040 447.480 255.300 ;
        RECT 448.140 255.040 448.400 255.300 ;
        RECT 446.760 241.100 447.020 241.360 ;
        RECT 448.140 241.100 448.400 241.360 ;
        RECT 446.760 193.160 447.020 193.420 ;
        RECT 447.680 193.160 447.940 193.420 ;
        RECT 445.840 130.940 446.100 131.200 ;
        RECT 446.300 130.940 446.560 131.200 ;
        RECT 445.840 106.800 446.100 107.060 ;
        RECT 447.220 106.800 447.480 107.060 ;
        RECT 446.760 41.520 447.020 41.780 ;
        RECT 447.220 41.520 447.480 41.780 ;
        RECT 442.620 5.480 442.880 5.740 ;
        RECT 446.760 5.480 447.020 5.740 ;
      LAYER met2 ;
        RECT 1024.590 1600.380 1024.870 1604.000 ;
        RECT 1024.580 1600.000 1024.870 1600.380 ;
        RECT 1024.580 1593.230 1024.720 1600.000 ;
        RECT 1024.520 1592.910 1024.780 1593.230 ;
        RECT 447.680 1592.230 447.940 1592.550 ;
        RECT 447.740 1511.370 447.880 1592.230 ;
        RECT 447.280 1511.230 447.880 1511.370 ;
        RECT 447.280 1510.690 447.420 1511.230 ;
        RECT 447.280 1510.550 447.880 1510.690 ;
        RECT 447.740 1463.090 447.880 1510.550 ;
        RECT 447.740 1462.950 448.340 1463.090 ;
        RECT 448.200 1462.410 448.340 1462.950 ;
        RECT 447.740 1462.270 448.340 1462.410 ;
        RECT 447.740 1414.810 447.880 1462.270 ;
        RECT 447.280 1414.670 447.880 1414.810 ;
        RECT 447.280 1414.130 447.420 1414.670 ;
        RECT 447.280 1413.990 447.880 1414.130 ;
        RECT 447.740 1366.530 447.880 1413.990 ;
        RECT 447.740 1366.390 448.340 1366.530 ;
        RECT 448.200 1269.290 448.340 1366.390 ;
        RECT 447.740 1269.150 448.340 1269.290 ;
        RECT 447.740 1221.690 447.880 1269.150 ;
        RECT 447.280 1221.550 447.880 1221.690 ;
        RECT 447.280 1221.010 447.420 1221.550 ;
        RECT 447.280 1220.870 447.880 1221.010 ;
        RECT 447.740 1173.410 447.880 1220.870 ;
        RECT 447.740 1173.270 448.340 1173.410 ;
        RECT 448.200 1076.170 448.340 1173.270 ;
        RECT 447.740 1076.030 448.340 1076.170 ;
        RECT 447.740 1014.550 447.880 1076.030 ;
        RECT 446.760 1014.230 447.020 1014.550 ;
        RECT 447.680 1014.230 447.940 1014.550 ;
        RECT 446.820 980.210 446.960 1014.230 ;
        RECT 446.760 979.890 447.020 980.210 ;
        RECT 447.220 979.210 447.480 979.530 ;
        RECT 447.280 869.710 447.420 979.210 ;
        RECT 447.220 869.390 447.480 869.710 ;
        RECT 448.140 869.390 448.400 869.710 ;
        RECT 448.200 835.450 448.340 869.390 ;
        RECT 447.740 835.310 448.340 835.450 ;
        RECT 447.740 834.770 447.880 835.310 ;
        RECT 447.280 834.630 447.880 834.770 ;
        RECT 447.280 787.430 447.420 834.630 ;
        RECT 447.220 787.110 447.480 787.430 ;
        RECT 447.220 786.430 447.480 786.750 ;
        RECT 447.280 785.810 447.420 786.430 ;
        RECT 447.280 785.670 447.880 785.810 ;
        RECT 447.740 772.810 447.880 785.670 ;
        RECT 446.300 772.490 446.560 772.810 ;
        RECT 447.680 772.490 447.940 772.810 ;
        RECT 446.360 724.725 446.500 772.490 ;
        RECT 446.290 724.355 446.570 724.725 ;
        RECT 447.210 724.355 447.490 724.725 ;
        RECT 447.280 690.190 447.420 724.355 ;
        RECT 447.220 689.870 447.480 690.190 ;
        RECT 447.680 689.190 447.940 689.510 ;
        RECT 447.740 642.250 447.880 689.190 ;
        RECT 447.680 641.930 447.940 642.250 ;
        RECT 447.220 641.250 447.480 641.570 ;
        RECT 447.280 620.490 447.420 641.250 ;
        RECT 447.220 620.170 447.480 620.490 ;
        RECT 448.140 620.170 448.400 620.490 ;
        RECT 448.200 593.630 448.340 620.170 ;
        RECT 448.140 593.310 448.400 593.630 ;
        RECT 447.680 592.630 447.940 592.950 ;
        RECT 447.740 545.690 447.880 592.630 ;
        RECT 447.680 545.370 447.940 545.690 ;
        RECT 447.220 544.690 447.480 545.010 ;
        RECT 447.280 524.270 447.420 544.690 ;
        RECT 446.300 523.950 446.560 524.270 ;
        RECT 447.220 523.950 447.480 524.270 ;
        RECT 446.360 476.330 446.500 523.950 ;
        RECT 446.300 476.010 446.560 476.330 ;
        RECT 446.760 476.010 447.020 476.330 ;
        RECT 446.820 447.170 446.960 476.010 ;
        RECT 446.820 447.030 447.880 447.170 ;
        RECT 447.740 400.850 447.880 447.030 ;
        RECT 447.680 400.530 447.940 400.850 ;
        RECT 447.680 399.850 447.940 400.170 ;
        RECT 447.740 351.970 447.880 399.850 ;
        RECT 447.280 351.830 447.880 351.970 ;
        RECT 447.280 351.290 447.420 351.830 ;
        RECT 447.280 351.150 447.880 351.290 ;
        RECT 447.740 255.410 447.880 351.150 ;
        RECT 447.280 255.330 447.880 255.410 ;
        RECT 447.220 255.270 447.880 255.330 ;
        RECT 447.220 255.010 447.480 255.270 ;
        RECT 448.140 255.010 448.400 255.330 ;
        RECT 447.280 254.855 447.420 255.010 ;
        RECT 448.200 241.390 448.340 255.010 ;
        RECT 446.760 241.070 447.020 241.390 ;
        RECT 448.140 241.070 448.400 241.390 ;
        RECT 446.820 193.450 446.960 241.070 ;
        RECT 446.760 193.130 447.020 193.450 ;
        RECT 447.680 193.130 447.940 193.450 ;
        RECT 447.740 158.965 447.880 193.130 ;
        RECT 447.670 158.595 447.950 158.965 ;
        RECT 446.290 131.395 446.570 131.765 ;
        RECT 446.360 131.230 446.500 131.395 ;
        RECT 445.840 130.910 446.100 131.230 ;
        RECT 446.300 130.910 446.560 131.230 ;
        RECT 445.900 107.090 446.040 130.910 ;
        RECT 445.840 106.770 446.100 107.090 ;
        RECT 447.220 106.770 447.480 107.090 ;
        RECT 447.280 41.810 447.420 106.770 ;
        RECT 446.760 41.490 447.020 41.810 ;
        RECT 447.220 41.490 447.480 41.810 ;
        RECT 446.820 5.770 446.960 41.490 ;
        RECT 442.620 5.450 442.880 5.770 ;
        RECT 446.760 5.450 447.020 5.770 ;
        RECT 442.680 2.400 442.820 5.450 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 446.290 724.400 446.570 724.680 ;
        RECT 447.210 724.400 447.490 724.680 ;
        RECT 447.670 158.640 447.950 158.920 ;
        RECT 446.290 131.440 446.570 131.720 ;
      LAYER met3 ;
        RECT 446.265 724.690 446.595 724.705 ;
        RECT 447.185 724.690 447.515 724.705 ;
        RECT 446.265 724.390 447.515 724.690 ;
        RECT 446.265 724.375 446.595 724.390 ;
        RECT 447.185 724.375 447.515 724.390 ;
        RECT 446.470 158.930 446.850 158.940 ;
        RECT 447.645 158.930 447.975 158.945 ;
        RECT 446.470 158.630 447.975 158.930 ;
        RECT 446.470 158.620 446.850 158.630 ;
        RECT 447.645 158.615 447.975 158.630 ;
        RECT 446.265 131.740 446.595 131.745 ;
        RECT 446.265 131.730 446.850 131.740 ;
        RECT 446.040 131.430 446.850 131.730 ;
        RECT 446.265 131.420 446.850 131.430 ;
        RECT 446.265 131.415 446.595 131.420 ;
      LAYER via3 ;
        RECT 446.500 158.620 446.820 158.940 ;
        RECT 446.500 131.420 446.820 131.740 ;
      LAYER met4 ;
        RECT 446.495 158.615 446.825 158.945 ;
        RECT 446.510 131.745 446.810 158.615 ;
        RECT 446.495 131.415 446.825 131.745 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1054.030 1600.450 1054.310 1604.000 ;
        RECT 1048.960 1600.310 1054.310 1600.450 ;
        RECT 1048.960 18.205 1049.100 1600.310 ;
        RECT 1054.030 1600.000 1054.310 1600.310 ;
        RECT 460.550 17.835 460.830 18.205 ;
        RECT 1048.890 17.835 1049.170 18.205 ;
        RECT 460.620 2.400 460.760 17.835 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 460.550 17.880 460.830 18.160 ;
        RECT 1048.890 17.880 1049.170 18.160 ;
      LAYER met3 ;
        RECT 460.525 18.170 460.855 18.185 ;
        RECT 1048.865 18.170 1049.195 18.185 ;
        RECT 460.525 17.870 1049.195 18.170 ;
        RECT 460.525 17.855 460.855 17.870 ;
        RECT 1048.865 17.855 1049.195 17.870 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 1592.460 482.930 1592.520 ;
        RECT 1082.910 1592.460 1083.230 1592.520 ;
        RECT 482.610 1592.320 1083.230 1592.460 ;
        RECT 482.610 1592.260 482.930 1592.320 ;
        RECT 1082.910 1592.260 1083.230 1592.320 ;
        RECT 478.470 18.940 478.790 19.000 ;
        RECT 482.610 18.940 482.930 19.000 ;
        RECT 478.470 18.800 482.930 18.940 ;
        RECT 478.470 18.740 478.790 18.800 ;
        RECT 482.610 18.740 482.930 18.800 ;
      LAYER via ;
        RECT 482.640 1592.260 482.900 1592.520 ;
        RECT 1082.940 1592.260 1083.200 1592.520 ;
        RECT 478.500 18.740 478.760 19.000 ;
        RECT 482.640 18.740 482.900 19.000 ;
      LAYER met2 ;
        RECT 1083.010 1600.380 1083.290 1604.000 ;
        RECT 1083.000 1600.000 1083.290 1600.380 ;
        RECT 1083.000 1592.550 1083.140 1600.000 ;
        RECT 482.640 1592.230 482.900 1592.550 ;
        RECT 1082.940 1592.230 1083.200 1592.550 ;
        RECT 482.700 19.030 482.840 1592.230 ;
        RECT 478.500 18.710 478.760 19.030 ;
        RECT 482.640 18.710 482.900 19.030 ;
        RECT 478.560 2.400 478.700 18.710 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.450 1600.450 1112.730 1604.000 ;
        RECT 1111.060 1600.310 1112.730 1600.450 ;
        RECT 1111.060 17.525 1111.200 1600.310 ;
        RECT 1112.450 1600.000 1112.730 1600.310 ;
        RECT 496.430 17.155 496.710 17.525 ;
        RECT 1110.990 17.155 1111.270 17.525 ;
        RECT 496.500 2.400 496.640 17.155 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 496.430 17.200 496.710 17.480 ;
        RECT 1110.990 17.200 1111.270 17.480 ;
      LAYER met3 ;
        RECT 496.405 17.490 496.735 17.505 ;
        RECT 1110.965 17.490 1111.295 17.505 ;
        RECT 496.405 17.190 1111.295 17.490 ;
        RECT 496.405 17.175 496.735 17.190 ;
        RECT 1110.965 17.175 1111.295 17.190 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 1591.440 517.430 1591.500 ;
        RECT 1141.330 1591.440 1141.650 1591.500 ;
        RECT 517.110 1591.300 1141.650 1591.440 ;
        RECT 517.110 1591.240 517.430 1591.300 ;
        RECT 1141.330 1591.240 1141.650 1591.300 ;
        RECT 513.890 19.280 514.210 19.340 ;
        RECT 517.110 19.280 517.430 19.340 ;
        RECT 513.890 19.140 517.430 19.280 ;
        RECT 513.890 19.080 514.210 19.140 ;
        RECT 517.110 19.080 517.430 19.140 ;
      LAYER via ;
        RECT 517.140 1591.240 517.400 1591.500 ;
        RECT 1141.360 1591.240 1141.620 1591.500 ;
        RECT 513.920 19.080 514.180 19.340 ;
        RECT 517.140 19.080 517.400 19.340 ;
      LAYER met2 ;
        RECT 1141.430 1600.380 1141.710 1604.000 ;
        RECT 1141.420 1600.000 1141.710 1600.380 ;
        RECT 1141.420 1591.530 1141.560 1600.000 ;
        RECT 517.140 1591.210 517.400 1591.530 ;
        RECT 1141.360 1591.210 1141.620 1591.530 ;
        RECT 517.200 19.370 517.340 1591.210 ;
        RECT 513.920 19.050 514.180 19.370 ;
        RECT 517.140 19.050 517.400 19.370 ;
        RECT 513.980 2.400 514.120 19.050 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.810 1591.100 538.130 1591.160 ;
        RECT 1170.770 1591.100 1171.090 1591.160 ;
        RECT 537.810 1590.960 1171.090 1591.100 ;
        RECT 537.810 1590.900 538.130 1590.960 ;
        RECT 1170.770 1590.900 1171.090 1590.960 ;
        RECT 531.830 17.920 532.150 17.980 ;
        RECT 537.810 17.920 538.130 17.980 ;
        RECT 531.830 17.780 538.130 17.920 ;
        RECT 531.830 17.720 532.150 17.780 ;
        RECT 537.810 17.720 538.130 17.780 ;
      LAYER via ;
        RECT 537.840 1590.900 538.100 1591.160 ;
        RECT 1170.800 1590.900 1171.060 1591.160 ;
        RECT 531.860 17.720 532.120 17.980 ;
        RECT 537.840 17.720 538.100 17.980 ;
      LAYER met2 ;
        RECT 1170.870 1600.380 1171.150 1604.000 ;
        RECT 1170.860 1600.000 1171.150 1600.380 ;
        RECT 1170.860 1591.190 1171.000 1600.000 ;
        RECT 537.840 1590.870 538.100 1591.190 ;
        RECT 1170.800 1590.870 1171.060 1591.190 ;
        RECT 537.900 18.010 538.040 1590.870 ;
        RECT 531.860 17.690 532.120 18.010 ;
        RECT 537.840 17.690 538.100 18.010 ;
        RECT 531.920 2.400 532.060 17.690 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 580.130 18.940 580.450 19.000 ;
        RECT 1193.770 18.940 1194.090 19.000 ;
        RECT 580.130 18.800 1194.090 18.940 ;
        RECT 580.130 18.740 580.450 18.800 ;
        RECT 1193.770 18.740 1194.090 18.800 ;
        RECT 549.770 17.920 550.090 17.980 ;
        RECT 568.630 17.920 568.950 17.980 ;
        RECT 549.770 17.780 568.950 17.920 ;
        RECT 549.770 17.720 550.090 17.780 ;
        RECT 568.630 17.720 568.950 17.780 ;
        RECT 570.470 17.920 570.790 17.980 ;
        RECT 580.130 17.920 580.450 17.980 ;
        RECT 570.470 17.780 580.450 17.920 ;
        RECT 570.470 17.720 570.790 17.780 ;
        RECT 580.130 17.720 580.450 17.780 ;
      LAYER via ;
        RECT 580.160 18.740 580.420 19.000 ;
        RECT 1193.800 18.740 1194.060 19.000 ;
        RECT 549.800 17.720 550.060 17.980 ;
        RECT 568.660 17.720 568.920 17.980 ;
        RECT 570.500 17.720 570.760 17.980 ;
        RECT 580.160 17.720 580.420 17.980 ;
      LAYER met2 ;
        RECT 1199.850 1600.450 1200.130 1604.000 ;
        RECT 1193.860 1600.310 1200.130 1600.450 ;
        RECT 1193.860 19.030 1194.000 1600.310 ;
        RECT 1199.850 1600.000 1200.130 1600.310 ;
        RECT 568.720 18.630 570.700 18.770 ;
        RECT 580.160 18.710 580.420 19.030 ;
        RECT 1193.800 18.710 1194.060 19.030 ;
        RECT 568.720 18.010 568.860 18.630 ;
        RECT 570.560 18.010 570.700 18.630 ;
        RECT 580.220 18.010 580.360 18.710 ;
        RECT 549.800 17.690 550.060 18.010 ;
        RECT 568.660 17.690 568.920 18.010 ;
        RECT 570.500 17.690 570.760 18.010 ;
        RECT 580.160 17.690 580.420 18.010 ;
        RECT 549.860 2.400 550.000 17.690 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 1590.420 572.630 1590.480 ;
        RECT 1229.190 1590.420 1229.510 1590.480 ;
        RECT 572.310 1590.280 1229.510 1590.420 ;
        RECT 572.310 1590.220 572.630 1590.280 ;
        RECT 1229.190 1590.220 1229.510 1590.280 ;
        RECT 567.710 18.940 568.030 19.000 ;
        RECT 572.310 18.940 572.630 19.000 ;
        RECT 567.710 18.800 572.630 18.940 ;
        RECT 567.710 18.740 568.030 18.800 ;
        RECT 572.310 18.740 572.630 18.800 ;
      LAYER via ;
        RECT 572.340 1590.220 572.600 1590.480 ;
        RECT 1229.220 1590.220 1229.480 1590.480 ;
        RECT 567.740 18.740 568.000 19.000 ;
        RECT 572.340 18.740 572.600 19.000 ;
      LAYER met2 ;
        RECT 1229.290 1600.380 1229.570 1604.000 ;
        RECT 1229.280 1600.000 1229.570 1600.380 ;
        RECT 1229.280 1590.510 1229.420 1600.000 ;
        RECT 572.340 1590.190 572.600 1590.510 ;
        RECT 1229.220 1590.190 1229.480 1590.510 ;
        RECT 572.400 19.030 572.540 1590.190 ;
        RECT 567.740 18.710 568.000 19.030 ;
        RECT 572.340 18.710 572.600 19.030 ;
        RECT 567.800 2.400 567.940 18.710 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 18.260 585.970 18.320 ;
        RECT 585.650 18.120 602.900 18.260 ;
        RECT 585.650 18.060 585.970 18.120 ;
        RECT 602.760 17.920 602.900 18.120 ;
        RECT 1255.870 17.920 1256.190 17.980 ;
        RECT 602.760 17.780 613.940 17.920 ;
        RECT 613.800 17.580 613.940 17.780 ;
        RECT 615.180 17.780 1256.190 17.920 ;
        RECT 615.180 17.580 615.320 17.780 ;
        RECT 1255.870 17.720 1256.190 17.780 ;
        RECT 613.800 17.440 615.320 17.580 ;
      LAYER via ;
        RECT 585.680 18.060 585.940 18.320 ;
        RECT 1255.900 17.720 1256.160 17.980 ;
      LAYER met2 ;
        RECT 1258.270 1600.450 1258.550 1604.000 ;
        RECT 1255.960 1600.310 1258.550 1600.450 ;
        RECT 585.680 18.030 585.940 18.350 ;
        RECT 585.740 2.400 585.880 18.030 ;
        RECT 1255.960 18.010 1256.100 1600.310 ;
        RECT 1258.270 1600.000 1258.550 1600.310 ;
        RECT 1255.900 17.690 1256.160 18.010 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 91.610 19.620 91.930 19.680 ;
        RECT 448.110 19.620 448.430 19.680 ;
        RECT 91.610 19.480 448.430 19.620 ;
        RECT 91.610 19.420 91.930 19.480 ;
        RECT 448.110 19.420 448.430 19.480 ;
      LAYER via ;
        RECT 91.640 19.420 91.900 19.680 ;
        RECT 448.140 19.420 448.400 19.680 ;
      LAYER met2 ;
        RECT 450.510 1600.450 450.790 1604.000 ;
        RECT 448.660 1600.310 450.790 1600.450 ;
        RECT 448.660 20.810 448.800 1600.310 ;
        RECT 450.510 1600.000 450.790 1600.310 ;
        RECT 448.200 20.670 448.800 20.810 ;
        RECT 448.200 19.710 448.340 20.670 ;
        RECT 91.640 19.390 91.900 19.710 ;
        RECT 448.140 19.390 448.400 19.710 ;
        RECT 91.700 2.400 91.840 19.390 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 603.130 18.260 603.450 18.320 ;
        RECT 606.810 18.260 607.130 18.320 ;
        RECT 603.130 18.120 607.130 18.260 ;
        RECT 603.130 18.060 603.450 18.120 ;
        RECT 606.810 18.060 607.130 18.120 ;
      LAYER via ;
        RECT 603.160 18.060 603.420 18.320 ;
        RECT 606.840 18.060 607.100 18.320 ;
      LAYER met2 ;
        RECT 1287.710 1600.380 1287.990 1604.000 ;
        RECT 1287.700 1600.000 1287.990 1600.380 ;
        RECT 1287.700 1591.045 1287.840 1600.000 ;
        RECT 606.830 1590.675 607.110 1591.045 ;
        RECT 1287.630 1590.675 1287.910 1591.045 ;
        RECT 606.900 18.350 607.040 1590.675 ;
        RECT 603.160 18.030 603.420 18.350 ;
        RECT 606.840 18.030 607.100 18.350 ;
        RECT 603.220 2.400 603.360 18.030 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 606.830 1590.720 607.110 1591.000 ;
        RECT 1287.630 1590.720 1287.910 1591.000 ;
      LAYER met3 ;
        RECT 606.805 1591.010 607.135 1591.025 ;
        RECT 1287.605 1591.010 1287.935 1591.025 ;
        RECT 606.805 1590.710 1287.935 1591.010 ;
        RECT 606.805 1590.695 607.135 1590.710 ;
        RECT 1287.605 1590.695 1287.935 1590.710 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 621.070 17.580 621.390 17.640 ;
        RECT 1311.070 17.580 1311.390 17.640 ;
        RECT 621.070 17.440 1311.390 17.580 ;
        RECT 621.070 17.380 621.390 17.440 ;
        RECT 1311.070 17.380 1311.390 17.440 ;
      LAYER via ;
        RECT 621.100 17.380 621.360 17.640 ;
        RECT 1311.100 17.380 1311.360 17.640 ;
      LAYER met2 ;
        RECT 1316.690 1600.450 1316.970 1604.000 ;
        RECT 1311.160 1600.310 1316.970 1600.450 ;
        RECT 1311.160 17.670 1311.300 1600.310 ;
        RECT 1316.690 1600.000 1316.970 1600.310 ;
        RECT 621.100 17.350 621.360 17.670 ;
        RECT 1311.100 17.350 1311.360 17.670 ;
        RECT 621.160 2.400 621.300 17.350 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 477.550 19.280 477.870 19.340 ;
        RECT 139.080 19.140 477.870 19.280 ;
        RECT 115.530 18.940 115.850 19.000 ;
        RECT 139.080 18.940 139.220 19.140 ;
        RECT 477.550 19.080 477.870 19.140 ;
        RECT 115.530 18.800 139.220 18.940 ;
        RECT 115.530 18.740 115.850 18.800 ;
      LAYER via ;
        RECT 115.560 18.740 115.820 19.000 ;
        RECT 477.580 19.080 477.840 19.340 ;
      LAYER met2 ;
        RECT 489.610 1600.450 489.890 1604.000 ;
        RECT 483.160 1600.310 489.890 1600.450 ;
        RECT 483.160 19.565 483.300 1600.310 ;
        RECT 489.610 1600.000 489.890 1600.310 ;
        RECT 477.570 19.195 477.850 19.565 ;
        RECT 483.090 19.195 483.370 19.565 ;
        RECT 477.580 19.050 477.840 19.195 ;
        RECT 115.560 18.710 115.820 19.030 ;
        RECT 115.620 2.400 115.760 18.710 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 477.570 19.240 477.850 19.520 ;
        RECT 483.090 19.240 483.370 19.520 ;
      LAYER met3 ;
        RECT 477.545 19.530 477.875 19.545 ;
        RECT 483.065 19.530 483.395 19.545 ;
        RECT 477.545 19.230 483.395 19.530 ;
        RECT 477.545 19.215 477.875 19.230 ;
        RECT 483.065 19.215 483.395 19.230 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.570 19.280 517.890 19.340 ;
        RECT 524.470 19.280 524.790 19.340 ;
        RECT 478.100 19.140 483.300 19.280 ;
        RECT 139.450 18.940 139.770 19.000 ;
        RECT 478.100 18.940 478.240 19.140 ;
        RECT 139.450 18.800 478.240 18.940 ;
        RECT 483.160 18.940 483.300 19.140 ;
        RECT 517.570 19.140 524.790 19.280 ;
        RECT 517.570 19.080 517.890 19.140 ;
        RECT 524.470 19.080 524.790 19.140 ;
        RECT 512.970 18.940 513.290 19.000 ;
        RECT 483.160 18.800 513.290 18.940 ;
        RECT 139.450 18.740 139.770 18.800 ;
        RECT 512.970 18.740 513.290 18.800 ;
      LAYER via ;
        RECT 139.480 18.740 139.740 19.000 ;
        RECT 517.600 19.080 517.860 19.340 ;
        RECT 524.500 19.080 524.760 19.340 ;
        RECT 513.000 18.740 513.260 19.000 ;
      LAYER met2 ;
        RECT 528.250 1600.450 528.530 1604.000 ;
        RECT 524.560 1600.310 528.530 1600.450 ;
        RECT 512.990 19.195 513.270 19.565 ;
        RECT 517.590 19.195 517.870 19.565 ;
        RECT 524.560 19.370 524.700 1600.310 ;
        RECT 528.250 1600.000 528.530 1600.310 ;
        RECT 513.060 19.030 513.200 19.195 ;
        RECT 517.600 19.050 517.860 19.195 ;
        RECT 524.500 19.050 524.760 19.370 ;
        RECT 139.480 18.710 139.740 19.030 ;
        RECT 513.000 18.710 513.260 19.030 ;
        RECT 139.540 2.400 139.680 18.710 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 512.990 19.240 513.270 19.520 ;
        RECT 517.590 19.240 517.870 19.520 ;
      LAYER met3 ;
        RECT 512.965 19.530 513.295 19.545 ;
        RECT 517.565 19.530 517.895 19.545 ;
        RECT 512.965 19.230 517.895 19.530 ;
        RECT 512.965 19.215 513.295 19.230 ;
        RECT 517.565 19.215 517.895 19.230 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 541.030 19.280 541.350 19.340 ;
        RECT 530.540 19.140 541.350 19.280 ;
        RECT 157.390 18.600 157.710 18.660 ;
        RECT 530.540 18.600 530.680 19.140 ;
        RECT 541.030 19.080 541.350 19.140 ;
        RECT 157.390 18.460 530.680 18.600 ;
        RECT 542.410 18.600 542.730 18.660 ;
        RECT 552.070 18.600 552.390 18.660 ;
        RECT 542.410 18.460 552.390 18.600 ;
        RECT 157.390 18.400 157.710 18.460 ;
        RECT 542.410 18.400 542.730 18.460 ;
        RECT 552.070 18.400 552.390 18.460 ;
      LAYER via ;
        RECT 157.420 18.400 157.680 18.660 ;
        RECT 541.060 19.080 541.320 19.340 ;
        RECT 542.440 18.400 542.700 18.660 ;
        RECT 552.100 18.400 552.360 18.660 ;
      LAYER met2 ;
        RECT 557.690 1600.450 557.970 1604.000 ;
        RECT 552.160 1600.310 557.970 1600.450 ;
        RECT 541.060 19.050 541.320 19.370 ;
        RECT 541.120 18.770 541.260 19.050 ;
        RECT 541.120 18.690 542.640 18.770 ;
        RECT 552.160 18.690 552.300 1600.310 ;
        RECT 557.690 1600.000 557.970 1600.310 ;
        RECT 157.420 18.370 157.680 18.690 ;
        RECT 541.120 18.630 542.700 18.690 ;
        RECT 542.440 18.370 542.700 18.630 ;
        RECT 552.100 18.370 552.360 18.690 ;
        RECT 157.480 2.400 157.620 18.370 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 570.010 18.260 570.330 18.320 ;
        RECT 570.010 18.120 580.820 18.260 ;
        RECT 570.010 18.060 570.330 18.120 ;
        RECT 580.680 17.920 580.820 18.120 ;
        RECT 586.570 17.920 586.890 17.980 ;
        RECT 580.680 17.780 586.890 17.920 ;
        RECT 586.570 17.720 586.890 17.780 ;
        RECT 174.870 17.580 175.190 17.640 ;
        RECT 568.170 17.580 568.490 17.640 ;
        RECT 174.870 17.440 568.490 17.580 ;
        RECT 174.870 17.380 175.190 17.440 ;
        RECT 568.170 17.380 568.490 17.440 ;
      LAYER via ;
        RECT 570.040 18.060 570.300 18.320 ;
        RECT 586.600 17.720 586.860 17.980 ;
        RECT 174.900 17.380 175.160 17.640 ;
        RECT 568.200 17.380 568.460 17.640 ;
      LAYER met2 ;
        RECT 586.670 1600.380 586.950 1604.000 ;
        RECT 586.660 1600.000 586.950 1600.380 ;
        RECT 570.040 18.090 570.300 18.350 ;
        RECT 569.180 18.030 570.300 18.090 ;
        RECT 569.180 17.950 570.240 18.030 ;
        RECT 586.660 18.010 586.800 1600.000 ;
        RECT 174.900 17.350 175.160 17.670 ;
        RECT 568.200 17.410 568.460 17.670 ;
        RECT 569.180 17.410 569.320 17.950 ;
        RECT 586.600 17.690 586.860 18.010 ;
        RECT 568.200 17.350 569.320 17.410 ;
        RECT 174.960 2.400 175.100 17.350 ;
        RECT 568.260 17.270 569.320 17.350 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.970 17.240 214.290 17.300 ;
        RECT 614.630 17.240 614.950 17.300 ;
        RECT 213.970 17.100 614.950 17.240 ;
        RECT 213.970 17.040 214.290 17.100 ;
        RECT 614.630 17.040 614.950 17.100 ;
        RECT 192.810 15.880 193.130 15.940 ;
        RECT 213.970 15.880 214.290 15.940 ;
        RECT 192.810 15.740 214.290 15.880 ;
        RECT 192.810 15.680 193.130 15.740 ;
        RECT 213.970 15.680 214.290 15.740 ;
      LAYER via ;
        RECT 214.000 17.040 214.260 17.300 ;
        RECT 614.660 17.040 614.920 17.300 ;
        RECT 192.840 15.680 193.100 15.940 ;
        RECT 214.000 15.680 214.260 15.940 ;
      LAYER met2 ;
        RECT 616.110 1600.450 616.390 1604.000 ;
        RECT 614.720 1600.310 616.390 1600.450 ;
        RECT 614.720 17.330 614.860 1600.310 ;
        RECT 616.110 1600.000 616.390 1600.310 ;
        RECT 214.000 17.010 214.260 17.330 ;
        RECT 614.660 17.010 614.920 17.330 ;
        RECT 214.060 15.970 214.200 17.010 ;
        RECT 192.840 15.650 193.100 15.970 ;
        RECT 214.000 15.650 214.260 15.970 ;
        RECT 192.900 2.400 193.040 15.650 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1592.120 213.830 1592.180 ;
        RECT 644.990 1592.120 645.310 1592.180 ;
        RECT 213.510 1591.980 645.310 1592.120 ;
        RECT 213.510 1591.920 213.830 1591.980 ;
        RECT 644.990 1591.920 645.310 1591.980 ;
        RECT 210.750 17.240 211.070 17.300 ;
        RECT 213.510 17.240 213.830 17.300 ;
        RECT 210.750 17.100 213.830 17.240 ;
        RECT 210.750 17.040 211.070 17.100 ;
        RECT 213.510 17.040 213.830 17.100 ;
      LAYER via ;
        RECT 213.540 1591.920 213.800 1592.180 ;
        RECT 645.020 1591.920 645.280 1592.180 ;
        RECT 210.780 17.040 211.040 17.300 ;
        RECT 213.540 17.040 213.800 17.300 ;
      LAYER met2 ;
        RECT 645.090 1600.380 645.370 1604.000 ;
        RECT 645.080 1600.000 645.370 1600.380 ;
        RECT 645.080 1592.210 645.220 1600.000 ;
        RECT 213.540 1591.890 213.800 1592.210 ;
        RECT 645.020 1591.890 645.280 1592.210 ;
        RECT 213.600 17.330 213.740 1591.890 ;
        RECT 210.780 17.010 211.040 17.330 ;
        RECT 213.540 17.010 213.800 17.330 ;
        RECT 210.840 2.400 210.980 17.010 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 228.690 14.520 229.010 14.580 ;
        RECT 669.830 14.520 670.150 14.580 ;
        RECT 228.690 14.380 670.150 14.520 ;
        RECT 228.690 14.320 229.010 14.380 ;
        RECT 669.830 14.320 670.150 14.380 ;
      LAYER via ;
        RECT 228.720 14.320 228.980 14.580 ;
        RECT 669.860 14.320 670.120 14.580 ;
      LAYER met2 ;
        RECT 674.530 1600.450 674.810 1604.000 ;
        RECT 669.920 1600.310 674.810 1600.450 ;
        RECT 669.920 14.610 670.060 1600.310 ;
        RECT 674.530 1600.000 674.810 1600.310 ;
        RECT 228.720 14.290 228.980 14.610 ;
        RECT 669.860 14.290 670.120 14.610 ;
        RECT 228.780 2.400 228.920 14.290 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 1592.460 55.130 1592.520 ;
        RECT 382.330 1592.460 382.650 1592.520 ;
        RECT 54.810 1592.320 382.650 1592.460 ;
        RECT 54.810 1592.260 55.130 1592.320 ;
        RECT 382.330 1592.260 382.650 1592.320 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 54.810 17.580 55.130 17.640 ;
        RECT 50.210 17.440 55.130 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 54.810 17.380 55.130 17.440 ;
      LAYER via ;
        RECT 54.840 1592.260 55.100 1592.520 ;
        RECT 382.360 1592.260 382.620 1592.520 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 54.840 17.380 55.100 17.640 ;
      LAYER met2 ;
        RECT 382.430 1600.380 382.710 1604.000 ;
        RECT 382.420 1600.000 382.710 1600.380 ;
        RECT 382.420 1592.550 382.560 1600.000 ;
        RECT 54.840 1592.230 55.100 1592.550 ;
        RECT 382.360 1592.230 382.620 1592.550 ;
        RECT 54.900 17.670 55.040 1592.230 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 54.840 17.350 55.100 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1588.040 255.230 1588.100 ;
        RECT 713.070 1588.040 713.390 1588.100 ;
        RECT 254.910 1587.900 713.390 1588.040 ;
        RECT 254.910 1587.840 255.230 1587.900 ;
        RECT 713.070 1587.840 713.390 1587.900 ;
        RECT 252.610 15.880 252.930 15.940 ;
        RECT 254.910 15.880 255.230 15.940 ;
        RECT 252.610 15.740 255.230 15.880 ;
        RECT 252.610 15.680 252.930 15.740 ;
        RECT 254.910 15.680 255.230 15.740 ;
      LAYER via ;
        RECT 254.940 1587.840 255.200 1588.100 ;
        RECT 713.100 1587.840 713.360 1588.100 ;
        RECT 252.640 15.680 252.900 15.940 ;
        RECT 254.940 15.680 255.200 15.940 ;
      LAYER met2 ;
        RECT 713.170 1600.380 713.450 1604.000 ;
        RECT 713.160 1600.000 713.450 1600.380 ;
        RECT 713.160 1588.130 713.300 1600.000 ;
        RECT 254.940 1587.810 255.200 1588.130 ;
        RECT 713.100 1587.810 713.360 1588.130 ;
        RECT 255.000 15.970 255.140 1587.810 ;
        RECT 252.640 15.650 252.900 15.970 ;
        RECT 254.940 15.650 255.200 15.970 ;
        RECT 252.700 2.400 252.840 15.650 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 270.090 15.200 270.410 15.260 ;
        RECT 738.370 15.200 738.690 15.260 ;
        RECT 270.090 15.060 738.690 15.200 ;
        RECT 270.090 15.000 270.410 15.060 ;
        RECT 738.370 15.000 738.690 15.060 ;
      LAYER via ;
        RECT 270.120 15.000 270.380 15.260 ;
        RECT 738.400 15.000 738.660 15.260 ;
      LAYER met2 ;
        RECT 742.610 1600.450 742.890 1604.000 ;
        RECT 738.460 1600.310 742.890 1600.450 ;
        RECT 738.460 15.290 738.600 1600.310 ;
        RECT 742.610 1600.000 742.890 1600.310 ;
        RECT 270.120 14.970 270.380 15.290 ;
        RECT 738.400 14.970 738.660 15.290 ;
        RECT 270.180 2.400 270.320 14.970 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 288.030 15.540 288.350 15.600 ;
        RECT 765.970 15.540 766.290 15.600 ;
        RECT 288.030 15.400 766.290 15.540 ;
        RECT 288.030 15.340 288.350 15.400 ;
        RECT 765.970 15.340 766.290 15.400 ;
      LAYER via ;
        RECT 288.060 15.340 288.320 15.600 ;
        RECT 766.000 15.340 766.260 15.600 ;
      LAYER met2 ;
        RECT 771.590 1600.450 771.870 1604.000 ;
        RECT 766.060 1600.310 771.870 1600.450 ;
        RECT 766.060 15.630 766.200 1600.310 ;
        RECT 771.590 1600.000 771.870 1600.310 ;
        RECT 288.060 15.310 288.320 15.630 ;
        RECT 766.000 15.310 766.260 15.630 ;
        RECT 288.120 2.400 288.260 15.310 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 1588.380 310.430 1588.440 ;
        RECT 800.930 1588.380 801.250 1588.440 ;
        RECT 310.110 1588.240 801.250 1588.380 ;
        RECT 310.110 1588.180 310.430 1588.240 ;
        RECT 800.930 1588.180 801.250 1588.240 ;
        RECT 305.970 16.900 306.290 16.960 ;
        RECT 310.110 16.900 310.430 16.960 ;
        RECT 305.970 16.760 310.430 16.900 ;
        RECT 305.970 16.700 306.290 16.760 ;
        RECT 310.110 16.700 310.430 16.760 ;
      LAYER via ;
        RECT 310.140 1588.180 310.400 1588.440 ;
        RECT 800.960 1588.180 801.220 1588.440 ;
        RECT 306.000 16.700 306.260 16.960 ;
        RECT 310.140 16.700 310.400 16.960 ;
      LAYER met2 ;
        RECT 801.030 1600.380 801.310 1604.000 ;
        RECT 801.020 1600.000 801.310 1600.380 ;
        RECT 801.020 1588.470 801.160 1600.000 ;
        RECT 310.140 1588.150 310.400 1588.470 ;
        RECT 800.960 1588.150 801.220 1588.470 ;
        RECT 310.200 16.990 310.340 1588.150 ;
        RECT 306.000 16.670 306.260 16.990 ;
        RECT 310.140 16.670 310.400 16.990 ;
        RECT 306.060 2.400 306.200 16.670 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 1588.720 324.230 1588.780 ;
        RECT 829.910 1588.720 830.230 1588.780 ;
        RECT 323.910 1588.580 830.230 1588.720 ;
        RECT 323.910 1588.520 324.230 1588.580 ;
        RECT 829.910 1588.520 830.230 1588.580 ;
      LAYER via ;
        RECT 323.940 1588.520 324.200 1588.780 ;
        RECT 829.940 1588.520 830.200 1588.780 ;
      LAYER met2 ;
        RECT 830.010 1600.380 830.290 1604.000 ;
        RECT 830.000 1600.000 830.290 1600.380 ;
        RECT 830.000 1588.810 830.140 1600.000 ;
        RECT 323.940 1588.490 324.200 1588.810 ;
        RECT 829.940 1588.490 830.200 1588.810 ;
        RECT 324.000 2.400 324.140 1588.490 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 341.390 16.900 341.710 16.960 ;
        RECT 341.390 16.760 376.120 16.900 ;
        RECT 341.390 16.700 341.710 16.760 ;
        RECT 375.980 16.560 376.120 16.760 ;
        RECT 855.670 16.560 855.990 16.620 ;
        RECT 375.980 16.420 855.990 16.560 ;
        RECT 855.670 16.360 855.990 16.420 ;
      LAYER via ;
        RECT 341.420 16.700 341.680 16.960 ;
        RECT 855.700 16.360 855.960 16.620 ;
      LAYER met2 ;
        RECT 859.450 1600.450 859.730 1604.000 ;
        RECT 855.760 1600.310 859.730 1600.450 ;
        RECT 341.420 16.670 341.680 16.990 ;
        RECT 341.480 2.400 341.620 16.670 ;
        RECT 855.760 16.650 855.900 1600.310 ;
        RECT 859.450 1600.000 859.730 1600.310 ;
        RECT 855.700 16.330 855.960 16.650 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 1589.400 365.170 1589.460 ;
        RECT 888.330 1589.400 888.650 1589.460 ;
        RECT 364.850 1589.260 888.650 1589.400 ;
        RECT 364.850 1589.200 365.170 1589.260 ;
        RECT 888.330 1589.200 888.650 1589.260 ;
        RECT 359.330 20.640 359.650 20.700 ;
        RECT 364.850 20.640 365.170 20.700 ;
        RECT 359.330 20.500 365.170 20.640 ;
        RECT 359.330 20.440 359.650 20.500 ;
        RECT 364.850 20.440 365.170 20.500 ;
      LAYER via ;
        RECT 364.880 1589.200 365.140 1589.460 ;
        RECT 888.360 1589.200 888.620 1589.460 ;
        RECT 359.360 20.440 359.620 20.700 ;
        RECT 364.880 20.440 365.140 20.700 ;
      LAYER met2 ;
        RECT 888.430 1600.380 888.710 1604.000 ;
        RECT 888.420 1600.000 888.710 1600.380 ;
        RECT 888.420 1589.490 888.560 1600.000 ;
        RECT 364.880 1589.170 365.140 1589.490 ;
        RECT 888.360 1589.170 888.620 1589.490 ;
        RECT 364.940 20.730 365.080 1589.170 ;
        RECT 359.360 20.410 359.620 20.730 ;
        RECT 364.880 20.410 365.140 20.730 ;
        RECT 359.420 2.400 359.560 20.410 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 917.870 1600.380 918.150 1604.000 ;
        RECT 917.860 1600.000 918.150 1600.380 ;
        RECT 917.860 18.885 918.000 1600.000 ;
        RECT 377.290 18.515 377.570 18.885 ;
        RECT 917.790 18.515 918.070 18.885 ;
        RECT 377.360 2.400 377.500 18.515 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 377.290 18.560 377.570 18.840 ;
        RECT 917.790 18.560 918.070 18.840 ;
      LAYER met3 ;
        RECT 377.265 18.850 377.595 18.865 ;
        RECT 917.765 18.850 918.095 18.865 ;
        RECT 377.265 18.550 918.095 18.850 ;
        RECT 377.265 18.535 377.595 18.550 ;
        RECT 917.765 18.535 918.095 18.550 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 1590.080 400.130 1590.140 ;
        RECT 946.750 1590.080 947.070 1590.140 ;
        RECT 399.810 1589.940 947.070 1590.080 ;
        RECT 399.810 1589.880 400.130 1589.940 ;
        RECT 946.750 1589.880 947.070 1589.940 ;
        RECT 395.210 20.300 395.530 20.360 ;
        RECT 399.810 20.300 400.130 20.360 ;
        RECT 395.210 20.160 400.130 20.300 ;
        RECT 395.210 20.100 395.530 20.160 ;
        RECT 399.810 20.100 400.130 20.160 ;
      LAYER via ;
        RECT 399.840 1589.880 400.100 1590.140 ;
        RECT 946.780 1589.880 947.040 1590.140 ;
        RECT 395.240 20.100 395.500 20.360 ;
        RECT 399.840 20.100 400.100 20.360 ;
      LAYER met2 ;
        RECT 946.850 1600.380 947.130 1604.000 ;
        RECT 946.840 1600.000 947.130 1600.380 ;
        RECT 946.840 1590.170 946.980 1600.000 ;
        RECT 399.840 1589.850 400.100 1590.170 ;
        RECT 946.780 1589.850 947.040 1590.170 ;
        RECT 399.900 20.390 400.040 1589.850 ;
        RECT 395.240 20.070 395.500 20.390 ;
        RECT 399.840 20.070 400.100 20.390 ;
        RECT 395.300 2.400 395.440 20.070 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 414.070 20.640 414.390 20.700 ;
        RECT 430.170 20.640 430.490 20.700 ;
        RECT 414.070 20.500 430.490 20.640 ;
        RECT 414.070 20.440 414.390 20.500 ;
        RECT 430.170 20.440 430.490 20.500 ;
        RECT 447.650 20.300 447.970 20.360 ;
        RECT 972.970 20.300 973.290 20.360 ;
        RECT 447.650 20.160 973.290 20.300 ;
        RECT 447.650 20.100 447.970 20.160 ;
        RECT 972.970 20.100 973.290 20.160 ;
      LAYER via ;
        RECT 414.100 20.440 414.360 20.700 ;
        RECT 430.200 20.440 430.460 20.700 ;
        RECT 447.680 20.100 447.940 20.360 ;
        RECT 973.000 20.100 973.260 20.360 ;
      LAYER met2 ;
        RECT 975.830 1600.450 976.110 1604.000 ;
        RECT 973.060 1600.310 976.110 1600.450 ;
        RECT 414.100 20.410 414.360 20.730 ;
        RECT 430.190 20.555 430.470 20.925 ;
        RECT 447.670 20.555 447.950 20.925 ;
        RECT 430.200 20.410 430.460 20.555 ;
        RECT 414.160 20.130 414.300 20.410 ;
        RECT 447.740 20.390 447.880 20.555 ;
        RECT 973.060 20.390 973.200 1600.310 ;
        RECT 975.830 1600.000 976.110 1600.310 ;
        RECT 413.240 19.990 414.300 20.130 ;
        RECT 447.680 20.070 447.940 20.390 ;
        RECT 973.000 20.070 973.260 20.390 ;
        RECT 413.240 2.400 413.380 19.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 430.190 20.600 430.470 20.880 ;
        RECT 447.670 20.600 447.950 20.880 ;
      LAYER met3 ;
        RECT 430.165 20.890 430.495 20.905 ;
        RECT 447.645 20.890 447.975 20.905 ;
        RECT 430.165 20.590 447.975 20.890 ;
        RECT 430.165 20.575 430.495 20.590 ;
        RECT 447.645 20.575 447.975 20.590 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 74.130 19.960 74.450 20.020 ;
        RECT 420.970 19.960 421.290 20.020 ;
        RECT 74.130 19.820 421.290 19.960 ;
        RECT 74.130 19.760 74.450 19.820 ;
        RECT 420.970 19.760 421.290 19.820 ;
      LAYER via ;
        RECT 74.160 19.760 74.420 20.020 ;
        RECT 421.000 19.760 421.260 20.020 ;
      LAYER met2 ;
        RECT 421.070 1600.380 421.350 1604.000 ;
        RECT 421.060 1600.000 421.350 1600.380 ;
        RECT 421.060 20.050 421.200 1600.000 ;
        RECT 74.160 19.730 74.420 20.050 ;
        RECT 421.000 19.730 421.260 20.050 ;
        RECT 74.220 2.400 74.360 19.730 ;
        RECT 74.010 -4.800 74.570 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 441.210 1593.480 441.530 1593.540 ;
        RECT 1005.170 1593.480 1005.490 1593.540 ;
        RECT 441.210 1593.340 1005.490 1593.480 ;
        RECT 441.210 1593.280 441.530 1593.340 ;
        RECT 1005.170 1593.280 1005.490 1593.340 ;
        RECT 434.310 1592.460 434.630 1592.520 ;
        RECT 441.210 1592.460 441.530 1592.520 ;
        RECT 434.310 1592.320 441.530 1592.460 ;
        RECT 434.310 1592.260 434.630 1592.320 ;
        RECT 441.210 1592.260 441.530 1592.320 ;
        RECT 434.310 1318.560 434.630 1318.820 ;
        RECT 434.400 1318.140 434.540 1318.560 ;
        RECT 434.310 1317.880 434.630 1318.140 ;
        RECT 434.310 1139.040 434.630 1139.300 ;
        RECT 434.400 1138.620 434.540 1139.040 ;
        RECT 434.310 1138.360 434.630 1138.620 ;
        RECT 434.310 904.440 434.630 904.700 ;
        RECT 434.400 904.020 434.540 904.440 ;
        RECT 434.310 903.760 434.630 904.020 ;
        RECT 434.310 849.360 434.630 849.620 ;
        RECT 434.400 848.940 434.540 849.360 ;
        RECT 434.310 848.680 434.630 848.940 ;
        RECT 430.630 28.120 430.950 28.180 ;
        RECT 434.310 28.120 434.630 28.180 ;
        RECT 430.630 27.980 434.630 28.120 ;
        RECT 430.630 27.920 430.950 27.980 ;
        RECT 434.310 27.920 434.630 27.980 ;
      LAYER via ;
        RECT 441.240 1593.280 441.500 1593.540 ;
        RECT 1005.200 1593.280 1005.460 1593.540 ;
        RECT 434.340 1592.260 434.600 1592.520 ;
        RECT 441.240 1592.260 441.500 1592.520 ;
        RECT 434.340 1318.560 434.600 1318.820 ;
        RECT 434.340 1317.880 434.600 1318.140 ;
        RECT 434.340 1139.040 434.600 1139.300 ;
        RECT 434.340 1138.360 434.600 1138.620 ;
        RECT 434.340 904.440 434.600 904.700 ;
        RECT 434.340 903.760 434.600 904.020 ;
        RECT 434.340 849.360 434.600 849.620 ;
        RECT 434.340 848.680 434.600 848.940 ;
        RECT 430.660 27.920 430.920 28.180 ;
        RECT 434.340 27.920 434.600 28.180 ;
      LAYER met2 ;
        RECT 1005.270 1600.380 1005.550 1604.000 ;
        RECT 1005.260 1600.000 1005.550 1600.380 ;
        RECT 1005.260 1593.570 1005.400 1600.000 ;
        RECT 441.240 1593.250 441.500 1593.570 ;
        RECT 1005.200 1593.250 1005.460 1593.570 ;
        RECT 441.300 1592.550 441.440 1593.250 ;
        RECT 434.340 1592.230 434.600 1592.550 ;
        RECT 441.240 1592.230 441.500 1592.550 ;
        RECT 434.400 1318.850 434.540 1592.230 ;
        RECT 434.340 1318.530 434.600 1318.850 ;
        RECT 434.340 1317.850 434.600 1318.170 ;
        RECT 434.400 1139.330 434.540 1317.850 ;
        RECT 434.340 1139.010 434.600 1139.330 ;
        RECT 434.340 1138.330 434.600 1138.650 ;
        RECT 434.400 904.730 434.540 1138.330 ;
        RECT 434.340 904.410 434.600 904.730 ;
        RECT 434.340 903.730 434.600 904.050 ;
        RECT 434.400 849.650 434.540 903.730 ;
        RECT 434.340 849.330 434.600 849.650 ;
        RECT 434.340 848.650 434.600 848.970 ;
        RECT 434.400 28.210 434.540 848.650 ;
        RECT 430.660 27.890 430.920 28.210 ;
        RECT 434.340 27.890 434.600 28.210 ;
        RECT 430.720 2.400 430.860 27.890 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 448.570 19.960 448.890 20.020 ;
        RECT 466.050 19.960 466.370 20.020 ;
        RECT 448.570 19.820 466.370 19.960 ;
        RECT 448.570 19.760 448.890 19.820 ;
        RECT 466.050 19.760 466.370 19.820 ;
        RECT 469.270 19.620 469.590 19.680 ;
        RECT 1028.170 19.620 1028.490 19.680 ;
        RECT 469.270 19.480 1028.490 19.620 ;
        RECT 469.270 19.420 469.590 19.480 ;
        RECT 1028.170 19.420 1028.490 19.480 ;
      LAYER via ;
        RECT 448.600 19.760 448.860 20.020 ;
        RECT 466.080 19.760 466.340 20.020 ;
        RECT 469.300 19.420 469.560 19.680 ;
        RECT 1028.200 19.420 1028.460 19.680 ;
      LAYER met2 ;
        RECT 1034.250 1600.450 1034.530 1604.000 ;
        RECT 1028.260 1600.310 1034.530 1600.450 ;
        RECT 448.600 19.730 448.860 20.050 ;
        RECT 466.080 19.730 466.340 20.050 ;
        RECT 448.660 2.400 448.800 19.730 ;
        RECT 466.140 19.565 466.280 19.730 ;
        RECT 1028.260 19.710 1028.400 1600.310 ;
        RECT 1034.250 1600.000 1034.530 1600.310 ;
        RECT 469.300 19.565 469.560 19.710 ;
        RECT 466.070 19.195 466.350 19.565 ;
        RECT 469.290 19.195 469.570 19.565 ;
        RECT 1028.200 19.390 1028.460 19.710 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 466.070 19.240 466.350 19.520 ;
        RECT 469.290 19.240 469.570 19.520 ;
      LAYER met3 ;
        RECT 466.045 19.530 466.375 19.545 ;
        RECT 469.265 19.530 469.595 19.545 ;
        RECT 466.045 19.230 469.595 19.530 ;
        RECT 466.045 19.215 466.375 19.230 ;
        RECT 469.265 19.215 469.595 19.230 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 472.950 1592.800 473.270 1592.860 ;
        RECT 1063.590 1592.800 1063.910 1592.860 ;
        RECT 472.950 1592.660 1063.910 1592.800 ;
        RECT 472.950 1592.600 473.270 1592.660 ;
        RECT 1063.590 1592.600 1063.910 1592.660 ;
        RECT 468.810 1591.440 469.130 1591.500 ;
        RECT 472.950 1591.440 473.270 1591.500 ;
        RECT 468.810 1591.300 473.270 1591.440 ;
        RECT 468.810 1591.240 469.130 1591.300 ;
        RECT 472.950 1591.240 473.270 1591.300 ;
      LAYER via ;
        RECT 472.980 1592.600 473.240 1592.860 ;
        RECT 1063.620 1592.600 1063.880 1592.860 ;
        RECT 468.840 1591.240 469.100 1591.500 ;
        RECT 472.980 1591.240 473.240 1591.500 ;
      LAYER met2 ;
        RECT 1063.690 1600.380 1063.970 1604.000 ;
        RECT 1063.680 1600.000 1063.970 1600.380 ;
        RECT 1063.680 1592.890 1063.820 1600.000 ;
        RECT 472.980 1592.570 473.240 1592.890 ;
        RECT 1063.620 1592.570 1063.880 1592.890 ;
        RECT 473.040 1591.530 473.180 1592.570 ;
        RECT 468.840 1591.210 469.100 1591.530 ;
        RECT 472.980 1591.210 473.240 1591.530 ;
        RECT 468.900 3.130 469.040 1591.210 ;
        RECT 466.600 2.990 469.040 3.130 ;
        RECT 466.600 2.400 466.740 2.990 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 484.450 19.280 484.770 19.340 ;
        RECT 1090.270 19.280 1090.590 19.340 ;
        RECT 484.450 19.140 513.660 19.280 ;
        RECT 484.450 19.080 484.770 19.140 ;
        RECT 513.520 18.940 513.660 19.140 ;
        RECT 541.580 19.140 1090.590 19.280 ;
        RECT 529.990 18.940 530.310 19.000 ;
        RECT 513.520 18.800 530.310 18.940 ;
        RECT 529.990 18.740 530.310 18.800 ;
        RECT 530.910 18.940 531.230 19.000 ;
        RECT 541.580 18.940 541.720 19.140 ;
        RECT 1090.270 19.080 1090.590 19.140 ;
        RECT 530.910 18.800 541.720 18.940 ;
        RECT 530.910 18.740 531.230 18.800 ;
      LAYER via ;
        RECT 484.480 19.080 484.740 19.340 ;
        RECT 530.020 18.740 530.280 19.000 ;
        RECT 530.940 18.740 531.200 19.000 ;
        RECT 1090.300 19.080 1090.560 19.340 ;
      LAYER met2 ;
        RECT 1092.670 1600.450 1092.950 1604.000 ;
        RECT 1090.360 1600.310 1092.950 1600.450 ;
        RECT 1090.360 19.370 1090.500 1600.310 ;
        RECT 1092.670 1600.000 1092.950 1600.310 ;
        RECT 484.480 19.050 484.740 19.370 ;
        RECT 1090.300 19.050 1090.560 19.370 ;
        RECT 484.540 2.400 484.680 19.050 ;
        RECT 530.020 18.940 530.280 19.030 ;
        RECT 530.940 18.940 531.200 19.030 ;
        RECT 530.020 18.800 531.200 18.940 ;
        RECT 530.020 18.710 530.280 18.800 ;
        RECT 530.940 18.710 531.200 18.800 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 538.270 1591.780 538.590 1591.840 ;
        RECT 1122.010 1591.780 1122.330 1591.840 ;
        RECT 538.270 1591.640 1122.330 1591.780 ;
        RECT 538.270 1591.580 538.590 1591.640 ;
        RECT 1122.010 1591.580 1122.330 1591.640 ;
        RECT 503.310 1590.760 503.630 1590.820 ;
        RECT 503.310 1590.620 509.980 1590.760 ;
        RECT 503.310 1590.560 503.630 1590.620 ;
        RECT 509.840 1590.420 509.980 1590.620 ;
        RECT 538.270 1590.420 538.590 1590.480 ;
        RECT 509.840 1590.280 538.590 1590.420 ;
        RECT 538.270 1590.220 538.590 1590.280 ;
      LAYER via ;
        RECT 538.300 1591.580 538.560 1591.840 ;
        RECT 1122.040 1591.580 1122.300 1591.840 ;
        RECT 503.340 1590.560 503.600 1590.820 ;
        RECT 538.300 1590.220 538.560 1590.480 ;
      LAYER met2 ;
        RECT 1122.110 1600.380 1122.390 1604.000 ;
        RECT 1122.100 1600.000 1122.390 1600.380 ;
        RECT 1122.100 1591.870 1122.240 1600.000 ;
        RECT 538.300 1591.550 538.560 1591.870 ;
        RECT 1122.040 1591.550 1122.300 1591.870 ;
        RECT 503.340 1590.530 503.600 1590.850 ;
        RECT 503.400 3.130 503.540 1590.530 ;
        RECT 538.360 1590.510 538.500 1591.550 ;
        RECT 538.300 1590.190 538.560 1590.510 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.090 1600.450 1151.370 1604.000 ;
        RECT 1145.560 1600.310 1151.370 1600.450 ;
        RECT 1145.560 16.845 1145.700 1600.310 ;
        RECT 1151.090 1600.000 1151.370 1600.310 ;
        RECT 519.890 16.475 520.170 16.845 ;
        RECT 1145.490 16.475 1145.770 16.845 ;
        RECT 519.960 2.400 520.100 16.475 ;
        RECT 519.750 -4.800 520.310 2.400 ;
      LAYER via2 ;
        RECT 519.890 16.520 520.170 16.800 ;
        RECT 1145.490 16.520 1145.770 16.800 ;
      LAYER met3 ;
        RECT 519.865 16.810 520.195 16.825 ;
        RECT 1145.465 16.810 1145.795 16.825 ;
        RECT 519.865 16.510 1145.795 16.810 ;
        RECT 519.865 16.495 520.195 16.510 ;
        RECT 1145.465 16.495 1145.795 16.510 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.350 1590.760 537.670 1590.820 ;
        RECT 1180.430 1590.760 1180.750 1590.820 ;
        RECT 537.350 1590.620 1180.750 1590.760 ;
        RECT 537.350 1590.560 537.670 1590.620 ;
        RECT 1180.430 1590.560 1180.750 1590.620 ;
      LAYER via ;
        RECT 537.380 1590.560 537.640 1590.820 ;
        RECT 1180.460 1590.560 1180.720 1590.820 ;
      LAYER met2 ;
        RECT 1180.530 1600.380 1180.810 1604.000 ;
        RECT 1180.520 1600.000 1180.810 1600.380 ;
        RECT 1180.520 1590.850 1180.660 1600.000 ;
        RECT 537.380 1590.530 537.640 1590.850 ;
        RECT 1180.460 1590.530 1180.720 1590.850 ;
        RECT 537.440 17.410 537.580 1590.530 ;
        RECT 537.440 17.270 538.040 17.410 ;
        RECT 537.900 2.400 538.040 17.270 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 555.750 18.600 556.070 18.660 ;
        RECT 1207.570 18.600 1207.890 18.660 ;
        RECT 555.750 18.460 1207.890 18.600 ;
        RECT 555.750 18.400 556.070 18.460 ;
        RECT 1207.570 18.400 1207.890 18.460 ;
      LAYER via ;
        RECT 555.780 18.400 556.040 18.660 ;
        RECT 1207.600 18.400 1207.860 18.660 ;
      LAYER met2 ;
        RECT 1209.510 1600.450 1209.790 1604.000 ;
        RECT 1207.660 1600.310 1209.790 1600.450 ;
        RECT 1207.660 18.690 1207.800 1600.310 ;
        RECT 1209.510 1600.000 1209.790 1600.310 ;
        RECT 555.780 18.370 556.040 18.690 ;
        RECT 1207.600 18.370 1207.860 18.690 ;
        RECT 555.840 2.400 555.980 18.370 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 573.690 18.940 574.010 19.000 ;
        RECT 579.210 18.940 579.530 19.000 ;
        RECT 573.690 18.800 579.530 18.940 ;
        RECT 573.690 18.740 574.010 18.800 ;
        RECT 579.210 18.740 579.530 18.800 ;
      LAYER via ;
        RECT 573.720 18.740 573.980 19.000 ;
        RECT 579.240 18.740 579.500 19.000 ;
      LAYER met2 ;
        RECT 1238.950 1600.380 1239.230 1604.000 ;
        RECT 1238.940 1600.000 1239.230 1600.380 ;
        RECT 1238.940 1591.725 1239.080 1600.000 ;
        RECT 579.230 1591.355 579.510 1591.725 ;
        RECT 1238.870 1591.355 1239.150 1591.725 ;
        RECT 579.300 19.030 579.440 1591.355 ;
        RECT 573.720 18.710 573.980 19.030 ;
        RECT 579.240 18.710 579.500 19.030 ;
        RECT 573.780 2.400 573.920 18.710 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 579.230 1591.400 579.510 1591.680 ;
        RECT 1238.870 1591.400 1239.150 1591.680 ;
      LAYER met3 ;
        RECT 579.205 1591.690 579.535 1591.705 ;
        RECT 1238.845 1591.690 1239.175 1591.705 ;
        RECT 579.205 1591.390 1239.175 1591.690 ;
        RECT 579.205 1591.375 579.535 1591.390 ;
        RECT 1238.845 1591.375 1239.175 1591.390 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 614.170 18.260 614.490 18.320 ;
        RECT 1262.770 18.260 1263.090 18.320 ;
        RECT 614.170 18.120 1263.090 18.260 ;
        RECT 614.170 18.060 614.490 18.120 ;
        RECT 1262.770 18.060 1263.090 18.120 ;
        RECT 591.170 17.920 591.490 17.980 ;
        RECT 591.170 17.780 602.440 17.920 ;
        RECT 591.170 17.720 591.490 17.780 ;
        RECT 602.300 17.580 602.440 17.780 ;
        RECT 613.250 17.580 613.570 17.640 ;
        RECT 602.300 17.440 613.570 17.580 ;
        RECT 613.250 17.380 613.570 17.440 ;
      LAYER via ;
        RECT 614.200 18.060 614.460 18.320 ;
        RECT 1262.800 18.060 1263.060 18.320 ;
        RECT 591.200 17.720 591.460 17.980 ;
        RECT 613.280 17.380 613.540 17.640 ;
      LAYER met2 ;
        RECT 1267.930 1600.450 1268.210 1604.000 ;
        RECT 1262.860 1600.310 1268.210 1600.450 ;
        RECT 1262.860 18.350 1263.000 1600.310 ;
        RECT 1267.930 1600.000 1268.210 1600.310 ;
        RECT 614.200 18.030 614.460 18.350 ;
        RECT 1262.800 18.030 1263.060 18.350 ;
        RECT 591.200 17.690 591.460 18.010 ;
        RECT 591.260 2.400 591.400 17.690 ;
        RECT 613.280 17.410 613.540 17.670 ;
        RECT 614.260 17.410 614.400 18.030 ;
        RECT 613.280 17.350 614.400 17.410 ;
        RECT 613.340 17.270 614.400 17.350 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 1591.440 103.430 1591.500 ;
        RECT 460.070 1591.440 460.390 1591.500 ;
        RECT 103.110 1591.300 460.390 1591.440 ;
        RECT 103.110 1591.240 103.430 1591.300 ;
        RECT 460.070 1591.240 460.390 1591.300 ;
        RECT 97.590 17.580 97.910 17.640 ;
        RECT 103.110 17.580 103.430 17.640 ;
        RECT 97.590 17.440 103.430 17.580 ;
        RECT 97.590 17.380 97.910 17.440 ;
        RECT 103.110 17.380 103.430 17.440 ;
      LAYER via ;
        RECT 103.140 1591.240 103.400 1591.500 ;
        RECT 460.100 1591.240 460.360 1591.500 ;
        RECT 97.620 17.380 97.880 17.640 ;
        RECT 103.140 17.380 103.400 17.640 ;
      LAYER met2 ;
        RECT 460.170 1600.380 460.450 1604.000 ;
        RECT 460.160 1600.000 460.450 1600.380 ;
        RECT 460.160 1591.530 460.300 1600.000 ;
        RECT 103.140 1591.210 103.400 1591.530 ;
        RECT 460.100 1591.210 460.360 1591.530 ;
        RECT 103.200 17.670 103.340 1591.210 ;
        RECT 97.620 17.350 97.880 17.670 ;
        RECT 103.140 17.350 103.400 17.670 ;
        RECT 97.680 2.400 97.820 17.350 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 609.110 18.260 609.430 18.320 ;
        RECT 613.710 18.260 614.030 18.320 ;
        RECT 609.110 18.120 614.030 18.260 ;
        RECT 609.110 18.060 609.430 18.120 ;
        RECT 613.710 18.060 614.030 18.120 ;
      LAYER via ;
        RECT 609.140 18.060 609.400 18.320 ;
        RECT 613.740 18.060 614.000 18.320 ;
      LAYER met2 ;
        RECT 1297.370 1600.380 1297.650 1604.000 ;
        RECT 1297.360 1600.000 1297.650 1600.380 ;
        RECT 1297.360 1590.365 1297.500 1600.000 ;
        RECT 613.730 1589.995 614.010 1590.365 ;
        RECT 1297.290 1589.995 1297.570 1590.365 ;
        RECT 613.800 18.350 613.940 1589.995 ;
        RECT 609.140 18.030 609.400 18.350 ;
        RECT 613.740 18.030 614.000 18.350 ;
        RECT 609.200 2.400 609.340 18.030 ;
        RECT 608.990 -4.800 609.550 2.400 ;
      LAYER via2 ;
        RECT 613.730 1590.040 614.010 1590.320 ;
        RECT 1297.290 1590.040 1297.570 1590.320 ;
      LAYER met3 ;
        RECT 613.705 1590.330 614.035 1590.345 ;
        RECT 1297.265 1590.330 1297.595 1590.345 ;
        RECT 613.705 1590.030 1297.595 1590.330 ;
        RECT 613.705 1590.015 614.035 1590.030 ;
        RECT 1297.265 1590.015 1297.595 1590.030 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.050 17.240 627.370 17.300 ;
        RECT 1324.870 17.240 1325.190 17.300 ;
        RECT 627.050 17.100 1325.190 17.240 ;
        RECT 627.050 17.040 627.370 17.100 ;
        RECT 1324.870 17.040 1325.190 17.100 ;
      LAYER via ;
        RECT 627.080 17.040 627.340 17.300 ;
        RECT 1324.900 17.040 1325.160 17.300 ;
      LAYER met2 ;
        RECT 1326.350 1600.450 1326.630 1604.000 ;
        RECT 1324.960 1600.310 1326.630 1600.450 ;
        RECT 1324.960 17.330 1325.100 1600.310 ;
        RECT 1326.350 1600.000 1326.630 1600.310 ;
        RECT 627.080 17.010 627.340 17.330 ;
        RECT 1324.900 17.010 1325.160 17.330 ;
        RECT 627.140 2.400 627.280 17.010 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 1590.760 124.130 1590.820 ;
        RECT 499.170 1590.760 499.490 1590.820 ;
        RECT 123.810 1590.620 499.490 1590.760 ;
        RECT 123.810 1590.560 124.130 1590.620 ;
        RECT 499.170 1590.560 499.490 1590.620 ;
        RECT 121.510 17.580 121.830 17.640 ;
        RECT 123.810 17.580 124.130 17.640 ;
        RECT 121.510 17.440 124.130 17.580 ;
        RECT 121.510 17.380 121.830 17.440 ;
        RECT 123.810 17.380 124.130 17.440 ;
      LAYER via ;
        RECT 123.840 1590.560 124.100 1590.820 ;
        RECT 499.200 1590.560 499.460 1590.820 ;
        RECT 121.540 17.380 121.800 17.640 ;
        RECT 123.840 17.380 124.100 17.640 ;
      LAYER met2 ;
        RECT 499.270 1600.380 499.550 1604.000 ;
        RECT 499.260 1600.000 499.550 1600.380 ;
        RECT 499.260 1590.850 499.400 1600.000 ;
        RECT 123.840 1590.530 124.100 1590.850 ;
        RECT 499.200 1590.530 499.460 1590.850 ;
        RECT 123.900 17.670 124.040 1590.530 ;
        RECT 121.540 17.350 121.800 17.670 ;
        RECT 123.840 17.350 124.100 17.670 ;
        RECT 121.600 2.400 121.740 17.350 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 375.980 1593.000 424.420 1593.140 ;
        RECT 227.310 1592.800 227.630 1592.860 ;
        RECT 276.070 1592.800 276.390 1592.860 ;
        RECT 227.310 1592.660 276.390 1592.800 ;
        RECT 227.310 1592.600 227.630 1592.660 ;
        RECT 276.070 1592.600 276.390 1592.660 ;
        RECT 323.910 1592.800 324.230 1592.860 ;
        RECT 375.980 1592.800 376.120 1593.000 ;
        RECT 323.910 1592.660 376.120 1592.800 ;
        RECT 424.280 1592.800 424.420 1593.000 ;
        RECT 472.030 1592.800 472.350 1592.860 ;
        RECT 424.280 1592.660 472.350 1592.800 ;
        RECT 323.910 1592.600 324.230 1592.660 ;
        RECT 472.030 1592.600 472.350 1592.660 ;
        RECT 472.030 1591.780 472.350 1591.840 ;
        RECT 537.810 1591.780 538.130 1591.840 ;
        RECT 472.030 1591.640 538.130 1591.780 ;
        RECT 472.030 1591.580 472.350 1591.640 ;
        RECT 537.810 1591.580 538.130 1591.640 ;
        RECT 323.910 1589.200 324.230 1589.460 ;
        RECT 210.290 1589.060 210.610 1589.120 ;
        RECT 227.310 1589.060 227.630 1589.120 ;
        RECT 210.290 1588.920 227.630 1589.060 ;
        RECT 210.290 1588.860 210.610 1588.920 ;
        RECT 227.310 1588.860 227.630 1588.920 ;
        RECT 276.070 1589.060 276.390 1589.120 ;
        RECT 324.000 1589.060 324.140 1589.200 ;
        RECT 276.070 1588.920 324.140 1589.060 ;
        RECT 276.070 1588.860 276.390 1588.920 ;
        RECT 145.430 15.200 145.750 15.260 ;
        RECT 145.430 15.060 187.520 15.200 ;
        RECT 145.430 15.000 145.750 15.060 ;
        RECT 187.380 14.520 187.520 15.060 ;
        RECT 210.290 14.520 210.610 14.580 ;
        RECT 187.380 14.380 210.610 14.520 ;
        RECT 210.290 14.320 210.610 14.380 ;
      LAYER via ;
        RECT 227.340 1592.600 227.600 1592.860 ;
        RECT 276.100 1592.600 276.360 1592.860 ;
        RECT 323.940 1592.600 324.200 1592.860 ;
        RECT 472.060 1592.600 472.320 1592.860 ;
        RECT 472.060 1591.580 472.320 1591.840 ;
        RECT 537.840 1591.580 538.100 1591.840 ;
        RECT 323.940 1589.200 324.200 1589.460 ;
        RECT 210.320 1588.860 210.580 1589.120 ;
        RECT 227.340 1588.860 227.600 1589.120 ;
        RECT 276.100 1588.860 276.360 1589.120 ;
        RECT 145.460 15.000 145.720 15.260 ;
        RECT 210.320 14.320 210.580 14.580 ;
      LAYER met2 ;
        RECT 537.910 1600.380 538.190 1604.000 ;
        RECT 537.900 1600.000 538.190 1600.380 ;
        RECT 227.340 1592.570 227.600 1592.890 ;
        RECT 276.100 1592.570 276.360 1592.890 ;
        RECT 323.940 1592.570 324.200 1592.890 ;
        RECT 472.060 1592.570 472.320 1592.890 ;
        RECT 227.400 1589.150 227.540 1592.570 ;
        RECT 276.160 1589.150 276.300 1592.570 ;
        RECT 324.000 1589.490 324.140 1592.570 ;
        RECT 472.120 1591.870 472.260 1592.570 ;
        RECT 537.900 1591.870 538.040 1600.000 ;
        RECT 472.060 1591.550 472.320 1591.870 ;
        RECT 537.840 1591.550 538.100 1591.870 ;
        RECT 323.940 1589.170 324.200 1589.490 ;
        RECT 210.320 1588.830 210.580 1589.150 ;
        RECT 227.340 1588.830 227.600 1589.150 ;
        RECT 276.100 1588.830 276.360 1589.150 ;
        RECT 145.460 14.970 145.720 15.290 ;
        RECT 145.520 2.400 145.660 14.970 ;
        RECT 210.380 14.610 210.520 1588.830 ;
        RECT 210.320 14.290 210.580 14.610 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 565.870 18.940 566.190 19.000 ;
        RECT 542.040 18.800 566.190 18.940 ;
        RECT 531.370 18.600 531.690 18.660 ;
        RECT 542.040 18.600 542.180 18.800 ;
        RECT 565.870 18.740 566.190 18.800 ;
        RECT 531.370 18.460 542.180 18.600 ;
        RECT 531.370 18.400 531.690 18.460 ;
        RECT 163.370 17.920 163.690 17.980 ;
        RECT 531.370 17.920 531.690 17.980 ;
        RECT 163.370 17.780 531.690 17.920 ;
        RECT 163.370 17.720 163.690 17.780 ;
        RECT 531.370 17.720 531.690 17.780 ;
      LAYER via ;
        RECT 531.400 18.400 531.660 18.660 ;
        RECT 565.900 18.740 566.160 19.000 ;
        RECT 163.400 17.720 163.660 17.980 ;
        RECT 531.400 17.720 531.660 17.980 ;
      LAYER met2 ;
        RECT 567.350 1600.450 567.630 1604.000 ;
        RECT 565.960 1600.310 567.630 1600.450 ;
        RECT 565.960 19.030 566.100 1600.310 ;
        RECT 567.350 1600.000 567.630 1600.310 ;
        RECT 565.900 18.710 566.160 19.030 ;
        RECT 531.400 18.370 531.660 18.690 ;
        RECT 531.460 18.010 531.600 18.370 ;
        RECT 163.400 17.690 163.660 18.010 ;
        RECT 531.400 17.690 531.660 18.010 ;
        RECT 163.460 2.400 163.600 17.690 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 180.850 18.260 181.170 18.320 ;
        RECT 180.850 18.120 569.320 18.260 ;
        RECT 180.850 18.060 181.170 18.120 ;
        RECT 569.180 17.580 569.320 18.120 ;
        RECT 593.470 17.580 593.790 17.640 ;
        RECT 569.180 17.440 593.790 17.580 ;
        RECT 593.470 17.380 593.790 17.440 ;
      LAYER via ;
        RECT 180.880 18.060 181.140 18.320 ;
        RECT 593.500 17.380 593.760 17.640 ;
      LAYER met2 ;
        RECT 596.330 1600.450 596.610 1604.000 ;
        RECT 593.560 1600.310 596.610 1600.450 ;
        RECT 180.880 18.030 181.140 18.350 ;
        RECT 180.940 2.400 181.080 18.030 ;
        RECT 593.560 17.670 593.700 1600.310 ;
        RECT 596.330 1600.000 596.610 1600.310 ;
        RECT 593.500 17.350 593.760 17.670 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 1587.360 200.030 1587.420 ;
        RECT 623.830 1587.360 624.150 1587.420 ;
        RECT 199.710 1587.220 624.150 1587.360 ;
        RECT 199.710 1587.160 200.030 1587.220 ;
        RECT 623.830 1587.160 624.150 1587.220 ;
      LAYER via ;
        RECT 199.740 1587.160 200.000 1587.420 ;
        RECT 623.860 1587.160 624.120 1587.420 ;
      LAYER met2 ;
        RECT 625.770 1600.450 626.050 1604.000 ;
        RECT 623.920 1600.310 626.050 1600.450 ;
        RECT 623.920 1587.450 624.060 1600.310 ;
        RECT 625.770 1600.000 626.050 1600.310 ;
        RECT 199.740 1587.130 200.000 1587.450 ;
        RECT 623.860 1587.130 624.120 1587.450 ;
        RECT 199.800 16.730 199.940 1587.130 ;
        RECT 198.880 16.590 199.940 16.730 ;
        RECT 198.880 2.400 199.020 16.590 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 216.730 14.180 217.050 14.240 ;
        RECT 649.130 14.180 649.450 14.240 ;
        RECT 216.730 14.040 620.840 14.180 ;
        RECT 216.730 13.980 217.050 14.040 ;
        RECT 620.700 13.840 620.840 14.040 ;
        RECT 639.100 14.040 649.450 14.180 ;
        RECT 639.100 13.840 639.240 14.040 ;
        RECT 649.130 13.980 649.450 14.040 ;
        RECT 620.700 13.700 639.240 13.840 ;
      LAYER via ;
        RECT 216.760 13.980 217.020 14.240 ;
        RECT 649.160 13.980 649.420 14.240 ;
      LAYER met2 ;
        RECT 654.750 1600.450 655.030 1604.000 ;
        RECT 649.220 1600.310 655.030 1600.450 ;
        RECT 649.220 14.270 649.360 1600.310 ;
        RECT 654.750 1600.000 655.030 1600.310 ;
        RECT 216.760 13.950 217.020 14.270 ;
        RECT 649.160 13.950 649.420 14.270 ;
        RECT 216.820 2.400 216.960 13.950 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 1587.700 240.970 1587.760 ;
        RECT 684.090 1587.700 684.410 1587.760 ;
        RECT 240.650 1587.560 684.410 1587.700 ;
        RECT 240.650 1587.500 240.970 1587.560 ;
        RECT 684.090 1587.500 684.410 1587.560 ;
        RECT 234.670 15.880 234.990 15.940 ;
        RECT 240.650 15.880 240.970 15.940 ;
        RECT 234.670 15.740 240.970 15.880 ;
        RECT 234.670 15.680 234.990 15.740 ;
        RECT 240.650 15.680 240.970 15.740 ;
      LAYER via ;
        RECT 240.680 1587.500 240.940 1587.760 ;
        RECT 684.120 1587.500 684.380 1587.760 ;
        RECT 234.700 15.680 234.960 15.940 ;
        RECT 240.680 15.680 240.940 15.940 ;
      LAYER met2 ;
        RECT 684.190 1600.380 684.470 1604.000 ;
        RECT 684.180 1600.000 684.470 1600.380 ;
        RECT 684.180 1587.790 684.320 1600.000 ;
        RECT 240.680 1587.470 240.940 1587.790 ;
        RECT 684.120 1587.470 684.380 1587.790 ;
        RECT 240.740 15.970 240.880 1587.470 ;
        RECT 234.700 15.650 234.960 15.970 ;
        RECT 240.680 15.650 240.940 15.970 ;
        RECT 234.760 2.400 234.900 15.650 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 161.990 1590.080 162.310 1590.140 ;
        RECT 391.990 1590.080 392.310 1590.140 ;
        RECT 161.990 1589.940 392.310 1590.080 ;
        RECT 161.990 1589.880 162.310 1589.940 ;
        RECT 391.990 1589.880 392.310 1589.940 ;
        RECT 56.190 17.240 56.510 17.300 ;
        RECT 161.990 17.240 162.310 17.300 ;
        RECT 56.190 17.100 162.310 17.240 ;
        RECT 56.190 17.040 56.510 17.100 ;
        RECT 161.990 17.040 162.310 17.100 ;
      LAYER via ;
        RECT 162.020 1589.880 162.280 1590.140 ;
        RECT 392.020 1589.880 392.280 1590.140 ;
        RECT 56.220 17.040 56.480 17.300 ;
        RECT 162.020 17.040 162.280 17.300 ;
      LAYER met2 ;
        RECT 392.090 1600.380 392.370 1604.000 ;
        RECT 392.080 1600.000 392.370 1600.380 ;
        RECT 392.080 1590.170 392.220 1600.000 ;
        RECT 162.020 1589.850 162.280 1590.170 ;
        RECT 392.020 1589.850 392.280 1590.170 ;
        RECT 162.080 17.330 162.220 1589.850 ;
        RECT 56.220 17.010 56.480 17.330 ;
        RECT 162.020 17.010 162.280 17.330 ;
        RECT 56.280 2.400 56.420 17.010 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 1591.780 82.730 1591.840 ;
        RECT 431.090 1591.780 431.410 1591.840 ;
        RECT 82.410 1591.640 431.410 1591.780 ;
        RECT 82.410 1591.580 82.730 1591.640 ;
        RECT 431.090 1591.580 431.410 1591.640 ;
        RECT 80.110 17.580 80.430 17.640 ;
        RECT 82.410 17.580 82.730 17.640 ;
        RECT 80.110 17.440 82.730 17.580 ;
        RECT 80.110 17.380 80.430 17.440 ;
        RECT 82.410 17.380 82.730 17.440 ;
      LAYER via ;
        RECT 82.440 1591.580 82.700 1591.840 ;
        RECT 431.120 1591.580 431.380 1591.840 ;
        RECT 80.140 17.380 80.400 17.640 ;
        RECT 82.440 17.380 82.700 17.640 ;
      LAYER met2 ;
        RECT 431.190 1600.380 431.470 1604.000 ;
        RECT 431.180 1600.000 431.470 1600.380 ;
        RECT 431.180 1591.870 431.320 1600.000 ;
        RECT 82.440 1591.550 82.700 1591.870 ;
        RECT 431.120 1591.550 431.380 1591.870 ;
        RECT 82.500 17.670 82.640 1591.550 ;
        RECT 80.140 17.350 80.400 17.670 ;
        RECT 82.440 17.350 82.700 17.670 ;
        RECT 80.200 2.400 80.340 17.350 ;
        RECT 79.990 -4.800 80.550 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 1591.100 109.870 1591.160 ;
        RECT 469.730 1591.100 470.050 1591.160 ;
        RECT 109.550 1590.960 470.050 1591.100 ;
        RECT 109.550 1590.900 109.870 1590.960 ;
        RECT 469.730 1590.900 470.050 1590.960 ;
        RECT 103.570 17.580 103.890 17.640 ;
        RECT 109.550 17.580 109.870 17.640 ;
        RECT 103.570 17.440 109.870 17.580 ;
        RECT 103.570 17.380 103.890 17.440 ;
        RECT 109.550 17.380 109.870 17.440 ;
      LAYER via ;
        RECT 109.580 1590.900 109.840 1591.160 ;
        RECT 469.760 1590.900 470.020 1591.160 ;
        RECT 103.600 17.380 103.860 17.640 ;
        RECT 109.580 17.380 109.840 17.640 ;
      LAYER met2 ;
        RECT 469.830 1600.380 470.110 1604.000 ;
        RECT 469.820 1600.000 470.110 1600.380 ;
        RECT 469.820 1591.190 469.960 1600.000 ;
        RECT 109.580 1590.870 109.840 1591.190 ;
        RECT 469.760 1590.870 470.020 1591.190 ;
        RECT 109.640 17.670 109.780 1590.870 ;
        RECT 103.600 17.350 103.860 17.670 ;
        RECT 109.580 17.350 109.840 17.670 ;
        RECT 103.660 2.400 103.800 17.350 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 130.710 1590.420 131.030 1590.480 ;
        RECT 508.830 1590.420 509.150 1590.480 ;
        RECT 130.710 1590.280 509.150 1590.420 ;
        RECT 130.710 1590.220 131.030 1590.280 ;
        RECT 508.830 1590.220 509.150 1590.280 ;
        RECT 127.490 17.580 127.810 17.640 ;
        RECT 130.710 17.580 131.030 17.640 ;
        RECT 127.490 17.440 131.030 17.580 ;
        RECT 127.490 17.380 127.810 17.440 ;
        RECT 130.710 17.380 131.030 17.440 ;
      LAYER via ;
        RECT 130.740 1590.220 131.000 1590.480 ;
        RECT 508.860 1590.220 509.120 1590.480 ;
        RECT 127.520 17.380 127.780 17.640 ;
        RECT 130.740 17.380 131.000 17.640 ;
      LAYER met2 ;
        RECT 508.930 1600.380 509.210 1604.000 ;
        RECT 508.920 1600.000 509.210 1600.380 ;
        RECT 508.920 1590.510 509.060 1600.000 ;
        RECT 130.740 1590.190 131.000 1590.510 ;
        RECT 508.860 1590.190 509.120 1590.510 ;
        RECT 130.800 17.670 130.940 1590.190 ;
        RECT 127.520 17.350 127.780 17.670 ;
        RECT 130.740 17.350 131.000 17.670 ;
        RECT 127.580 2.400 127.720 17.350 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 196.490 1589.740 196.810 1589.800 ;
        RECT 343.230 1589.740 343.550 1589.800 ;
        RECT 196.490 1589.600 343.550 1589.740 ;
        RECT 196.490 1589.540 196.810 1589.600 ;
        RECT 343.230 1589.540 343.550 1589.600 ;
        RECT 26.290 15.880 26.610 15.940 ;
        RECT 26.290 15.740 188.900 15.880 ;
        RECT 26.290 15.680 26.610 15.740 ;
        RECT 188.760 15.540 188.900 15.740 ;
        RECT 196.490 15.540 196.810 15.600 ;
        RECT 188.760 15.400 196.810 15.540 ;
        RECT 196.490 15.340 196.810 15.400 ;
      LAYER via ;
        RECT 196.520 1589.540 196.780 1589.800 ;
        RECT 343.260 1589.540 343.520 1589.800 ;
        RECT 26.320 15.680 26.580 15.940 ;
        RECT 196.520 15.340 196.780 15.600 ;
      LAYER met2 ;
        RECT 343.330 1600.380 343.610 1604.000 ;
        RECT 343.320 1600.000 343.610 1600.380 ;
        RECT 343.320 1589.830 343.460 1600.000 ;
        RECT 196.520 1589.510 196.780 1589.830 ;
        RECT 343.260 1589.510 343.520 1589.830 ;
        RECT 26.320 15.650 26.580 15.970 ;
        RECT 26.380 2.400 26.520 15.650 ;
        RECT 196.580 15.630 196.720 1589.510 ;
        RECT 196.520 15.310 196.780 15.630 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 16.900 32.590 16.960 ;
        RECT 32.270 16.760 305.740 16.900 ;
        RECT 32.270 16.700 32.590 16.760 ;
        RECT 305.600 16.560 305.740 16.760 ;
        RECT 351.970 16.560 352.290 16.620 ;
        RECT 305.600 16.420 352.290 16.560 ;
        RECT 351.970 16.360 352.290 16.420 ;
      LAYER via ;
        RECT 32.300 16.700 32.560 16.960 ;
        RECT 352.000 16.360 352.260 16.620 ;
      LAYER met2 ;
        RECT 352.990 1600.450 353.270 1604.000 ;
        RECT 352.060 1600.310 353.270 1600.450 ;
        RECT 32.300 16.670 32.560 16.990 ;
        RECT 32.360 2.400 32.500 16.670 ;
        RECT 352.060 16.650 352.200 1600.310 ;
        RECT 352.990 1600.000 353.270 1600.310 ;
        RECT 352.000 16.330 352.260 16.650 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.480 3243.600 684.050 3244.660 ;
        RECT 1331.480 3243.600 1334.050 3244.660 ;
        RECT 1931.480 3243.600 1934.050 3244.660 ;
        RECT 1702.430 1611.575 1705.000 1612.635 ;
      LAYER via3 ;
        RECT 682.500 3243.620 684.020 3244.630 ;
        RECT 1332.500 3243.620 1334.020 3244.630 ;
        RECT 1932.500 3243.620 1934.020 3244.630 ;
        RECT 1702.460 1611.605 1703.980 1612.615 ;
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 364.020 3271.235 367.020 3529.000 ;
        RECT 382.020 3271.235 385.020 3538.400 ;
        RECT 400.020 3271.235 403.020 3547.800 ;
        RECT 418.020 3271.235 421.020 3557.200 ;
        RECT 544.020 3271.235 547.020 3529.000 ;
        RECT 562.020 3271.235 565.020 3538.400 ;
        RECT 580.020 3271.235 583.020 3547.800 ;
        RECT 598.020 3271.235 601.020 3557.200 ;
        RECT 682.470 2803.670 684.070 3244.680 ;
        RECT 382.020 2715.000 385.020 2785.000 ;
        RECT 400.020 2715.000 403.020 2785.000 ;
        RECT 418.020 2715.000 421.020 2785.000 ;
        RECT 562.020 2715.000 565.020 2785.000 ;
        RECT 580.020 2715.000 583.020 2785.000 ;
        RECT 598.020 2715.000 601.020 2785.000 ;
        RECT 724.020 2715.000 727.020 3529.000 ;
        RECT 742.020 2715.000 745.020 3538.400 ;
        RECT 760.020 2715.000 763.020 3547.800 ;
        RECT 778.020 2715.000 781.020 3557.200 ;
        RECT 904.020 2715.000 907.020 3529.000 ;
        RECT 922.020 2715.000 925.020 3538.400 ;
        RECT 940.020 3271.235 943.020 3547.800 ;
        RECT 958.020 3271.235 961.020 3557.200 ;
        RECT 1084.020 3271.235 1087.020 3529.000 ;
        RECT 1102.020 3271.235 1105.020 3538.400 ;
        RECT 1120.020 3271.235 1123.020 3547.800 ;
        RECT 1138.020 3271.235 1141.020 3557.200 ;
        RECT 1264.020 3271.235 1267.020 3529.000 ;
        RECT 1282.020 3271.235 1285.020 3538.400 ;
        RECT 1300.020 3271.235 1303.020 3547.800 ;
        RECT 1318.020 3271.235 1321.020 3557.200 ;
        RECT 1332.470 2803.670 1334.070 3244.680 ;
        RECT 940.020 2715.000 943.020 2785.000 ;
        RECT 958.020 2715.000 961.020 2785.000 ;
        RECT 1102.020 2715.000 1105.020 2785.000 ;
        RECT 1120.020 2715.000 1123.020 2785.000 ;
        RECT 1138.020 2715.000 1141.020 2785.000 ;
        RECT 1282.020 2715.000 1285.020 2785.000 ;
        RECT 1300.020 2715.000 1303.020 2785.000 ;
        RECT 1318.020 2715.000 1321.020 2785.000 ;
        RECT 321.040 1610.640 322.640 2688.240 ;
        RECT 364.020 -9.320 367.020 1585.000 ;
        RECT 382.020 -18.720 385.020 1585.000 ;
        RECT 400.020 -28.120 403.020 1585.000 ;
        RECT 418.020 -37.520 421.020 1585.000 ;
        RECT 544.020 -9.320 547.020 1585.000 ;
        RECT 562.020 -18.720 565.020 1585.000 ;
        RECT 580.020 -28.120 583.020 1585.000 ;
        RECT 598.020 -37.520 601.020 1585.000 ;
        RECT 724.020 -9.320 727.020 1585.000 ;
        RECT 742.020 -18.720 745.020 1585.000 ;
        RECT 760.020 -28.120 763.020 1585.000 ;
        RECT 778.020 -37.520 781.020 1585.000 ;
        RECT 904.020 -9.320 907.020 1585.000 ;
        RECT 922.020 -18.720 925.020 1585.000 ;
        RECT 940.020 -28.120 943.020 1585.000 ;
        RECT 958.020 -37.520 961.020 1585.000 ;
        RECT 1084.020 -9.320 1087.020 1585.000 ;
        RECT 1102.020 -18.720 1105.020 1585.000 ;
        RECT 1120.020 -28.120 1123.020 1585.000 ;
        RECT 1138.020 -37.520 1141.020 1585.000 ;
        RECT 1264.020 -9.320 1267.020 1585.000 ;
        RECT 1282.020 -18.720 1285.020 1585.000 ;
        RECT 1300.020 -28.120 1303.020 1585.000 ;
        RECT 1318.020 -37.520 1321.020 1585.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1624.020 3271.235 1627.020 3529.000 ;
        RECT 1642.020 3271.235 1645.020 3538.400 ;
        RECT 1660.020 3271.235 1663.020 3547.800 ;
        RECT 1678.020 3271.235 1681.020 3557.200 ;
        RECT 1804.020 3271.235 1807.020 3529.000 ;
        RECT 1822.020 3271.235 1825.020 3538.400 ;
        RECT 1840.020 3271.235 1843.020 3547.800 ;
        RECT 1858.020 3271.235 1861.020 3557.200 ;
        RECT 1932.470 2803.670 1934.070 3244.680 ;
        RECT 1624.020 -9.320 1627.020 2785.000 ;
        RECT 1642.020 -18.720 1645.020 2785.000 ;
        RECT 1660.020 -28.120 1663.020 2785.000 ;
        RECT 1678.020 -37.520 1681.020 2785.000 ;
        RECT 1804.020 2071.235 1807.020 2785.000 ;
        RECT 1822.020 2071.235 1825.020 2785.000 ;
        RECT 1840.020 2071.235 1843.020 2785.000 ;
        RECT 1858.020 2071.235 1861.020 2785.000 ;
        RECT 1984.020 2071.235 1987.020 3529.000 ;
        RECT 2002.020 2071.235 2005.020 3538.400 ;
        RECT 2020.020 2071.235 2023.020 3547.800 ;
        RECT 2038.020 2071.235 2041.020 3557.200 ;
        RECT 1702.410 1611.555 1704.010 2052.565 ;
        RECT 1804.020 -9.320 1807.020 1585.000 ;
        RECT 1822.020 -18.720 1825.020 1585.000 ;
        RECT 1840.020 -28.120 1843.020 1585.000 ;
        RECT 1858.020 -37.520 1861.020 1585.000 ;
        RECT 1984.020 -9.320 1987.020 1585.000 ;
        RECT 2002.020 -18.720 2005.020 1585.000 ;
        RECT 2020.020 -28.120 2023.020 1585.000 ;
        RECT 2038.020 -37.520 2041.020 1585.000 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2344.020 -9.320 2347.020 3529.000 ;
        RECT 2362.020 -18.720 2365.020 3538.400 ;
        RECT 2380.020 -28.120 2383.020 3547.800 ;
        RECT 2398.020 -37.520 2401.020 3557.200 ;
        RECT 2524.020 -9.320 2527.020 3529.000 ;
        RECT 2542.020 -18.720 2545.020 3538.400 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 682.680 3125.090 683.860 3126.270 ;
        RECT 682.680 3123.490 683.860 3124.670 ;
        RECT 682.680 3107.090 683.860 3108.270 ;
        RECT 682.680 3105.490 683.860 3106.670 ;
        RECT 682.680 3089.090 683.860 3090.270 ;
        RECT 682.680 3087.490 683.860 3088.670 ;
        RECT 682.680 3071.090 683.860 3072.270 ;
        RECT 682.680 3069.490 683.860 3070.670 ;
        RECT 682.680 2945.090 683.860 2946.270 ;
        RECT 682.680 2943.490 683.860 2944.670 ;
        RECT 682.680 2927.090 683.860 2928.270 ;
        RECT 682.680 2925.490 683.860 2926.670 ;
        RECT 682.680 2909.090 683.860 2910.270 ;
        RECT 682.680 2907.490 683.860 2908.670 ;
        RECT 682.680 2891.090 683.860 2892.270 ;
        RECT 682.680 2889.490 683.860 2890.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 1332.680 3125.090 1333.860 3126.270 ;
        RECT 1332.680 3123.490 1333.860 3124.670 ;
        RECT 1332.680 3107.090 1333.860 3108.270 ;
        RECT 1332.680 3105.490 1333.860 3106.670 ;
        RECT 1332.680 3089.090 1333.860 3090.270 ;
        RECT 1332.680 3087.490 1333.860 3088.670 ;
        RECT 1332.680 3071.090 1333.860 3072.270 ;
        RECT 1332.680 3069.490 1333.860 3070.670 ;
        RECT 1332.680 2945.090 1333.860 2946.270 ;
        RECT 1332.680 2943.490 1333.860 2944.670 ;
        RECT 1332.680 2927.090 1333.860 2928.270 ;
        RECT 1332.680 2925.490 1333.860 2926.670 ;
        RECT 1332.680 2909.090 1333.860 2910.270 ;
        RECT 1332.680 2907.490 1333.860 2908.670 ;
        RECT 1332.680 2891.090 1333.860 2892.270 ;
        RECT 1332.680 2889.490 1333.860 2890.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 321.250 2585.090 322.430 2586.270 ;
        RECT 321.250 2583.490 322.430 2584.670 ;
        RECT 321.250 2567.090 322.430 2568.270 ;
        RECT 321.250 2565.490 322.430 2566.670 ;
        RECT 321.250 2549.090 322.430 2550.270 ;
        RECT 321.250 2547.490 322.430 2548.670 ;
        RECT 321.250 2531.090 322.430 2532.270 ;
        RECT 321.250 2529.490 322.430 2530.670 ;
        RECT 321.250 2405.090 322.430 2406.270 ;
        RECT 321.250 2403.490 322.430 2404.670 ;
        RECT 321.250 2387.090 322.430 2388.270 ;
        RECT 321.250 2385.490 322.430 2386.670 ;
        RECT 321.250 2369.090 322.430 2370.270 ;
        RECT 321.250 2367.490 322.430 2368.670 ;
        RECT 321.250 2351.090 322.430 2352.270 ;
        RECT 321.250 2349.490 322.430 2350.670 ;
        RECT 321.250 2225.090 322.430 2226.270 ;
        RECT 321.250 2223.490 322.430 2224.670 ;
        RECT 321.250 2207.090 322.430 2208.270 ;
        RECT 321.250 2205.490 322.430 2206.670 ;
        RECT 321.250 2189.090 322.430 2190.270 ;
        RECT 321.250 2187.490 322.430 2188.670 ;
        RECT 321.250 2171.090 322.430 2172.270 ;
        RECT 321.250 2169.490 322.430 2170.670 ;
        RECT 321.250 2045.090 322.430 2046.270 ;
        RECT 321.250 2043.490 322.430 2044.670 ;
        RECT 321.250 2027.090 322.430 2028.270 ;
        RECT 321.250 2025.490 322.430 2026.670 ;
        RECT 321.250 2009.090 322.430 2010.270 ;
        RECT 321.250 2007.490 322.430 2008.670 ;
        RECT 321.250 1991.090 322.430 1992.270 ;
        RECT 321.250 1989.490 322.430 1990.670 ;
        RECT 321.250 1865.090 322.430 1866.270 ;
        RECT 321.250 1863.490 322.430 1864.670 ;
        RECT 321.250 1847.090 322.430 1848.270 ;
        RECT 321.250 1845.490 322.430 1846.670 ;
        RECT 321.250 1829.090 322.430 1830.270 ;
        RECT 321.250 1827.490 322.430 1828.670 ;
        RECT 321.250 1811.090 322.430 1812.270 ;
        RECT 321.250 1809.490 322.430 1810.670 ;
        RECT 321.250 1685.090 322.430 1686.270 ;
        RECT 321.250 1683.490 322.430 1684.670 ;
        RECT 321.250 1667.090 322.430 1668.270 ;
        RECT 321.250 1665.490 322.430 1666.670 ;
        RECT 321.250 1649.090 322.430 1650.270 ;
        RECT 321.250 1647.490 322.430 1648.670 ;
        RECT 321.250 1631.090 322.430 1632.270 ;
        RECT 321.250 1629.490 322.430 1630.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1932.680 3125.090 1933.860 3126.270 ;
        RECT 1932.680 3123.490 1933.860 3124.670 ;
        RECT 1932.680 3107.090 1933.860 3108.270 ;
        RECT 1932.680 3105.490 1933.860 3106.670 ;
        RECT 1932.680 3089.090 1933.860 3090.270 ;
        RECT 1932.680 3087.490 1933.860 3088.670 ;
        RECT 1932.680 3071.090 1933.860 3072.270 ;
        RECT 1932.680 3069.490 1933.860 3070.670 ;
        RECT 1932.680 2945.090 1933.860 2946.270 ;
        RECT 1932.680 2943.490 1933.860 2944.670 ;
        RECT 1932.680 2927.090 1933.860 2928.270 ;
        RECT 1932.680 2925.490 1933.860 2926.670 ;
        RECT 1932.680 2909.090 1933.860 2910.270 ;
        RECT 1932.680 2907.490 1933.860 2908.670 ;
        RECT 1932.680 2891.090 1933.860 2892.270 ;
        RECT 1932.680 2889.490 1933.860 2890.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1702.620 2045.090 1703.800 2046.270 ;
        RECT 1702.620 2043.490 1703.800 2044.670 ;
        RECT 1702.620 2027.090 1703.800 2028.270 ;
        RECT 1702.620 2025.490 1703.800 2026.670 ;
        RECT 1702.620 2009.090 1703.800 2010.270 ;
        RECT 1702.620 2007.490 1703.800 2008.670 ;
        RECT 1702.620 1991.090 1703.800 1992.270 ;
        RECT 1702.620 1989.490 1703.800 1990.670 ;
        RECT 1702.620 1865.090 1703.800 1866.270 ;
        RECT 1702.620 1863.490 1703.800 1864.670 ;
        RECT 1702.620 1847.090 1703.800 1848.270 ;
        RECT 1702.620 1845.490 1703.800 1846.670 ;
        RECT 1702.620 1829.090 1703.800 1830.270 ;
        RECT 1702.620 1827.490 1703.800 1828.670 ;
        RECT 1702.620 1811.090 1703.800 1812.270 ;
        RECT 1702.620 1809.490 1703.800 1810.670 ;
        RECT 1702.620 1685.090 1703.800 1686.270 ;
        RECT 1702.620 1683.490 1703.800 1684.670 ;
        RECT 1702.620 1667.090 1703.800 1668.270 ;
        RECT 1702.620 1665.490 1703.800 1666.670 ;
        RECT 1702.620 1649.090 1703.800 1650.270 ;
        RECT 1702.620 1647.490 1703.800 1648.670 ;
        RECT 1702.620 1631.090 1703.800 1632.270 ;
        RECT 1702.620 1629.490 1703.800 1630.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 682.470 3126.380 684.070 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 1332.470 3126.380 1334.070 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1932.470 3126.380 1934.070 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 682.470 3123.370 684.070 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 1332.470 3123.370 1334.070 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1932.470 3123.370 1934.070 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 682.470 3108.380 684.070 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 1332.470 3108.380 1334.070 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1932.470 3108.380 1934.070 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 682.470 3105.370 684.070 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 1332.470 3105.370 1334.070 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1932.470 3105.370 1934.070 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 682.470 3090.380 684.070 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1332.470 3090.380 1334.070 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1932.470 3090.380 1934.070 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 682.470 3087.370 684.070 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1332.470 3087.370 1334.070 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1932.470 3087.370 1934.070 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 682.470 3072.380 684.070 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1332.470 3072.380 1334.070 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1932.470 3072.380 1934.070 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 682.470 3069.370 684.070 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1332.470 3069.370 1334.070 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1932.470 3069.370 1934.070 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 682.470 2946.380 684.070 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 1332.470 2946.380 1334.070 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1932.470 2946.380 1934.070 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 682.470 2943.370 684.070 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 1332.470 2943.370 1334.070 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1932.470 2943.370 1934.070 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 682.470 2928.380 684.070 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 1332.470 2928.380 1334.070 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1932.470 2928.380 1934.070 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 682.470 2925.370 684.070 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 1332.470 2925.370 1334.070 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1932.470 2925.370 1934.070 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 682.470 2910.380 684.070 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1332.470 2910.380 1334.070 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1932.470 2910.380 1934.070 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 682.470 2907.370 684.070 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1332.470 2907.370 1334.070 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1932.470 2907.370 1934.070 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 682.470 2892.380 684.070 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1332.470 2892.380 1334.070 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1932.470 2892.380 1934.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 682.470 2889.370 684.070 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1332.470 2889.370 1334.070 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1932.470 2889.370 1934.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 321.040 2586.380 322.640 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 321.040 2583.370 322.640 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 321.040 2568.380 322.640 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 321.040 2565.370 322.640 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 321.040 2550.380 322.640 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 321.040 2547.370 322.640 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 321.040 2532.380 322.640 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 321.040 2529.370 322.640 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 321.040 2406.380 322.640 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 321.040 2403.370 322.640 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 321.040 2388.380 322.640 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 321.040 2385.370 322.640 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 321.040 2370.380 322.640 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 321.040 2367.370 322.640 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 321.040 2352.380 322.640 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 321.040 2349.370 322.640 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 321.040 2226.380 322.640 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 321.040 2223.370 322.640 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 321.040 2208.380 322.640 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 321.040 2205.370 322.640 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 321.040 2190.380 322.640 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 321.040 2187.370 322.640 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 321.040 2172.380 322.640 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 321.040 2169.370 322.640 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 321.040 2046.380 322.640 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1702.410 2046.380 1704.010 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 321.040 2043.370 322.640 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1702.410 2043.370 1704.010 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 321.040 2028.380 322.640 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1702.410 2028.380 1704.010 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 321.040 2025.370 322.640 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1702.410 2025.370 1704.010 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 321.040 2010.380 322.640 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1702.410 2010.380 1704.010 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 321.040 2007.370 322.640 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1702.410 2007.370 1704.010 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 321.040 1992.380 322.640 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1702.410 1992.380 1704.010 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 321.040 1989.370 322.640 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1702.410 1989.370 1704.010 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 321.040 1866.380 322.640 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1702.410 1866.380 1704.010 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 321.040 1863.370 322.640 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1702.410 1863.370 1704.010 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 321.040 1848.380 322.640 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1702.410 1848.380 1704.010 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 321.040 1845.370 322.640 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1702.410 1845.370 1704.010 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 321.040 1830.380 322.640 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1702.410 1830.380 1704.010 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 321.040 1827.370 322.640 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1702.410 1827.370 1704.010 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 321.040 1812.380 322.640 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1702.410 1812.380 1704.010 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 321.040 1809.370 322.640 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1702.410 1809.370 1704.010 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 321.040 1686.380 322.640 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1702.410 1686.380 1704.010 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 321.040 1683.370 322.640 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1702.410 1683.370 1704.010 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 321.040 1668.380 322.640 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1702.410 1668.380 1704.010 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 321.040 1665.370 322.640 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1702.410 1665.370 1704.010 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 321.040 1650.380 322.640 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1702.410 1650.380 1704.010 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 321.040 1647.370 322.640 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1702.410 1647.370 1704.010 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 321.040 1632.380 322.640 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1702.410 1632.380 1704.010 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 321.040 1629.370 322.640 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1702.410 1629.370 1704.010 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 681.040 3251.235 686.300 3252.140 ;
        RECT 1331.040 3251.235 1336.300 3252.140 ;
        RECT 1931.040 3251.235 1936.300 3252.140 ;
        RECT 681.480 3250.400 686.300 3251.235 ;
        RECT 1331.480 3250.400 1336.300 3251.235 ;
        RECT 1931.480 3250.400 1936.300 3251.235 ;
        RECT 1700.180 1605.000 1705.000 1605.835 ;
        RECT 1700.180 1604.095 1705.440 1605.000 ;
      LAYER via3 ;
        RECT 684.720 3250.440 686.240 3252.050 ;
        RECT 1334.720 3250.440 1336.240 3252.050 ;
        RECT 1934.720 3250.440 1936.240 3252.050 ;
        RECT 1700.240 1604.185 1701.760 1605.795 ;
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 292.020 3271.235 295.020 3538.400 ;
        RECT 310.020 3271.235 313.020 3547.800 ;
        RECT 328.020 3271.235 331.020 3557.200 ;
        RECT 454.020 3271.235 457.020 3529.000 ;
        RECT 472.020 3271.235 475.020 3538.400 ;
        RECT 490.020 3271.235 493.020 3547.800 ;
        RECT 508.020 3271.235 511.020 3557.200 ;
        RECT 634.020 3271.235 637.020 3529.000 ;
        RECT 652.020 3271.235 655.020 3538.400 ;
        RECT 670.020 3271.235 673.020 3547.800 ;
        RECT 688.020 3271.235 691.020 3557.200 ;
        RECT 684.690 2804.060 686.310 3252.140 ;
        RECT 814.020 2715.000 817.020 3529.000 ;
        RECT 832.020 2715.000 835.020 3538.400 ;
        RECT 850.020 2715.000 853.020 3547.800 ;
        RECT 868.020 2715.000 871.020 3557.200 ;
        RECT 994.020 3271.235 997.020 3529.000 ;
        RECT 1012.020 3271.235 1015.020 3538.400 ;
        RECT 1030.020 3271.235 1033.020 3547.800 ;
        RECT 1048.020 3271.235 1051.020 3557.200 ;
        RECT 1174.020 3271.235 1177.020 3529.000 ;
        RECT 1192.020 3271.235 1195.020 3538.400 ;
        RECT 1210.020 3271.235 1213.020 3547.800 ;
        RECT 1228.020 3271.235 1231.020 3557.200 ;
        RECT 1334.690 2804.060 1336.310 3252.140 ;
        RECT 1354.020 2715.000 1357.020 3529.000 ;
        RECT 1372.020 2715.000 1375.020 3538.400 ;
        RECT 1390.020 2715.000 1393.020 3547.800 ;
        RECT 1408.020 2715.000 1411.020 3557.200 ;
        RECT 1534.020 3271.235 1537.020 3529.000 ;
        RECT 1552.020 3271.235 1555.020 3538.400 ;
        RECT 1570.020 3271.235 1573.020 3547.800 ;
        RECT 1588.020 3271.235 1591.020 3557.200 ;
        RECT 1714.020 3271.235 1717.020 3529.000 ;
        RECT 1732.020 3271.235 1735.020 3538.400 ;
        RECT 1750.020 3271.235 1753.020 3547.800 ;
        RECT 1768.020 3271.235 1771.020 3557.200 ;
        RECT 1894.020 3271.235 1897.020 3529.000 ;
        RECT 1912.020 3271.235 1915.020 3538.400 ;
        RECT 1930.020 3271.235 1933.020 3547.800 ;
        RECT 1948.020 3271.235 1951.020 3557.200 ;
        RECT 1934.690 2804.060 1936.310 3252.140 ;
        RECT 397.840 1610.640 399.440 2688.240 ;
        RECT 292.020 -18.720 295.020 1585.000 ;
        RECT 310.020 -28.120 313.020 1585.000 ;
        RECT 328.020 -37.520 331.020 1585.000 ;
        RECT 454.020 -9.320 457.020 1585.000 ;
        RECT 472.020 -18.720 475.020 1585.000 ;
        RECT 490.020 -28.120 493.020 1585.000 ;
        RECT 508.020 -37.520 511.020 1585.000 ;
        RECT 634.020 -9.320 637.020 1585.000 ;
        RECT 652.020 -18.720 655.020 1585.000 ;
        RECT 670.020 -28.120 673.020 1585.000 ;
        RECT 688.020 -37.520 691.020 1585.000 ;
        RECT 814.020 -9.320 817.020 1585.000 ;
        RECT 832.020 -18.720 835.020 1585.000 ;
        RECT 850.020 -28.120 853.020 1585.000 ;
        RECT 868.020 -37.520 871.020 1585.000 ;
        RECT 994.020 -9.320 997.020 1585.000 ;
        RECT 1012.020 -18.720 1015.020 1585.000 ;
        RECT 1030.020 -28.120 1033.020 1585.000 ;
        RECT 1048.020 -37.520 1051.020 1585.000 ;
        RECT 1174.020 -9.320 1177.020 1585.000 ;
        RECT 1192.020 -18.720 1195.020 1585.000 ;
        RECT 1210.020 -28.120 1213.020 1585.000 ;
        RECT 1228.020 -37.520 1231.020 1585.000 ;
        RECT 1354.020 -9.320 1357.020 1585.000 ;
        RECT 1372.020 -18.720 1375.020 1585.000 ;
        RECT 1390.020 -28.120 1393.020 1585.000 ;
        RECT 1408.020 -37.520 1411.020 1585.000 ;
        RECT 1534.020 -9.320 1537.020 2785.000 ;
        RECT 1552.020 -18.720 1555.020 2785.000 ;
        RECT 1570.020 -28.120 1573.020 2785.000 ;
        RECT 1588.020 -37.520 1591.020 2785.000 ;
        RECT 1714.020 2071.235 1717.020 2785.000 ;
        RECT 1732.020 2071.235 1735.020 2785.000 ;
        RECT 1750.020 2071.235 1753.020 2785.000 ;
        RECT 1768.020 2071.235 1771.020 2785.000 ;
        RECT 1894.020 2071.235 1897.020 2785.000 ;
        RECT 1912.020 2071.235 1915.020 2785.000 ;
        RECT 1930.020 2071.235 1933.020 2785.000 ;
        RECT 1948.020 2071.235 1951.020 2785.000 ;
        RECT 2074.020 2071.235 2077.020 3529.000 ;
        RECT 2092.020 2071.235 2095.020 3538.400 ;
        RECT 1700.170 1604.095 1701.790 2052.175 ;
        RECT 1714.020 -9.320 1717.020 1585.000 ;
        RECT 1732.020 -18.720 1735.020 1585.000 ;
        RECT 1750.020 -28.120 1753.020 1585.000 ;
        RECT 1768.020 -37.520 1771.020 1585.000 ;
        RECT 1894.020 -9.320 1897.020 1585.000 ;
        RECT 1912.020 -18.720 1915.020 1585.000 ;
        RECT 1930.020 -28.120 1933.020 1585.000 ;
        RECT 1948.020 -37.520 1951.020 1585.000 ;
        RECT 2074.020 -9.320 2077.020 1585.000 ;
        RECT 2092.020 -18.720 2095.020 1585.000 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2308.020 -37.520 2311.020 3557.200 ;
        RECT 2434.020 -9.320 2437.020 3529.000 ;
        RECT 2452.020 -18.720 2455.020 3538.400 ;
        RECT 2470.020 -28.120 2473.020 3547.800 ;
        RECT 2488.020 -37.520 2491.020 3557.200 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 684.910 3215.090 686.090 3216.270 ;
        RECT 684.910 3213.490 686.090 3214.670 ;
        RECT 684.910 3197.090 686.090 3198.270 ;
        RECT 684.910 3195.490 686.090 3196.670 ;
        RECT 684.910 3179.090 686.090 3180.270 ;
        RECT 684.910 3177.490 686.090 3178.670 ;
        RECT 684.910 3161.090 686.090 3162.270 ;
        RECT 684.910 3159.490 686.090 3160.670 ;
        RECT 684.910 3035.090 686.090 3036.270 ;
        RECT 684.910 3033.490 686.090 3034.670 ;
        RECT 684.910 3017.090 686.090 3018.270 ;
        RECT 684.910 3015.490 686.090 3016.670 ;
        RECT 684.910 2999.090 686.090 3000.270 ;
        RECT 684.910 2997.490 686.090 2998.670 ;
        RECT 684.910 2981.090 686.090 2982.270 ;
        RECT 684.910 2979.490 686.090 2980.670 ;
        RECT 684.910 2855.090 686.090 2856.270 ;
        RECT 684.910 2853.490 686.090 2854.670 ;
        RECT 684.910 2837.090 686.090 2838.270 ;
        RECT 684.910 2835.490 686.090 2836.670 ;
        RECT 684.910 2819.090 686.090 2820.270 ;
        RECT 684.910 2817.490 686.090 2818.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 1334.910 3215.090 1336.090 3216.270 ;
        RECT 1334.910 3213.490 1336.090 3214.670 ;
        RECT 1334.910 3197.090 1336.090 3198.270 ;
        RECT 1334.910 3195.490 1336.090 3196.670 ;
        RECT 1334.910 3179.090 1336.090 3180.270 ;
        RECT 1334.910 3177.490 1336.090 3178.670 ;
        RECT 1334.910 3161.090 1336.090 3162.270 ;
        RECT 1334.910 3159.490 1336.090 3160.670 ;
        RECT 1334.910 3035.090 1336.090 3036.270 ;
        RECT 1334.910 3033.490 1336.090 3034.670 ;
        RECT 1334.910 3017.090 1336.090 3018.270 ;
        RECT 1334.910 3015.490 1336.090 3016.670 ;
        RECT 1334.910 2999.090 1336.090 3000.270 ;
        RECT 1334.910 2997.490 1336.090 2998.670 ;
        RECT 1334.910 2981.090 1336.090 2982.270 ;
        RECT 1334.910 2979.490 1336.090 2980.670 ;
        RECT 1334.910 2855.090 1336.090 2856.270 ;
        RECT 1334.910 2853.490 1336.090 2854.670 ;
        RECT 1334.910 2837.090 1336.090 2838.270 ;
        RECT 1334.910 2835.490 1336.090 2836.670 ;
        RECT 1334.910 2819.090 1336.090 2820.270 ;
        RECT 1334.910 2817.490 1336.090 2818.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1934.910 3215.090 1936.090 3216.270 ;
        RECT 1934.910 3213.490 1936.090 3214.670 ;
        RECT 1934.910 3197.090 1936.090 3198.270 ;
        RECT 1934.910 3195.490 1936.090 3196.670 ;
        RECT 1934.910 3179.090 1936.090 3180.270 ;
        RECT 1934.910 3177.490 1936.090 3178.670 ;
        RECT 1934.910 3161.090 1936.090 3162.270 ;
        RECT 1934.910 3159.490 1936.090 3160.670 ;
        RECT 1934.910 3035.090 1936.090 3036.270 ;
        RECT 1934.910 3033.490 1936.090 3034.670 ;
        RECT 1934.910 3017.090 1936.090 3018.270 ;
        RECT 1934.910 3015.490 1936.090 3016.670 ;
        RECT 1934.910 2999.090 1936.090 3000.270 ;
        RECT 1934.910 2997.490 1936.090 2998.670 ;
        RECT 1934.910 2981.090 1936.090 2982.270 ;
        RECT 1934.910 2979.490 1936.090 2980.670 ;
        RECT 1934.910 2855.090 1936.090 2856.270 ;
        RECT 1934.910 2853.490 1936.090 2854.670 ;
        RECT 1934.910 2837.090 1936.090 2838.270 ;
        RECT 1934.910 2835.490 1936.090 2836.670 ;
        RECT 1934.910 2819.090 1936.090 2820.270 ;
        RECT 1934.910 2817.490 1936.090 2818.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 398.050 2675.090 399.230 2676.270 ;
        RECT 398.050 2673.490 399.230 2674.670 ;
        RECT 398.050 2657.090 399.230 2658.270 ;
        RECT 398.050 2655.490 399.230 2656.670 ;
        RECT 398.050 2639.090 399.230 2640.270 ;
        RECT 398.050 2637.490 399.230 2638.670 ;
        RECT 398.050 2621.090 399.230 2622.270 ;
        RECT 398.050 2619.490 399.230 2620.670 ;
        RECT 398.050 2495.090 399.230 2496.270 ;
        RECT 398.050 2493.490 399.230 2494.670 ;
        RECT 398.050 2477.090 399.230 2478.270 ;
        RECT 398.050 2475.490 399.230 2476.670 ;
        RECT 398.050 2459.090 399.230 2460.270 ;
        RECT 398.050 2457.490 399.230 2458.670 ;
        RECT 398.050 2441.090 399.230 2442.270 ;
        RECT 398.050 2439.490 399.230 2440.670 ;
        RECT 398.050 2315.090 399.230 2316.270 ;
        RECT 398.050 2313.490 399.230 2314.670 ;
        RECT 398.050 2297.090 399.230 2298.270 ;
        RECT 398.050 2295.490 399.230 2296.670 ;
        RECT 398.050 2279.090 399.230 2280.270 ;
        RECT 398.050 2277.490 399.230 2278.670 ;
        RECT 398.050 2261.090 399.230 2262.270 ;
        RECT 398.050 2259.490 399.230 2260.670 ;
        RECT 398.050 2135.090 399.230 2136.270 ;
        RECT 398.050 2133.490 399.230 2134.670 ;
        RECT 398.050 2117.090 399.230 2118.270 ;
        RECT 398.050 2115.490 399.230 2116.670 ;
        RECT 398.050 2099.090 399.230 2100.270 ;
        RECT 398.050 2097.490 399.230 2098.670 ;
        RECT 398.050 2081.090 399.230 2082.270 ;
        RECT 398.050 2079.490 399.230 2080.670 ;
        RECT 398.050 1955.090 399.230 1956.270 ;
        RECT 398.050 1953.490 399.230 1954.670 ;
        RECT 398.050 1937.090 399.230 1938.270 ;
        RECT 398.050 1935.490 399.230 1936.670 ;
        RECT 398.050 1919.090 399.230 1920.270 ;
        RECT 398.050 1917.490 399.230 1918.670 ;
        RECT 398.050 1901.090 399.230 1902.270 ;
        RECT 398.050 1899.490 399.230 1900.670 ;
        RECT 398.050 1775.090 399.230 1776.270 ;
        RECT 398.050 1773.490 399.230 1774.670 ;
        RECT 398.050 1757.090 399.230 1758.270 ;
        RECT 398.050 1755.490 399.230 1756.670 ;
        RECT 398.050 1739.090 399.230 1740.270 ;
        RECT 398.050 1737.490 399.230 1738.670 ;
        RECT 398.050 1721.090 399.230 1722.270 ;
        RECT 398.050 1719.490 399.230 1720.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1700.390 1955.090 1701.570 1956.270 ;
        RECT 1700.390 1953.490 1701.570 1954.670 ;
        RECT 1700.390 1937.090 1701.570 1938.270 ;
        RECT 1700.390 1935.490 1701.570 1936.670 ;
        RECT 1700.390 1919.090 1701.570 1920.270 ;
        RECT 1700.390 1917.490 1701.570 1918.670 ;
        RECT 1700.390 1901.090 1701.570 1902.270 ;
        RECT 1700.390 1899.490 1701.570 1900.670 ;
        RECT 1700.390 1775.090 1701.570 1776.270 ;
        RECT 1700.390 1773.490 1701.570 1774.670 ;
        RECT 1700.390 1757.090 1701.570 1758.270 ;
        RECT 1700.390 1755.490 1701.570 1756.670 ;
        RECT 1700.390 1739.090 1701.570 1740.270 ;
        RECT 1700.390 1737.490 1701.570 1738.670 ;
        RECT 1700.390 1721.090 1701.570 1722.270 ;
        RECT 1700.390 1719.490 1701.570 1720.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 684.690 3216.380 686.310 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1334.690 3216.380 1336.310 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1934.690 3216.380 1936.310 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 684.690 3213.370 686.310 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1334.690 3213.370 1336.310 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1934.690 3213.370 1936.310 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 684.690 3198.380 686.310 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1334.690 3198.380 1336.310 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1934.690 3198.380 1936.310 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 684.690 3195.370 686.310 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1334.690 3195.370 1336.310 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1934.690 3195.370 1936.310 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 684.690 3180.380 686.310 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1334.690 3180.380 1336.310 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1934.690 3180.380 1936.310 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 684.690 3177.370 686.310 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1334.690 3177.370 1336.310 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1934.690 3177.370 1936.310 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 684.690 3162.380 686.310 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 1334.690 3162.380 1336.310 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1934.690 3162.380 1936.310 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 684.690 3159.370 686.310 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 1334.690 3159.370 1336.310 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1934.690 3159.370 1936.310 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 684.690 3036.380 686.310 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1334.690 3036.380 1336.310 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1934.690 3036.380 1936.310 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 684.690 3033.370 686.310 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1334.690 3033.370 1336.310 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1934.690 3033.370 1936.310 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 684.690 3018.380 686.310 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1334.690 3018.380 1336.310 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1934.690 3018.380 1936.310 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 684.690 3015.370 686.310 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1334.690 3015.370 1336.310 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1934.690 3015.370 1936.310 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 684.690 3000.380 686.310 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1334.690 3000.380 1336.310 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1934.690 3000.380 1936.310 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 684.690 2997.370 686.310 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1334.690 2997.370 1336.310 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1934.690 2997.370 1936.310 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 684.690 2982.380 686.310 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 1334.690 2982.380 1336.310 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1934.690 2982.380 1936.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 684.690 2979.370 686.310 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 1334.690 2979.370 1336.310 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1934.690 2979.370 1936.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 684.690 2856.380 686.310 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1334.690 2856.380 1336.310 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1934.690 2856.380 1936.310 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 684.690 2853.370 686.310 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1334.690 2853.370 1336.310 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1934.690 2853.370 1936.310 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 684.690 2838.380 686.310 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1334.690 2838.380 1336.310 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1934.690 2838.380 1936.310 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 684.690 2835.370 686.310 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1334.690 2835.370 1336.310 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1934.690 2835.370 1936.310 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 684.690 2820.380 686.310 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1334.690 2820.380 1336.310 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1934.690 2820.380 1936.310 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 684.690 2817.370 686.310 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1334.690 2817.370 1336.310 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1934.690 2817.370 1936.310 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 397.840 2676.380 399.440 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 397.840 2673.370 399.440 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 397.840 2658.380 399.440 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 397.840 2655.370 399.440 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 397.840 2640.380 399.440 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 397.840 2637.370 399.440 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 397.840 2622.380 399.440 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 397.840 2619.370 399.440 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 397.840 2496.380 399.440 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 397.840 2493.370 399.440 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 397.840 2478.380 399.440 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 397.840 2475.370 399.440 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 397.840 2460.380 399.440 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 397.840 2457.370 399.440 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 397.840 2442.380 399.440 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 397.840 2439.370 399.440 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 397.840 2316.380 399.440 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 397.840 2313.370 399.440 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 397.840 2298.380 399.440 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 397.840 2295.370 399.440 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 397.840 2280.380 399.440 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 397.840 2277.370 399.440 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 397.840 2262.380 399.440 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 397.840 2259.370 399.440 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 397.840 2136.380 399.440 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 397.840 2133.370 399.440 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 397.840 2118.380 399.440 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 397.840 2115.370 399.440 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 397.840 2100.380 399.440 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 397.840 2097.370 399.440 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 397.840 2082.380 399.440 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 397.840 2079.370 399.440 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 397.840 1956.380 399.440 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1700.170 1956.380 1701.790 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 397.840 1953.370 399.440 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1700.170 1953.370 1701.790 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 397.840 1938.380 399.440 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1700.170 1938.380 1701.790 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 397.840 1935.370 399.440 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1700.170 1935.370 1701.790 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 397.840 1920.380 399.440 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1700.170 1920.380 1701.790 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 397.840 1917.370 399.440 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1700.170 1917.370 1701.790 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 397.840 1902.380 399.440 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1700.170 1902.380 1701.790 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 397.840 1899.370 399.440 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1700.170 1899.370 1701.790 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 397.840 1776.380 399.440 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1700.170 1776.380 1701.790 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 397.840 1773.370 399.440 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1700.170 1773.370 1701.790 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 397.840 1758.380 399.440 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1700.170 1758.380 1701.790 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 397.840 1755.370 399.440 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1700.170 1755.370 1701.790 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 397.840 1740.380 399.440 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1700.170 1740.380 1701.790 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 397.840 1737.370 399.440 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1700.170 1737.370 1701.790 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 397.840 1722.380 399.440 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1700.170 1722.380 1701.790 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 397.840 1719.370 399.440 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1700.170 1719.370 1701.790 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
        RECT 305.520 1610.795 1395.115 2688.085 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met1 ;
        RECT 1317.510 3266.960 1317.830 3267.020 ;
        RECT 1890.670 3266.960 1890.990 3267.020 ;
        RECT 1317.510 3266.820 1890.990 3266.960 ;
        RECT 1317.510 3266.760 1317.830 3266.820 ;
        RECT 1890.670 3266.760 1890.990 3266.820 ;
        RECT 696.970 3264.240 697.290 3264.300 ;
        RECT 1890.670 3264.240 1890.990 3264.300 ;
        RECT 1917.350 3264.240 1917.670 3264.300 ;
        RECT 1938.970 3264.240 1939.290 3264.300 ;
        RECT 676.360 3264.100 698.580 3264.240 ;
        RECT 646.370 3263.900 646.690 3263.960 ;
        RECT 668.450 3263.900 668.770 3263.960 ;
        RECT 676.360 3263.900 676.500 3264.100 ;
        RECT 696.970 3264.040 697.290 3264.100 ;
        RECT 646.370 3263.760 676.500 3263.900 ;
        RECT 698.440 3263.900 698.580 3264.100 ;
        RECT 1890.670 3264.100 1939.290 3264.240 ;
        RECT 1890.670 3264.040 1890.990 3264.100 ;
        RECT 1917.350 3264.040 1917.670 3264.100 ;
        RECT 1938.970 3264.040 1939.290 3264.100 ;
        RECT 1293.130 3263.900 1293.450 3263.960 ;
        RECT 1317.510 3263.900 1317.830 3263.960 ;
        RECT 698.440 3263.760 1317.830 3263.900 ;
        RECT 646.370 3263.700 646.690 3263.760 ;
        RECT 668.450 3263.700 668.770 3263.760 ;
        RECT 1293.130 3263.700 1293.450 3263.760 ;
        RECT 1317.510 3263.700 1317.830 3263.760 ;
        RECT 986.770 3254.720 987.090 3254.780 ;
        RECT 1034.610 3254.720 1034.930 3254.780 ;
        RECT 986.770 3254.580 1034.930 3254.720 ;
        RECT 986.770 3254.520 987.090 3254.580 ;
        RECT 1034.610 3254.520 1034.930 3254.580 ;
        RECT 976.190 3254.040 976.510 3254.100 ;
        RECT 986.770 3254.040 987.090 3254.100 ;
        RECT 976.190 3253.900 987.090 3254.040 ;
        RECT 976.190 3253.840 976.510 3253.900 ;
        RECT 986.770 3253.840 987.090 3253.900 ;
        RECT 1035.070 3253.020 1035.390 3253.080 ;
        RECT 1035.070 3252.880 1077.160 3253.020 ;
        RECT 1035.070 3252.820 1035.390 3252.880 ;
        RECT 1077.020 3252.680 1077.160 3252.880 ;
        RECT 1096.800 3252.880 1125.000 3253.020 ;
        RECT 1096.800 3252.680 1096.940 3252.880 ;
        RECT 886.580 3252.540 934.560 3252.680 ;
        RECT 1077.020 3252.540 1096.940 3252.680 ;
        RECT 688.230 3252.340 688.550 3252.400 ;
        RECT 737.910 3252.340 738.230 3252.400 ;
        RECT 688.230 3252.200 738.230 3252.340 ;
        RECT 688.230 3252.140 688.550 3252.200 ;
        RECT 737.910 3252.140 738.230 3252.200 ;
        RECT 738.370 3252.000 738.690 3252.060 ;
        RECT 786.210 3252.000 786.530 3252.060 ;
        RECT 738.370 3251.860 786.530 3252.000 ;
        RECT 738.370 3251.800 738.690 3251.860 ;
        RECT 786.210 3251.800 786.530 3251.860 ;
        RECT 786.670 3252.000 786.990 3252.060 ;
        RECT 786.670 3251.860 787.360 3252.000 ;
        RECT 786.670 3251.800 786.990 3251.860 ;
        RECT 787.220 3251.660 787.360 3251.860 ;
        RECT 820.710 3251.660 821.030 3251.720 ;
        RECT 787.220 3251.520 821.030 3251.660 ;
        RECT 820.710 3251.460 821.030 3251.520 ;
        RECT 821.170 3251.660 821.490 3251.720 ;
        RECT 821.170 3251.520 868.780 3251.660 ;
        RECT 821.170 3251.460 821.490 3251.520 ;
        RECT 868.640 3251.320 868.780 3251.520 ;
        RECT 886.580 3251.320 886.720 3252.540 ;
        RECT 934.420 3252.000 934.560 3252.540 ;
        RECT 1124.860 3252.340 1125.000 3252.880 ;
        RECT 1270.220 3252.880 1290.600 3253.020 ;
        RECT 1186.870 3252.680 1187.190 3252.740 ;
        RECT 1173.620 3252.540 1187.190 3252.680 ;
        RECT 1124.860 3252.200 1144.780 3252.340 ;
        RECT 976.190 3252.000 976.510 3252.060 ;
        RECT 934.420 3251.860 976.510 3252.000 ;
        RECT 1144.640 3252.000 1144.780 3252.200 ;
        RECT 1173.620 3252.000 1173.760 3252.540 ;
        RECT 1186.870 3252.480 1187.190 3252.540 ;
        RECT 1144.640 3251.860 1173.760 3252.000 ;
        RECT 1187.790 3252.000 1188.110 3252.060 ;
        RECT 1270.220 3252.000 1270.360 3252.880 ;
        RECT 1290.460 3252.340 1290.600 3252.880 ;
        RECT 1331.770 3252.340 1332.090 3252.400 ;
        RECT 1290.460 3252.200 1332.090 3252.340 ;
        RECT 1331.770 3252.140 1332.090 3252.200 ;
        RECT 1187.790 3251.860 1270.360 3252.000 ;
        RECT 976.190 3251.800 976.510 3251.860 ;
        RECT 1187.790 3251.800 1188.110 3251.860 ;
        RECT 1427.910 3251.660 1428.230 3251.720 ;
        RECT 1932.070 3251.660 1932.390 3251.720 ;
        RECT 1427.910 3251.520 1932.390 3251.660 ;
        RECT 1427.910 3251.460 1428.230 3251.520 ;
        RECT 1932.070 3251.460 1932.390 3251.520 ;
      LAYER met1 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met1 ;
        RECT 868.640 3251.180 886.720 3251.320 ;
      LAYER met1 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met1 ;
        RECT 1427.910 3250.980 1428.230 3251.040 ;
        RECT 1414.200 3250.840 1428.230 3250.980 ;
        RECT 1400.310 3250.640 1400.630 3250.700 ;
        RECT 1414.200 3250.640 1414.340 3250.840 ;
        RECT 1427.910 3250.780 1428.230 3250.840 ;
        RECT 1400.310 3250.500 1414.340 3250.640 ;
        RECT 1400.310 3250.440 1400.630 3250.500 ;
        RECT 1331.770 3250.300 1332.090 3250.360 ;
        RECT 1352.470 3250.300 1352.790 3250.360 ;
        RECT 1331.770 3250.160 1352.790 3250.300 ;
        RECT 1331.770 3250.100 1332.090 3250.160 ;
        RECT 1352.470 3250.100 1352.790 3250.160 ;
        RECT 1486.790 3229.560 1487.110 3229.620 ;
        RECT 1535.550 3229.560 1535.870 3229.620 ;
        RECT 1486.790 3229.420 1535.870 3229.560 ;
        RECT 1486.790 3229.360 1487.110 3229.420 ;
        RECT 1535.550 3229.360 1535.870 3229.420 ;
        RECT 1472.990 3222.420 1473.310 3222.480 ;
        RECT 1535.550 3222.420 1535.870 3222.480 ;
        RECT 1472.990 3222.280 1535.870 3222.420 ;
        RECT 1472.990 3222.220 1473.310 3222.280 ;
        RECT 1535.550 3222.220 1535.870 3222.280 ;
        RECT 1459.190 3215.620 1459.510 3215.680 ;
        RECT 1535.550 3215.620 1535.870 3215.680 ;
        RECT 1459.190 3215.480 1535.870 3215.620 ;
        RECT 1459.190 3215.420 1459.510 3215.480 ;
        RECT 1535.550 3215.420 1535.870 3215.480 ;
        RECT 1452.290 3208.820 1452.610 3208.880 ;
        RECT 1538.310 3208.820 1538.630 3208.880 ;
        RECT 1452.290 3208.680 1538.630 3208.820 ;
        RECT 1452.290 3208.620 1452.610 3208.680 ;
        RECT 1538.310 3208.620 1538.630 3208.680 ;
        RECT 1438.490 3201.680 1438.810 3201.740 ;
        RECT 1538.310 3201.680 1538.630 3201.740 ;
        RECT 1438.490 3201.540 1538.630 3201.680 ;
        RECT 1438.490 3201.480 1438.810 3201.540 ;
        RECT 1538.310 3201.480 1538.630 3201.540 ;
        RECT 1431.590 3194.880 1431.910 3194.940 ;
        RECT 1533.250 3194.880 1533.570 3194.940 ;
        RECT 1431.590 3194.740 1533.570 3194.880 ;
        RECT 1431.590 3194.680 1431.910 3194.740 ;
        RECT 1533.250 3194.680 1533.570 3194.740 ;
        RECT 1507.490 3188.080 1507.810 3188.140 ;
        RECT 1534.170 3188.080 1534.490 3188.140 ;
        RECT 1507.490 3187.940 1534.490 3188.080 ;
        RECT 1507.490 3187.880 1507.810 3187.940 ;
        RECT 1534.170 3187.880 1534.490 3187.940 ;
        RECT 1352.010 2946.680 1352.330 2946.740 ;
        RECT 1548.890 2946.680 1549.210 2946.740 ;
        RECT 1352.010 2946.540 1549.210 2946.680 ;
        RECT 1352.010 2946.480 1352.330 2946.540 ;
        RECT 1548.890 2946.480 1549.210 2946.540 ;
      LAYER met1 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met1 ;
        RECT 284.350 2804.560 284.670 2804.620 ;
        RECT 944.910 2804.560 945.230 2804.620 ;
        RECT 1528.190 2804.560 1528.510 2804.620 ;
        RECT 284.350 2804.420 1528.510 2804.560 ;
        RECT 284.350 2804.360 284.670 2804.420 ;
        RECT 944.910 2804.360 945.230 2804.420 ;
        RECT 1528.190 2804.360 1528.510 2804.420 ;
        RECT 1548.890 2801.160 1549.210 2801.220 ;
        RECT 1552.110 2801.160 1552.430 2801.220 ;
        RECT 1945.870 2801.160 1946.190 2801.220 ;
        RECT 1548.890 2801.020 1946.190 2801.160 ;
        RECT 1548.890 2800.960 1549.210 2801.020 ;
        RECT 1552.110 2800.960 1552.430 2801.020 ;
        RECT 1945.870 2800.960 1946.190 2801.020 ;
        RECT 310.110 2794.360 310.430 2794.420 ;
        RECT 986.770 2794.360 987.090 2794.420 ;
        RECT 310.110 2794.220 987.090 2794.360 ;
        RECT 310.110 2794.160 310.430 2794.220 ;
        RECT 986.770 2794.160 987.090 2794.220 ;
        RECT 1076.470 2794.360 1076.790 2794.420 ;
        RECT 1122.470 2794.360 1122.790 2794.420 ;
        RECT 1076.470 2794.220 1122.790 2794.360 ;
        RECT 1076.470 2794.160 1076.790 2794.220 ;
        RECT 1122.470 2794.160 1122.790 2794.220 ;
        RECT 1677.230 2794.360 1677.550 2794.420 ;
        RECT 1724.150 2794.360 1724.470 2794.420 ;
        RECT 1677.230 2794.220 1724.470 2794.360 ;
        RECT 1677.230 2794.160 1677.550 2794.220 ;
        RECT 1724.150 2794.160 1724.470 2794.220 ;
        RECT 337.250 2794.020 337.570 2794.080 ;
        RECT 1007.470 2794.020 1007.790 2794.080 ;
        RECT 337.250 2793.880 1007.790 2794.020 ;
        RECT 337.250 2793.820 337.570 2793.880 ;
        RECT 1007.470 2793.820 1007.790 2793.880 ;
        RECT 1642.270 2794.020 1642.590 2794.080 ;
        RECT 1690.110 2794.020 1690.430 2794.080 ;
        RECT 1642.270 2793.880 1690.430 2794.020 ;
        RECT 1642.270 2793.820 1642.590 2793.880 ;
        RECT 1690.110 2793.820 1690.430 2793.880 ;
        RECT 386.930 2793.680 387.250 2793.740 ;
        RECT 432.010 2793.680 432.330 2793.740 ;
        RECT 478.930 2793.680 479.250 2793.740 ;
        RECT 527.690 2793.680 528.010 2793.740 ;
        RECT 386.930 2793.540 528.010 2793.680 ;
        RECT 386.930 2793.480 387.250 2793.540 ;
        RECT 432.010 2793.480 432.330 2793.540 ;
        RECT 478.930 2793.480 479.250 2793.540 ;
        RECT 527.690 2793.480 528.010 2793.540 ;
        RECT 627.510 2793.680 627.830 2793.740 ;
        RECT 1041.970 2793.680 1042.290 2793.740 ;
        RECT 1048.410 2793.680 1048.730 2793.740 ;
        RECT 627.510 2793.540 1048.730 2793.680 ;
        RECT 627.510 2793.480 627.830 2793.540 ;
        RECT 1041.970 2793.480 1042.290 2793.540 ;
        RECT 1048.410 2793.480 1048.730 2793.540 ;
        RECT 1117.870 2793.680 1118.190 2793.740 ;
        RECT 1159.270 2793.680 1159.590 2793.740 ;
        RECT 1117.870 2793.540 1159.590 2793.680 ;
        RECT 1117.870 2793.480 1118.190 2793.540 ;
        RECT 1159.270 2793.480 1159.590 2793.540 ;
        RECT 1642.730 2793.680 1643.050 2793.740 ;
        RECT 1689.650 2793.680 1689.970 2793.740 ;
        RECT 1642.730 2793.540 1689.970 2793.680 ;
        RECT 1642.730 2793.480 1643.050 2793.540 ;
        RECT 1689.650 2793.480 1689.970 2793.540 ;
        RECT 380.030 2793.340 380.350 2793.400 ;
        RECT 421.430 2793.340 421.750 2793.400 ;
        RECT 466.510 2793.340 466.830 2793.400 ;
        RECT 380.030 2793.200 421.200 2793.340 ;
        RECT 380.030 2793.140 380.350 2793.200 ;
        RECT 421.060 2793.000 421.200 2793.200 ;
        RECT 421.430 2793.200 466.830 2793.340 ;
        RECT 421.430 2793.140 421.750 2793.200 ;
        RECT 466.510 2793.140 466.830 2793.200 ;
        RECT 489.050 2793.340 489.370 2793.400 ;
        RECT 665.690 2793.340 666.010 2793.400 ;
        RECT 489.050 2793.200 666.010 2793.340 ;
        RECT 489.050 2793.140 489.370 2793.200 ;
        RECT 665.690 2793.140 666.010 2793.200 ;
        RECT 1122.470 2793.340 1122.790 2793.400 ;
        RECT 1166.170 2793.340 1166.490 2793.400 ;
        RECT 1122.470 2793.200 1166.490 2793.340 ;
        RECT 1122.470 2793.140 1122.790 2793.200 ;
        RECT 1166.170 2793.140 1166.490 2793.200 ;
        RECT 1724.150 2793.340 1724.470 2793.400 ;
        RECT 1766.470 2793.340 1766.790 2793.400 ;
        RECT 1724.150 2793.200 1766.790 2793.340 ;
        RECT 1724.150 2793.140 1724.470 2793.200 ;
        RECT 1766.470 2793.140 1766.790 2793.200 ;
        RECT 426.030 2793.000 426.350 2793.060 ;
        RECT 474.330 2793.000 474.650 2793.060 ;
        RECT 519.410 2793.000 519.730 2793.060 ;
        RECT 520.790 2793.000 521.110 2793.060 ;
        RECT 421.060 2792.860 521.110 2793.000 ;
        RECT 426.030 2792.800 426.350 2792.860 ;
        RECT 474.330 2792.800 474.650 2792.860 ;
        RECT 519.410 2792.800 519.730 2792.860 ;
        RECT 520.790 2792.800 521.110 2792.860 ;
        RECT 524.010 2793.000 524.330 2793.060 ;
        RECT 686.850 2793.000 687.170 2793.060 ;
        RECT 524.010 2792.860 687.170 2793.000 ;
        RECT 524.010 2792.800 524.330 2792.860 ;
        RECT 686.850 2792.800 687.170 2792.860 ;
        RECT 1088.890 2793.000 1089.210 2793.060 ;
        RECT 1129.370 2793.000 1129.690 2793.060 ;
        RECT 1174.450 2793.000 1174.770 2793.060 ;
        RECT 1088.890 2792.860 1174.770 2793.000 ;
        RECT 1088.890 2792.800 1089.210 2792.860 ;
        RECT 1129.370 2792.800 1129.690 2792.860 ;
        RECT 1174.450 2792.800 1174.770 2792.860 ;
        RECT 1682.290 2793.000 1682.610 2793.060 ;
        RECT 1728.750 2793.000 1729.070 2793.060 ;
        RECT 1773.370 2793.000 1773.690 2793.060 ;
        RECT 1682.290 2792.860 1773.690 2793.000 ;
        RECT 1682.290 2792.800 1682.610 2792.860 ;
        RECT 1728.750 2792.800 1729.070 2792.860 ;
        RECT 1773.370 2792.800 1773.690 2792.860 ;
        RECT 397.970 2792.660 398.290 2792.720 ;
        RECT 444.430 2792.660 444.750 2792.720 ;
        RECT 490.430 2792.660 490.750 2792.720 ;
        RECT 397.970 2792.520 490.750 2792.660 ;
        RECT 397.970 2792.460 398.290 2792.520 ;
        RECT 444.430 2792.460 444.750 2792.520 ;
        RECT 490.430 2792.460 490.750 2792.520 ;
        RECT 497.790 2792.660 498.110 2792.720 ;
        RECT 541.490 2792.660 541.810 2792.720 ;
        RECT 497.790 2792.520 541.810 2792.660 ;
        RECT 497.790 2792.460 498.110 2792.520 ;
        RECT 541.490 2792.460 541.810 2792.520 ;
        RECT 1048.410 2792.660 1048.730 2792.720 ;
        RECT 1089.810 2792.660 1090.130 2792.720 ;
        RECT 1117.870 2792.660 1118.190 2792.720 ;
        RECT 1048.410 2792.520 1090.130 2792.660 ;
        RECT 1048.410 2792.460 1048.730 2792.520 ;
        RECT 1089.810 2792.460 1090.130 2792.520 ;
        RECT 1106.460 2792.520 1118.190 2792.660 ;
        RECT 392.450 2792.320 392.770 2792.380 ;
        RECT 439.370 2792.320 439.690 2792.380 ;
        RECT 484.910 2792.320 485.230 2792.380 ;
        RECT 534.590 2792.320 534.910 2792.380 ;
        RECT 392.450 2792.180 534.910 2792.320 ;
        RECT 392.450 2792.120 392.770 2792.180 ;
        RECT 439.370 2792.120 439.690 2792.180 ;
        RECT 484.910 2792.120 485.230 2792.180 ;
        RECT 534.590 2792.120 534.910 2792.180 ;
        RECT 542.410 2792.320 542.730 2792.380 ;
        RECT 720.890 2792.320 721.210 2792.380 ;
        RECT 542.410 2792.180 721.210 2792.320 ;
        RECT 542.410 2792.120 542.730 2792.180 ;
        RECT 720.890 2792.120 721.210 2792.180 ;
        RECT 1069.570 2792.320 1069.890 2792.380 ;
        RECT 1106.460 2792.320 1106.600 2792.520 ;
        RECT 1117.870 2792.460 1118.190 2792.520 ;
        RECT 1652.390 2792.660 1652.710 2792.720 ;
        RECT 1699.310 2792.660 1699.630 2792.720 ;
        RECT 1747.610 2792.660 1747.930 2792.720 ;
        RECT 1788.550 2792.660 1788.870 2792.720 ;
        RECT 1652.390 2792.520 1788.870 2792.660 ;
        RECT 1652.390 2792.460 1652.710 2792.520 ;
        RECT 1699.310 2792.460 1699.630 2792.520 ;
        RECT 1747.610 2792.460 1747.930 2792.520 ;
        RECT 1788.550 2792.460 1788.870 2792.520 ;
        RECT 1135.810 2792.320 1136.130 2792.380 ;
        RECT 1159.270 2792.320 1159.590 2792.380 ;
        RECT 1069.570 2792.180 1106.600 2792.320 ;
        RECT 1106.920 2792.180 1159.590 2792.320 ;
        RECT 1069.570 2792.120 1069.890 2792.180 ;
        RECT 403.950 2791.980 404.270 2792.040 ;
        RECT 449.030 2791.980 449.350 2792.040 ;
        RECT 497.790 2791.980 498.110 2792.040 ;
        RECT 502.850 2791.980 503.170 2792.040 ;
        RECT 403.950 2791.840 498.110 2791.980 ;
        RECT 403.950 2791.780 404.270 2791.840 ;
        RECT 449.030 2791.780 449.350 2791.840 ;
        RECT 497.790 2791.780 498.110 2791.840 ;
        RECT 501.560 2791.840 503.170 2791.980 ;
        RECT 363.010 2791.640 363.330 2791.700 ;
        RECT 409.470 2791.640 409.790 2791.700 ;
        RECT 455.470 2791.640 455.790 2791.700 ;
        RECT 363.010 2791.500 455.790 2791.640 ;
        RECT 363.010 2791.440 363.330 2791.500 ;
        RECT 409.470 2791.440 409.790 2791.500 ;
        RECT 455.470 2791.440 455.790 2791.500 ;
        RECT 462.370 2791.640 462.690 2791.700 ;
        RECT 489.970 2791.640 490.290 2791.700 ;
        RECT 462.370 2791.500 490.290 2791.640 ;
        RECT 462.370 2791.440 462.690 2791.500 ;
        RECT 489.970 2791.440 490.290 2791.500 ;
        RECT 490.430 2791.640 490.750 2791.700 ;
        RECT 501.560 2791.640 501.700 2791.840 ;
        RECT 502.850 2791.780 503.170 2791.840 ;
        RECT 509.750 2791.980 510.070 2792.040 ;
        RECT 700.190 2791.980 700.510 2792.040 ;
        RECT 509.750 2791.840 700.510 2791.980 ;
        RECT 509.750 2791.780 510.070 2791.840 ;
        RECT 700.190 2791.780 700.510 2791.840 ;
        RECT 1042.890 2791.980 1043.210 2792.040 ;
        RECT 1053.010 2791.980 1053.330 2792.040 ;
        RECT 1089.810 2791.980 1090.130 2792.040 ;
        RECT 1106.920 2791.980 1107.060 2792.180 ;
        RECT 1135.810 2792.120 1136.130 2792.180 ;
        RECT 1159.270 2792.120 1159.590 2792.180 ;
        RECT 1688.730 2792.320 1689.050 2792.380 ;
        RECT 1734.270 2792.320 1734.590 2792.380 ;
        RECT 1780.270 2792.320 1780.590 2792.380 ;
        RECT 1688.730 2792.180 1780.590 2792.320 ;
        RECT 1688.730 2792.120 1689.050 2792.180 ;
        RECT 1734.270 2792.120 1734.590 2792.180 ;
        RECT 1780.270 2792.120 1780.590 2792.180 ;
        RECT 1147.770 2791.980 1148.090 2792.040 ;
        RECT 1193.770 2791.980 1194.090 2792.040 ;
        RECT 1042.890 2791.840 1089.580 2791.980 ;
        RECT 1042.890 2791.780 1043.210 2791.840 ;
        RECT 1053.010 2791.780 1053.330 2791.840 ;
        RECT 490.430 2791.500 501.700 2791.640 ;
        RECT 501.930 2791.640 502.250 2791.700 ;
        RECT 700.650 2791.640 700.970 2791.700 ;
        RECT 501.930 2791.500 700.970 2791.640 ;
        RECT 490.430 2791.440 490.750 2791.500 ;
        RECT 501.930 2791.440 502.250 2791.500 ;
        RECT 700.650 2791.440 700.970 2791.500 ;
        RECT 1055.770 2791.640 1056.090 2791.700 ;
        RECT 1058.990 2791.640 1059.310 2791.700 ;
        RECT 1075.550 2791.640 1075.870 2791.700 ;
        RECT 1055.770 2791.500 1075.870 2791.640 ;
        RECT 1089.440 2791.640 1089.580 2791.840 ;
        RECT 1089.810 2791.840 1107.060 2791.980 ;
        RECT 1107.380 2791.840 1194.090 2791.980 ;
        RECT 1089.810 2791.780 1090.130 2791.840 ;
        RECT 1100.390 2791.640 1100.710 2791.700 ;
        RECT 1104.070 2791.640 1104.390 2791.700 ;
        RECT 1089.440 2791.500 1104.390 2791.640 ;
        RECT 1055.770 2791.440 1056.090 2791.500 ;
        RECT 1058.990 2791.440 1059.310 2791.500 ;
        RECT 1075.550 2791.440 1075.870 2791.500 ;
        RECT 1100.390 2791.440 1100.710 2791.500 ;
        RECT 1104.070 2791.440 1104.390 2791.500 ;
        RECT 1105.450 2791.640 1105.770 2791.700 ;
        RECT 1107.380 2791.640 1107.520 2791.840 ;
        RECT 1147.770 2791.780 1148.090 2791.840 ;
        RECT 1193.770 2791.780 1194.090 2791.840 ;
        RECT 1646.410 2791.980 1646.730 2792.040 ;
        RECT 1695.170 2791.980 1695.490 2792.040 ;
        RECT 1741.170 2791.980 1741.490 2792.040 ;
        RECT 1787.170 2791.980 1787.490 2792.040 ;
        RECT 1646.410 2791.840 1787.490 2791.980 ;
        RECT 1646.410 2791.780 1646.730 2791.840 ;
        RECT 1695.170 2791.780 1695.490 2791.840 ;
        RECT 1741.170 2791.780 1741.490 2791.840 ;
        RECT 1787.170 2791.780 1787.490 2791.840 ;
        RECT 1105.450 2791.500 1107.520 2791.640 ;
        RECT 1107.750 2791.640 1108.070 2791.700 ;
        RECT 1152.370 2791.640 1152.690 2791.700 ;
        RECT 1107.750 2791.500 1152.690 2791.640 ;
        RECT 1105.450 2791.440 1105.770 2791.500 ;
        RECT 1107.750 2791.440 1108.070 2791.500 ;
        RECT 1152.370 2791.440 1152.690 2791.500 ;
        RECT 1663.430 2791.640 1663.750 2791.700 ;
        RECT 1712.650 2791.640 1712.970 2791.700 ;
        RECT 1740.710 2791.640 1741.030 2791.700 ;
        RECT 1663.430 2791.500 1741.030 2791.640 ;
        RECT 1663.430 2791.440 1663.750 2791.500 ;
        RECT 1712.650 2791.440 1712.970 2791.500 ;
        RECT 1740.710 2791.440 1741.030 2791.500 ;
        RECT 406.250 2791.300 406.570 2791.360 ;
        RECT 727.790 2791.300 728.110 2791.360 ;
        RECT 1111.890 2791.300 1112.210 2791.360 ;
        RECT 1159.270 2791.300 1159.590 2791.360 ;
        RECT 406.250 2791.160 728.110 2791.300 ;
        RECT 406.250 2791.100 406.570 2791.160 ;
        RECT 727.790 2791.100 728.110 2791.160 ;
        RECT 1108.300 2791.160 1159.590 2791.300 ;
        RECT 384.170 2790.960 384.490 2791.020 ;
        RECT 707.090 2790.960 707.410 2791.020 ;
        RECT 384.170 2790.820 707.410 2790.960 ;
        RECT 384.170 2790.760 384.490 2790.820 ;
        RECT 707.090 2790.760 707.410 2790.820 ;
        RECT 1034.610 2790.960 1034.930 2791.020 ;
        RECT 1076.470 2790.960 1076.790 2791.020 ;
        RECT 1108.300 2790.960 1108.440 2791.160 ;
        RECT 1111.890 2791.100 1112.210 2791.160 ;
        RECT 1159.270 2791.100 1159.590 2791.160 ;
        RECT 1656.530 2791.300 1656.850 2791.360 ;
        RECT 1658.830 2791.300 1659.150 2791.360 ;
        RECT 1706.210 2791.300 1706.530 2791.360 ;
        RECT 1752.670 2791.300 1752.990 2791.360 ;
        RECT 1656.530 2791.160 1752.990 2791.300 ;
        RECT 1656.530 2791.100 1656.850 2791.160 ;
        RECT 1658.830 2791.100 1659.150 2791.160 ;
        RECT 1706.210 2791.100 1706.530 2791.160 ;
        RECT 1752.670 2791.100 1752.990 2791.160 ;
        RECT 1140.870 2790.960 1141.190 2791.020 ;
        RECT 1186.870 2790.960 1187.190 2791.020 ;
        RECT 1034.610 2790.820 1076.790 2790.960 ;
        RECT 1034.610 2790.760 1034.930 2790.820 ;
        RECT 1076.470 2790.760 1076.790 2790.820 ;
        RECT 1094.500 2790.820 1108.440 2790.960 ;
        RECT 1124.860 2790.820 1187.190 2790.960 ;
        RECT 368.990 2790.620 369.310 2790.680 ;
        RECT 414.070 2790.620 414.390 2790.680 ;
        RECT 368.990 2790.480 414.390 2790.620 ;
        RECT 368.990 2790.420 369.310 2790.480 ;
        RECT 414.070 2790.420 414.390 2790.480 ;
        RECT 419.130 2790.620 419.450 2790.680 ;
        RECT 762.290 2790.620 762.610 2790.680 ;
        RECT 419.130 2790.480 762.610 2790.620 ;
        RECT 419.130 2790.420 419.450 2790.480 ;
        RECT 762.290 2790.420 762.610 2790.480 ;
        RECT 397.050 2790.280 397.370 2790.340 ;
        RECT 741.590 2790.280 741.910 2790.340 ;
        RECT 397.050 2790.140 741.910 2790.280 ;
        RECT 397.050 2790.080 397.370 2790.140 ;
        RECT 741.590 2790.080 741.910 2790.140 ;
        RECT 371.290 2789.940 371.610 2790.000 ;
        RECT 679.490 2789.940 679.810 2790.000 ;
        RECT 371.290 2789.800 679.810 2789.940 ;
        RECT 371.290 2789.740 371.610 2789.800 ;
        RECT 679.490 2789.740 679.810 2789.800 ;
        RECT 1017.590 2789.940 1017.910 2790.000 ;
        RECT 1065.430 2789.940 1065.750 2790.000 ;
        RECT 1094.500 2789.940 1094.640 2790.820 ;
        RECT 1094.870 2790.280 1095.190 2790.340 ;
        RECT 1124.860 2790.280 1125.000 2790.820 ;
        RECT 1140.870 2790.760 1141.190 2790.820 ;
        RECT 1186.870 2790.760 1187.190 2790.820 ;
        RECT 1670.330 2790.960 1670.650 2791.020 ;
        RECT 1718.170 2790.960 1718.490 2791.020 ;
        RECT 1759.570 2790.960 1759.890 2791.020 ;
        RECT 1670.330 2790.820 1759.890 2790.960 ;
        RECT 1670.330 2790.760 1670.650 2790.820 ;
        RECT 1718.170 2790.760 1718.490 2790.820 ;
        RECT 1759.570 2790.760 1759.890 2790.820 ;
        RECT 1418.710 2790.620 1419.030 2790.680 ;
        RECT 1773.370 2790.620 1773.690 2790.680 ;
        RECT 1418.710 2790.480 1773.690 2790.620 ;
        RECT 1418.710 2790.420 1419.030 2790.480 ;
        RECT 1773.370 2790.420 1773.690 2790.480 ;
        RECT 1094.870 2790.140 1125.000 2790.280 ;
        RECT 1094.870 2790.080 1095.190 2790.140 ;
        RECT 1017.590 2789.800 1094.640 2789.940 ;
        RECT 1631.690 2789.940 1632.010 2790.000 ;
        RECT 1677.230 2789.940 1677.550 2790.000 ;
        RECT 1631.690 2789.800 1677.550 2789.940 ;
        RECT 1017.590 2789.740 1017.910 2789.800 ;
        RECT 1065.430 2789.740 1065.750 2789.800 ;
        RECT 1631.690 2789.740 1632.010 2789.800 ;
        RECT 1677.230 2789.740 1677.550 2789.800 ;
        RECT 414.070 2789.600 414.390 2789.660 ;
        RECT 462.370 2789.600 462.690 2789.660 ;
        RECT 414.070 2789.460 462.690 2789.600 ;
        RECT 414.070 2789.400 414.390 2789.460 ;
        RECT 462.370 2789.400 462.690 2789.460 ;
        RECT 468.810 2789.600 469.130 2789.660 ;
        RECT 636.250 2789.600 636.570 2789.660 ;
        RECT 468.810 2789.460 636.570 2789.600 ;
        RECT 468.810 2789.400 469.130 2789.460 ;
        RECT 636.250 2789.400 636.570 2789.460 ;
        RECT 648.210 2789.600 648.530 2789.660 ;
        RECT 1042.890 2789.600 1043.210 2789.660 ;
        RECT 648.210 2789.460 1043.210 2789.600 ;
        RECT 648.210 2789.400 648.530 2789.460 ;
        RECT 1042.890 2789.400 1043.210 2789.460 ;
        RECT 1514.390 2789.600 1514.710 2789.660 ;
        RECT 1587.070 2789.600 1587.390 2789.660 ;
        RECT 1514.390 2789.460 1587.390 2789.600 ;
        RECT 1514.390 2789.400 1514.710 2789.460 ;
        RECT 1587.070 2789.400 1587.390 2789.460 ;
        RECT 1617.890 2789.600 1618.210 2789.660 ;
        RECT 1663.430 2789.600 1663.750 2789.660 ;
        RECT 1617.890 2789.460 1663.750 2789.600 ;
        RECT 1617.890 2789.400 1618.210 2789.460 ;
        RECT 1663.430 2789.400 1663.750 2789.460 ;
        RECT 399.810 2789.260 400.130 2789.320 ;
        RECT 514.350 2789.260 514.670 2789.320 ;
        RECT 399.810 2789.120 514.670 2789.260 ;
        RECT 399.810 2789.060 400.130 2789.120 ;
        RECT 514.350 2789.060 514.670 2789.120 ;
        RECT 606.810 2789.260 607.130 2789.320 ;
        RECT 1030.470 2789.260 1030.790 2789.320 ;
        RECT 1034.610 2789.260 1034.930 2789.320 ;
        RECT 606.810 2789.120 1034.930 2789.260 ;
        RECT 606.810 2789.060 607.130 2789.120 ;
        RECT 1030.470 2789.060 1030.790 2789.120 ;
        RECT 1034.610 2789.060 1034.930 2789.120 ;
        RECT 1045.190 2789.260 1045.510 2789.320 ;
        RECT 1094.870 2789.260 1095.190 2789.320 ;
        RECT 1045.190 2789.120 1095.190 2789.260 ;
        RECT 1045.190 2789.060 1045.510 2789.120 ;
        RECT 1094.870 2789.060 1095.190 2789.120 ;
        RECT 1487.250 2789.260 1487.570 2789.320 ;
        RECT 1600.870 2789.260 1601.190 2789.320 ;
        RECT 1487.250 2789.120 1601.190 2789.260 ;
        RECT 1487.250 2789.060 1487.570 2789.120 ;
        RECT 1600.870 2789.060 1601.190 2789.120 ;
        RECT 1610.990 2789.260 1611.310 2789.320 ;
        RECT 1656.530 2789.260 1656.850 2789.320 ;
        RECT 1610.990 2789.120 1656.850 2789.260 ;
        RECT 1610.990 2789.060 1611.310 2789.120 ;
        RECT 1656.530 2789.060 1656.850 2789.120 ;
        RECT 330.810 2788.920 331.130 2788.980 ;
        RECT 1001.030 2788.920 1001.350 2788.980 ;
        RECT 330.810 2788.780 1001.350 2788.920 ;
        RECT 330.810 2788.720 331.130 2788.780 ;
        RECT 1001.030 2788.720 1001.350 2788.780 ;
        RECT 1010.690 2788.920 1011.010 2788.980 ;
        RECT 1055.770 2788.920 1056.090 2788.980 ;
        RECT 1010.690 2788.780 1056.090 2788.920 ;
        RECT 1010.690 2788.720 1011.010 2788.780 ;
        RECT 1055.770 2788.720 1056.090 2788.780 ;
        RECT 1624.790 2788.920 1625.110 2788.980 ;
        RECT 1670.330 2788.920 1670.650 2788.980 ;
        RECT 1624.790 2788.780 1670.650 2788.920 ;
        RECT 1624.790 2788.720 1625.110 2788.780 ;
        RECT 1670.330 2788.720 1670.650 2788.780 ;
        RECT 374.970 2788.580 375.290 2788.640 ;
        RECT 420.970 2788.580 421.290 2788.640 ;
        RECT 374.970 2788.440 421.290 2788.580 ;
        RECT 374.970 2788.380 375.290 2788.440 ;
        RECT 420.970 2788.380 421.290 2788.440 ;
        RECT 466.510 2788.580 466.830 2788.640 ;
        RECT 499.170 2788.580 499.490 2788.640 ;
        RECT 466.510 2788.440 499.490 2788.580 ;
        RECT 466.510 2788.380 466.830 2788.440 ;
        RECT 499.170 2788.380 499.490 2788.440 ;
        RECT 537.350 2788.580 537.670 2788.640 ;
        RECT 707.550 2788.580 707.870 2788.640 ;
        RECT 537.350 2788.440 707.870 2788.580 ;
        RECT 537.350 2788.380 537.670 2788.440 ;
        RECT 707.550 2788.380 707.870 2788.440 ;
        RECT 1024.490 2788.580 1024.810 2788.640 ;
        RECT 1069.570 2788.580 1069.890 2788.640 ;
        RECT 1024.490 2788.440 1069.890 2788.580 ;
        RECT 1024.490 2788.380 1024.810 2788.440 ;
        RECT 1069.570 2788.380 1069.890 2788.440 ;
        RECT 1418.250 2788.580 1418.570 2788.640 ;
        RECT 1759.570 2788.580 1759.890 2788.640 ;
        RECT 1418.250 2788.440 1759.890 2788.580 ;
        RECT 1418.250 2788.380 1418.570 2788.440 ;
        RECT 1759.570 2788.380 1759.890 2788.440 ;
        RECT 317.010 2788.240 317.330 2788.300 ;
        RECT 993.670 2788.240 993.990 2788.300 ;
        RECT 317.010 2788.100 993.990 2788.240 ;
        RECT 317.010 2788.040 317.330 2788.100 ;
        RECT 993.670 2788.040 993.990 2788.100 ;
        RECT 1038.290 2788.240 1038.610 2788.300 ;
        RECT 1088.890 2788.240 1089.210 2788.300 ;
        RECT 1038.290 2788.100 1089.210 2788.240 ;
        RECT 1038.290 2788.040 1038.610 2788.100 ;
        RECT 1088.890 2788.040 1089.210 2788.100 ;
        RECT 1417.790 2788.240 1418.110 2788.300 ;
        RECT 1766.470 2788.240 1766.790 2788.300 ;
        RECT 1417.790 2788.100 1766.790 2788.240 ;
        RECT 1417.790 2788.040 1418.110 2788.100 ;
        RECT 1766.470 2788.040 1766.790 2788.100 ;
        RECT 455.470 2787.900 455.790 2787.960 ;
        RECT 500.090 2787.900 500.410 2787.960 ;
        RECT 513.890 2787.900 514.210 2787.960 ;
        RECT 538.730 2787.900 539.050 2787.960 ;
        RECT 542.410 2787.900 542.730 2787.960 ;
        RECT 455.470 2787.760 500.410 2787.900 ;
        RECT 455.470 2787.700 455.790 2787.760 ;
        RECT 500.090 2787.700 500.410 2787.760 ;
        RECT 500.640 2787.760 514.210 2787.900 ;
        RECT 499.170 2787.560 499.490 2787.620 ;
        RECT 500.640 2787.560 500.780 2787.760 ;
        RECT 513.890 2787.700 514.210 2787.760 ;
        RECT 514.440 2787.760 542.730 2787.900 ;
        RECT 499.170 2787.420 500.780 2787.560 ;
        RECT 502.850 2787.560 503.170 2787.620 ;
        RECT 514.440 2787.560 514.580 2787.760 ;
        RECT 538.730 2787.700 539.050 2787.760 ;
        RECT 542.410 2787.700 542.730 2787.760 ;
        RECT 636.250 2787.900 636.570 2787.960 ;
        RECT 658.790 2787.900 659.110 2787.960 ;
        RECT 636.250 2787.760 659.110 2787.900 ;
        RECT 636.250 2787.700 636.570 2787.760 ;
        RECT 658.790 2787.700 659.110 2787.760 ;
        RECT 1638.590 2787.900 1638.910 2787.960 ;
        RECT 1682.290 2787.900 1682.610 2787.960 ;
        RECT 1638.590 2787.760 1682.610 2787.900 ;
        RECT 1638.590 2787.700 1638.910 2787.760 ;
        RECT 1682.290 2787.700 1682.610 2787.760 ;
        RECT 502.850 2787.420 514.580 2787.560 ;
        RECT 499.170 2787.360 499.490 2787.420 ;
        RECT 502.850 2787.360 503.170 2787.420 ;
        RECT 387.850 2728.740 388.170 2728.800 ;
        RECT 943.990 2728.740 944.310 2728.800 ;
        RECT 387.850 2728.600 944.310 2728.740 ;
        RECT 387.850 2728.540 388.170 2728.600 ;
        RECT 943.990 2728.540 944.310 2728.600 ;
        RECT 288.030 2725.340 288.350 2725.400 ;
        RECT 564.030 2725.340 564.350 2725.400 ;
        RECT 288.030 2725.200 564.350 2725.340 ;
        RECT 288.030 2725.140 288.350 2725.200 ;
        RECT 564.030 2725.140 564.350 2725.200 ;
        RECT 574.610 2725.340 574.930 2725.400 ;
        RECT 1010.690 2725.340 1011.010 2725.400 ;
        RECT 574.610 2725.200 1011.010 2725.340 ;
        RECT 574.610 2725.140 574.930 2725.200 ;
        RECT 1010.690 2725.140 1011.010 2725.200 ;
        RECT 448.110 2725.000 448.430 2725.060 ;
        RECT 886.030 2725.000 886.350 2725.060 ;
        RECT 448.110 2724.860 886.350 2725.000 ;
        RECT 448.110 2724.800 448.430 2724.860 ;
        RECT 886.030 2724.800 886.350 2724.860 ;
        RECT 461.910 2724.660 462.230 2724.720 ;
        RECT 906.730 2724.660 907.050 2724.720 ;
        RECT 461.910 2724.520 907.050 2724.660 ;
        RECT 461.910 2724.460 462.230 2724.520 ;
        RECT 906.730 2724.460 907.050 2724.520 ;
        RECT 481.230 2724.320 481.550 2724.380 ;
        RECT 941.690 2724.320 942.010 2724.380 ;
        RECT 481.230 2724.180 942.010 2724.320 ;
        RECT 481.230 2724.120 481.550 2724.180 ;
        RECT 941.690 2724.120 942.010 2724.180 ;
        RECT 455.010 2723.980 455.330 2724.040 ;
        RECT 896.150 2723.980 896.470 2724.040 ;
        RECT 455.010 2723.840 896.470 2723.980 ;
        RECT 455.010 2723.780 455.330 2723.840 ;
        RECT 896.150 2723.780 896.470 2723.840 ;
        RECT 482.610 2723.640 482.930 2723.700 ;
        RECT 948.130 2723.640 948.450 2723.700 ;
        RECT 482.610 2723.500 948.450 2723.640 ;
        RECT 482.610 2723.440 482.930 2723.500 ;
        RECT 948.130 2723.440 948.450 2723.500 ;
        RECT 470.650 2723.300 470.970 2723.360 ;
        RECT 942.150 2723.300 942.470 2723.360 ;
        RECT 470.650 2723.160 942.470 2723.300 ;
        RECT 470.650 2723.100 470.970 2723.160 ;
        RECT 942.150 2723.100 942.470 2723.160 ;
        RECT 449.950 2722.960 450.270 2723.020 ;
        RECT 943.070 2722.960 943.390 2723.020 ;
        RECT 449.950 2722.820 943.390 2722.960 ;
        RECT 449.950 2722.760 450.270 2722.820 ;
        RECT 943.070 2722.760 943.390 2722.820 ;
        RECT 285.270 2722.620 285.590 2722.680 ;
        RECT 512.510 2722.620 512.830 2722.680 ;
        RECT 285.270 2722.480 512.830 2722.620 ;
        RECT 285.270 2722.420 285.590 2722.480 ;
        RECT 512.510 2722.420 512.830 2722.480 ;
        RECT 517.110 2722.620 517.430 2722.680 ;
        RECT 1010.230 2722.620 1010.550 2722.680 ;
        RECT 517.110 2722.480 1010.550 2722.620 ;
        RECT 517.110 2722.420 517.430 2722.480 ;
        RECT 1010.230 2722.420 1010.550 2722.480 ;
        RECT 287.110 2722.280 287.430 2722.340 ;
        RECT 543.330 2722.280 543.650 2722.340 ;
        RECT 287.110 2722.140 543.650 2722.280 ;
        RECT 287.110 2722.080 287.430 2722.140 ;
        RECT 543.330 2722.080 543.650 2722.140 ;
        RECT 551.610 2722.280 551.930 2722.340 ;
        RECT 1060.830 2722.280 1061.150 2722.340 ;
        RECT 551.610 2722.140 1061.150 2722.280 ;
        RECT 551.610 2722.080 551.930 2722.140 ;
        RECT 1060.830 2722.080 1061.150 2722.140 ;
        RECT 408.550 2721.940 408.870 2722.000 ;
        RECT 979.870 2721.940 980.190 2722.000 ;
        RECT 408.550 2721.800 980.190 2721.940 ;
        RECT 408.550 2721.740 408.870 2721.800 ;
        RECT 979.870 2721.740 980.190 2721.800 ;
        RECT 434.310 2721.600 434.630 2721.660 ;
        RECT 865.330 2721.600 865.650 2721.660 ;
        RECT 434.310 2721.460 865.650 2721.600 ;
        RECT 434.310 2721.400 434.630 2721.460 ;
        RECT 865.330 2721.400 865.650 2721.460 ;
        RECT 441.210 2721.260 441.530 2721.320 ;
        RECT 875.450 2721.260 875.770 2721.320 ;
        RECT 441.210 2721.120 875.770 2721.260 ;
        RECT 441.210 2721.060 441.530 2721.120 ;
        RECT 875.450 2721.060 875.770 2721.120 ;
        RECT 433.850 2720.920 434.170 2720.980 ;
        RECT 854.750 2720.920 855.070 2720.980 ;
        RECT 433.850 2720.780 855.070 2720.920 ;
        RECT 433.850 2720.720 434.170 2720.780 ;
        RECT 854.750 2720.720 855.070 2720.780 ;
        RECT 427.410 2720.580 427.730 2720.640 ;
        RECT 844.170 2720.580 844.490 2720.640 ;
        RECT 427.410 2720.440 844.490 2720.580 ;
        RECT 427.410 2720.380 427.730 2720.440 ;
        RECT 844.170 2720.380 844.490 2720.440 ;
        RECT 365.310 2720.240 365.630 2720.300 ;
        RECT 740.670 2720.240 740.990 2720.300 ;
        RECT 365.310 2720.100 740.990 2720.240 ;
        RECT 365.310 2720.040 365.630 2720.100 ;
        RECT 740.670 2720.040 740.990 2720.100 ;
        RECT 514.350 2719.900 514.670 2719.960 ;
        RECT 802.770 2719.900 803.090 2719.960 ;
        RECT 514.350 2719.760 803.090 2719.900 ;
        RECT 514.350 2719.700 514.670 2719.760 ;
        RECT 802.770 2719.700 803.090 2719.760 ;
        RECT 287.570 2719.560 287.890 2719.620 ;
        RECT 553.910 2719.560 554.230 2719.620 ;
        RECT 287.570 2719.420 554.230 2719.560 ;
        RECT 287.570 2719.360 287.890 2719.420 ;
        RECT 553.910 2719.360 554.230 2719.420 ;
        RECT 286.650 2719.220 286.970 2719.280 ;
        RECT 533.210 2719.220 533.530 2719.280 ;
        RECT 286.650 2719.080 533.530 2719.220 ;
        RECT 286.650 2719.020 286.970 2719.080 ;
        RECT 533.210 2719.020 533.530 2719.080 ;
        RECT 286.190 2718.880 286.510 2718.940 ;
        RECT 522.630 2718.880 522.950 2718.940 ;
        RECT 286.190 2718.740 522.950 2718.880 ;
        RECT 286.190 2718.680 286.510 2718.740 ;
        RECT 522.630 2718.680 522.950 2718.740 ;
        RECT 358.410 2718.540 358.730 2718.600 ;
        RECT 377.270 2718.540 377.590 2718.600 ;
        RECT 358.410 2718.400 377.590 2718.540 ;
        RECT 358.410 2718.340 358.730 2718.400 ;
        RECT 377.270 2718.340 377.590 2718.400 ;
        RECT 379.110 2718.540 379.430 2718.600 ;
        RECT 761.370 2718.540 761.690 2718.600 ;
        RECT 379.110 2718.400 761.690 2718.540 ;
        RECT 379.110 2718.340 379.430 2718.400 ;
        RECT 761.370 2718.340 761.690 2718.400 ;
        RECT 762.290 2718.540 762.610 2718.600 ;
        RECT 834.050 2718.540 834.370 2718.600 ;
        RECT 762.290 2718.400 834.370 2718.540 ;
        RECT 762.290 2718.340 762.610 2718.400 ;
        RECT 834.050 2718.340 834.370 2718.400 ;
        RECT 1034.610 2718.540 1034.930 2718.600 ;
        RECT 1102.230 2718.540 1102.550 2718.600 ;
        RECT 1034.610 2718.400 1102.550 2718.540 ;
        RECT 1034.610 2718.340 1034.930 2718.400 ;
        RECT 1102.230 2718.340 1102.550 2718.400 ;
        RECT 1145.010 2718.540 1145.330 2718.600 ;
        RECT 1300.950 2718.540 1301.270 2718.600 ;
        RECT 1145.010 2718.400 1301.270 2718.540 ;
        RECT 1145.010 2718.340 1145.330 2718.400 ;
        RECT 1300.950 2718.340 1301.270 2718.400 ;
        RECT 392.910 2718.200 393.230 2718.260 ;
        RECT 782.070 2718.200 782.390 2718.260 ;
        RECT 392.910 2718.060 782.390 2718.200 ;
        RECT 392.910 2718.000 393.230 2718.060 ;
        RECT 782.070 2718.000 782.390 2718.060 ;
        RECT 1027.710 2718.200 1028.030 2718.260 ;
        RECT 1093.490 2718.200 1093.810 2718.260 ;
        RECT 1027.710 2718.060 1093.810 2718.200 ;
        RECT 1027.710 2718.000 1028.030 2718.060 ;
        RECT 1093.490 2718.000 1093.810 2718.060 ;
        RECT 1138.110 2718.200 1138.430 2718.260 ;
        RECT 1290.370 2718.200 1290.690 2718.260 ;
        RECT 1138.110 2718.060 1290.690 2718.200 ;
        RECT 1138.110 2718.000 1138.430 2718.060 ;
        RECT 1290.370 2718.000 1290.690 2718.060 ;
        RECT 305.050 2717.860 305.370 2717.920 ;
        RECT 310.110 2717.860 310.430 2717.920 ;
        RECT 305.050 2717.720 310.430 2717.860 ;
        RECT 305.050 2717.660 305.370 2717.720 ;
        RECT 310.110 2717.660 310.430 2717.720 ;
        RECT 351.050 2717.860 351.370 2717.920 ;
        RECT 356.570 2717.860 356.890 2717.920 ;
        RECT 351.050 2717.720 356.890 2717.860 ;
        RECT 351.050 2717.660 351.370 2717.720 ;
        RECT 356.570 2717.660 356.890 2717.720 ;
        RECT 413.610 2717.860 413.930 2717.920 ;
        RECT 823.470 2717.860 823.790 2717.920 ;
        RECT 413.610 2717.720 823.790 2717.860 ;
        RECT 413.610 2717.660 413.930 2717.720 ;
        RECT 823.470 2717.660 823.790 2717.720 ;
        RECT 1041.510 2717.860 1041.830 2717.920 ;
        RECT 1114.190 2717.860 1114.510 2717.920 ;
        RECT 1041.510 2717.720 1114.510 2717.860 ;
        RECT 1041.510 2717.660 1041.830 2717.720 ;
        RECT 1114.190 2717.660 1114.510 2717.720 ;
        RECT 1151.910 2717.860 1152.230 2717.920 ;
        RECT 1311.070 2717.860 1311.390 2717.920 ;
        RECT 1151.910 2717.720 1311.390 2717.860 ;
        RECT 1151.910 2717.660 1152.230 2717.720 ;
        RECT 1311.070 2717.660 1311.390 2717.720 ;
        RECT 636.710 2717.520 637.030 2717.580 ;
        RECT 1045.190 2717.520 1045.510 2717.580 ;
        RECT 636.710 2717.380 1045.510 2717.520 ;
        RECT 636.710 2717.320 637.030 2717.380 ;
        RECT 1045.190 2717.320 1045.510 2717.380 ;
        RECT 1048.410 2717.520 1048.730 2717.580 ;
        RECT 1122.470 2717.520 1122.790 2717.580 ;
        RECT 1048.410 2717.380 1122.790 2717.520 ;
        RECT 1048.410 2717.320 1048.730 2717.380 ;
        RECT 1122.470 2717.320 1122.790 2717.380 ;
        RECT 1158.810 2717.520 1159.130 2717.580 ;
        RECT 1321.650 2717.520 1321.970 2717.580 ;
        RECT 1158.810 2717.380 1321.970 2717.520 ;
        RECT 1158.810 2717.320 1159.130 2717.380 ;
        RECT 1321.650 2717.320 1321.970 2717.380 ;
        RECT 616.010 2717.180 616.330 2717.240 ;
        RECT 1038.290 2717.180 1038.610 2717.240 ;
        RECT 616.010 2717.040 1038.610 2717.180 ;
        RECT 616.010 2716.980 616.330 2717.040 ;
        RECT 1038.290 2716.980 1038.610 2717.040 ;
        RECT 1055.310 2717.180 1055.630 2717.240 ;
        RECT 1134.890 2717.180 1135.210 2717.240 ;
        RECT 1055.310 2717.040 1135.210 2717.180 ;
        RECT 1055.310 2716.980 1055.630 2717.040 ;
        RECT 1134.890 2716.980 1135.210 2717.040 ;
        RECT 1165.710 2717.180 1166.030 2717.240 ;
        RECT 1332.230 2717.180 1332.550 2717.240 ;
        RECT 1165.710 2717.040 1332.550 2717.180 ;
        RECT 1165.710 2716.980 1166.030 2717.040 ;
        RECT 1332.230 2716.980 1332.550 2717.040 ;
        RECT 595.310 2716.840 595.630 2716.900 ;
        RECT 1024.490 2716.840 1024.810 2716.900 ;
        RECT 595.310 2716.700 1024.810 2716.840 ;
        RECT 595.310 2716.640 595.630 2716.700 ;
        RECT 1024.490 2716.640 1024.810 2716.700 ;
        RECT 1062.210 2716.840 1062.530 2716.900 ;
        RECT 1155.590 2716.840 1155.910 2716.900 ;
        RECT 1062.210 2716.700 1155.910 2716.840 ;
        RECT 1062.210 2716.640 1062.530 2716.700 ;
        RECT 1155.590 2716.640 1155.910 2716.700 ;
        RECT 1165.250 2716.840 1165.570 2716.900 ;
        RECT 1342.350 2716.840 1342.670 2716.900 ;
        RECT 1165.250 2716.700 1342.670 2716.840 ;
        RECT 1165.250 2716.640 1165.570 2716.700 ;
        RECT 1342.350 2716.640 1342.670 2716.700 ;
        RECT 585.190 2716.500 585.510 2716.560 ;
        RECT 1017.590 2716.500 1017.910 2716.560 ;
        RECT 585.190 2716.360 1017.910 2716.500 ;
        RECT 585.190 2716.300 585.510 2716.360 ;
        RECT 1017.590 2716.300 1017.910 2716.360 ;
        RECT 1076.010 2716.500 1076.330 2716.560 ;
        RECT 1176.290 2716.500 1176.610 2716.560 ;
        RECT 1076.010 2716.360 1176.610 2716.500 ;
        RECT 1076.010 2716.300 1076.330 2716.360 ;
        RECT 1176.290 2716.300 1176.610 2716.360 ;
        RECT 1179.510 2716.500 1179.830 2716.560 ;
        RECT 1363.050 2716.500 1363.370 2716.560 ;
        RECT 1179.510 2716.360 1363.370 2716.500 ;
        RECT 1179.510 2716.300 1179.830 2716.360 ;
        RECT 1363.050 2716.300 1363.370 2716.360 ;
        RECT 468.350 2716.160 468.670 2716.220 ;
        RECT 916.850 2716.160 917.170 2716.220 ;
        RECT 468.350 2716.020 917.170 2716.160 ;
        RECT 468.350 2715.960 468.670 2716.020 ;
        RECT 916.850 2715.960 917.170 2716.020 ;
        RECT 1054.850 2716.160 1055.170 2716.220 ;
        RECT 1145.470 2716.160 1145.790 2716.220 ;
        RECT 1054.850 2716.020 1145.790 2716.160 ;
        RECT 1054.850 2715.960 1055.170 2716.020 ;
        RECT 1145.470 2715.960 1145.790 2716.020 ;
        RECT 1172.610 2716.160 1172.930 2716.220 ;
        RECT 1352.930 2716.160 1353.250 2716.220 ;
        RECT 1172.610 2716.020 1353.250 2716.160 ;
        RECT 1172.610 2715.960 1172.930 2716.020 ;
        RECT 1352.930 2715.960 1353.250 2716.020 ;
        RECT 284.810 2715.820 285.130 2715.880 ;
        RECT 398.430 2715.820 398.750 2715.880 ;
        RECT 284.810 2715.680 398.750 2715.820 ;
        RECT 284.810 2715.620 285.130 2715.680 ;
        RECT 398.430 2715.620 398.750 2715.680 ;
        RECT 475.710 2715.820 476.030 2715.880 ;
        RECT 937.550 2715.820 937.870 2715.880 ;
        RECT 475.710 2715.680 937.870 2715.820 ;
        RECT 475.710 2715.620 476.030 2715.680 ;
        RECT 937.550 2715.620 937.870 2715.680 ;
        RECT 1020.810 2715.820 1021.130 2715.880 ;
        RECT 1081.070 2715.820 1081.390 2715.880 ;
        RECT 1020.810 2715.680 1081.390 2715.820 ;
        RECT 1020.810 2715.620 1021.130 2715.680 ;
        RECT 1081.070 2715.620 1081.390 2715.680 ;
        RECT 1082.910 2715.820 1083.230 2715.880 ;
        RECT 1186.870 2715.820 1187.190 2715.880 ;
        RECT 1082.910 2715.680 1187.190 2715.820 ;
        RECT 1082.910 2715.620 1083.230 2715.680 ;
        RECT 1186.870 2715.620 1187.190 2715.680 ;
        RECT 1193.310 2715.820 1193.630 2715.880 ;
        RECT 1383.750 2715.820 1384.070 2715.880 ;
        RECT 1193.310 2715.680 1384.070 2715.820 ;
        RECT 1193.310 2715.620 1193.630 2715.680 ;
        RECT 1383.750 2715.620 1384.070 2715.680 ;
        RECT 337.710 2715.480 338.030 2715.540 ;
        RECT 491.810 2715.480 492.130 2715.540 ;
        RECT 337.710 2715.340 492.130 2715.480 ;
        RECT 337.710 2715.280 338.030 2715.340 ;
        RECT 491.810 2715.280 492.130 2715.340 ;
        RECT 496.410 2715.480 496.730 2715.540 ;
        RECT 968.830 2715.480 969.150 2715.540 ;
        RECT 496.410 2715.340 969.150 2715.480 ;
        RECT 496.410 2715.280 496.730 2715.340 ;
        RECT 968.830 2715.280 969.150 2715.340 ;
        RECT 1069.110 2715.480 1069.430 2715.540 ;
        RECT 1166.170 2715.480 1166.490 2715.540 ;
        RECT 1069.110 2715.340 1166.490 2715.480 ;
        RECT 1069.110 2715.280 1069.430 2715.340 ;
        RECT 1166.170 2715.280 1166.490 2715.340 ;
        RECT 1186.410 2715.480 1186.730 2715.540 ;
        RECT 1373.630 2715.480 1373.950 2715.540 ;
        RECT 1186.410 2715.340 1373.950 2715.480 ;
        RECT 1186.410 2715.280 1186.730 2715.340 ;
        RECT 1373.630 2715.280 1373.950 2715.340 ;
        RECT 285.730 2715.140 286.050 2715.200 ;
        RECT 501.930 2715.140 502.250 2715.200 ;
        RECT 285.730 2715.000 502.250 2715.140 ;
        RECT 285.730 2714.940 286.050 2715.000 ;
        RECT 501.930 2714.940 502.250 2715.000 ;
        RECT 510.210 2715.140 510.530 2715.200 ;
        RECT 989.530 2715.140 989.850 2715.200 ;
        RECT 510.210 2715.000 989.850 2715.140 ;
        RECT 510.210 2714.940 510.530 2715.000 ;
        RECT 989.530 2714.940 989.850 2715.000 ;
        RECT 1013.910 2715.140 1014.230 2715.200 ;
        RECT 1072.790 2715.140 1073.110 2715.200 ;
        RECT 1013.910 2715.000 1073.110 2715.140 ;
        RECT 1013.910 2714.940 1014.230 2715.000 ;
        RECT 1072.790 2714.940 1073.110 2715.000 ;
        RECT 1089.350 2715.140 1089.670 2715.200 ;
        RECT 1196.990 2715.140 1197.310 2715.200 ;
        RECT 1089.350 2715.000 1197.310 2715.140 ;
        RECT 1089.350 2714.940 1089.670 2715.000 ;
        RECT 1196.990 2714.940 1197.310 2715.000 ;
        RECT 1200.210 2715.140 1200.530 2715.200 ;
        RECT 1394.330 2715.140 1394.650 2715.200 ;
        RECT 1200.210 2715.000 1394.650 2715.140 ;
        RECT 1200.210 2714.940 1200.530 2715.000 ;
        RECT 1394.330 2714.940 1394.650 2715.000 ;
        RECT 520.790 2714.800 521.110 2714.860 ;
        RECT 688.690 2714.800 689.010 2714.860 ;
        RECT 1020.810 2714.800 1021.130 2714.860 ;
        RECT 520.790 2714.660 689.010 2714.800 ;
        RECT 520.790 2714.600 521.110 2714.660 ;
        RECT 688.690 2714.600 689.010 2714.660 ;
        RECT 699.820 2714.660 1021.130 2714.800 ;
        RECT 351.510 2714.460 351.830 2714.520 ;
        RECT 367.150 2714.460 367.470 2714.520 ;
        RECT 351.510 2714.320 367.470 2714.460 ;
        RECT 351.510 2714.260 351.830 2714.320 ;
        RECT 367.150 2714.260 367.470 2714.320 ;
        RECT 527.690 2714.460 528.010 2714.520 ;
        RECT 699.270 2714.460 699.590 2714.520 ;
        RECT 527.690 2714.320 699.590 2714.460 ;
        RECT 527.690 2714.260 528.010 2714.320 ;
        RECT 699.270 2714.260 699.590 2714.320 ;
        RECT 500.090 2714.120 500.410 2714.180 ;
        RECT 657.410 2714.120 657.730 2714.180 ;
        RECT 500.090 2713.980 657.730 2714.120 ;
        RECT 500.090 2713.920 500.410 2713.980 ;
        RECT 657.410 2713.920 657.730 2713.980 ;
        RECT 665.690 2714.120 666.010 2714.180 ;
        RECT 686.850 2714.120 687.170 2714.180 ;
        RECT 699.820 2714.120 699.960 2714.660 ;
        RECT 1020.810 2714.600 1021.130 2714.660 ;
        RECT 1131.210 2714.800 1131.530 2714.860 ;
        RECT 1280.250 2714.800 1280.570 2714.860 ;
        RECT 1131.210 2714.660 1280.570 2714.800 ;
        RECT 1131.210 2714.600 1131.530 2714.660 ;
        RECT 1280.250 2714.600 1280.570 2714.660 ;
        RECT 700.190 2714.460 700.510 2714.520 ;
        RECT 1000.110 2714.460 1000.430 2714.520 ;
        RECT 700.190 2714.320 1000.430 2714.460 ;
        RECT 700.190 2714.260 700.510 2714.320 ;
        RECT 1000.110 2714.260 1000.430 2714.320 ;
        RECT 1130.750 2714.460 1131.070 2714.520 ;
        RECT 1269.670 2714.460 1269.990 2714.520 ;
        RECT 1130.750 2714.320 1269.990 2714.460 ;
        RECT 1130.750 2714.260 1131.070 2714.320 ;
        RECT 1269.670 2714.260 1269.990 2714.320 ;
        RECT 958.710 2714.120 959.030 2714.180 ;
        RECT 665.690 2713.980 679.260 2714.120 ;
        RECT 665.690 2713.920 666.010 2713.980 ;
        RECT 513.890 2713.780 514.210 2713.840 ;
        RECT 678.570 2713.780 678.890 2713.840 ;
        RECT 513.890 2713.640 678.890 2713.780 ;
        RECT 679.120 2713.780 679.260 2713.980 ;
        RECT 686.850 2713.980 699.960 2714.120 ;
        RECT 700.280 2713.980 959.030 2714.120 ;
        RECT 686.850 2713.920 687.170 2713.980 ;
        RECT 700.280 2713.780 700.420 2713.980 ;
        RECT 958.710 2713.920 959.030 2713.980 ;
        RECT 1117.410 2714.120 1117.730 2714.180 ;
        RECT 1248.970 2714.120 1249.290 2714.180 ;
        RECT 1117.410 2713.980 1249.290 2714.120 ;
        RECT 1117.410 2713.920 1117.730 2713.980 ;
        RECT 1248.970 2713.920 1249.290 2713.980 ;
        RECT 679.120 2713.640 700.420 2713.780 ;
        RECT 700.650 2713.780 700.970 2713.840 ;
        RECT 979.410 2713.780 979.730 2713.840 ;
        RECT 700.650 2713.640 979.730 2713.780 ;
        RECT 513.890 2713.580 514.210 2713.640 ;
        RECT 678.570 2713.580 678.890 2713.640 ;
        RECT 700.650 2713.580 700.970 2713.640 ;
        RECT 979.410 2713.580 979.730 2713.640 ;
        RECT 1124.310 2713.780 1124.630 2713.840 ;
        RECT 1259.550 2713.780 1259.870 2713.840 ;
        RECT 1124.310 2713.640 1259.870 2713.780 ;
        RECT 1124.310 2713.580 1124.630 2713.640 ;
        RECT 1259.550 2713.580 1259.870 2713.640 ;
        RECT 658.790 2713.440 659.110 2713.500 ;
        RECT 927.430 2713.440 927.750 2713.500 ;
        RECT 658.790 2713.300 927.750 2713.440 ;
        RECT 658.790 2713.240 659.110 2713.300 ;
        RECT 927.430 2713.240 927.750 2713.300 ;
        RECT 1110.510 2713.440 1110.830 2713.500 ;
        RECT 1238.850 2713.440 1239.170 2713.500 ;
        RECT 1110.510 2713.300 1239.170 2713.440 ;
        RECT 1110.510 2713.240 1110.830 2713.300 ;
        RECT 1238.850 2713.240 1239.170 2713.300 ;
        RECT 541.490 2713.100 541.810 2713.160 ;
        RECT 730.090 2713.100 730.410 2713.160 ;
        RECT 813.350 2713.100 813.670 2713.160 ;
        RECT 541.490 2712.960 730.410 2713.100 ;
        RECT 541.490 2712.900 541.810 2712.960 ;
        RECT 730.090 2712.900 730.410 2712.960 ;
        RECT 730.640 2712.960 813.670 2713.100 ;
        RECT 325.750 2712.760 326.070 2712.820 ;
        RECT 330.810 2712.760 331.130 2712.820 ;
        RECT 325.750 2712.620 331.130 2712.760 ;
        RECT 325.750 2712.560 326.070 2712.620 ;
        RECT 330.810 2712.560 331.130 2712.620 ;
        RECT 542.410 2712.760 542.730 2712.820 ;
        RECT 719.970 2712.760 720.290 2712.820 ;
        RECT 542.410 2712.620 720.290 2712.760 ;
        RECT 542.410 2712.560 542.730 2712.620 ;
        RECT 719.970 2712.560 720.290 2712.620 ;
        RECT 727.790 2712.760 728.110 2712.820 ;
        RECT 730.640 2712.760 730.780 2712.960 ;
        RECT 813.350 2712.900 813.670 2712.960 ;
        RECT 1103.610 2713.100 1103.930 2713.160 ;
        RECT 1228.270 2713.100 1228.590 2713.160 ;
        RECT 1103.610 2712.960 1228.590 2713.100 ;
        RECT 1103.610 2712.900 1103.930 2712.960 ;
        RECT 1228.270 2712.900 1228.590 2712.960 ;
        RECT 727.790 2712.620 730.780 2712.760 ;
        RECT 741.590 2712.760 741.910 2712.820 ;
        RECT 792.650 2712.760 792.970 2712.820 ;
        RECT 741.590 2712.620 792.970 2712.760 ;
        RECT 727.790 2712.560 728.110 2712.620 ;
        RECT 741.590 2712.560 741.910 2712.620 ;
        RECT 792.650 2712.560 792.970 2712.620 ;
        RECT 1089.810 2712.760 1090.130 2712.820 ;
        RECT 1207.570 2712.760 1207.890 2712.820 ;
        RECT 1089.810 2712.620 1207.890 2712.760 ;
        RECT 1089.810 2712.560 1090.130 2712.620 ;
        RECT 1207.570 2712.560 1207.890 2712.620 ;
        RECT 534.590 2712.420 534.910 2712.480 ;
        RECT 709.390 2712.420 709.710 2712.480 ;
        RECT 771.950 2712.420 772.270 2712.480 ;
        RECT 534.590 2712.280 709.710 2712.420 ;
        RECT 534.590 2712.220 534.910 2712.280 ;
        RECT 709.390 2712.220 709.710 2712.280 ;
        RECT 709.940 2712.280 772.270 2712.420 ;
        RECT 506.990 2712.080 507.310 2712.140 ;
        RECT 667.990 2712.080 668.310 2712.140 ;
        RECT 506.990 2711.940 668.310 2712.080 ;
        RECT 506.990 2711.880 507.310 2711.940 ;
        RECT 667.990 2711.880 668.310 2711.940 ;
        RECT 679.490 2712.080 679.810 2712.140 ;
        RECT 707.090 2712.080 707.410 2712.140 ;
        RECT 709.940 2712.080 710.080 2712.280 ;
        RECT 771.950 2712.220 772.270 2712.280 ;
        RECT 1096.710 2712.420 1097.030 2712.480 ;
        RECT 1217.690 2712.420 1218.010 2712.480 ;
        RECT 1096.710 2712.280 1218.010 2712.420 ;
        RECT 1096.710 2712.220 1097.030 2712.280 ;
        RECT 1217.690 2712.220 1218.010 2712.280 ;
        RECT 750.790 2712.080 751.110 2712.140 ;
        RECT 679.490 2711.940 706.860 2712.080 ;
        RECT 679.490 2711.880 679.810 2711.940 ;
        RECT 706.720 2711.740 706.860 2711.940 ;
        RECT 707.090 2711.940 710.080 2712.080 ;
        RECT 710.400 2711.940 751.110 2712.080 ;
        RECT 707.090 2711.880 707.410 2711.940 ;
        RECT 710.400 2711.740 710.540 2711.940 ;
        RECT 750.790 2711.880 751.110 2711.940 ;
        RECT 706.720 2711.600 710.540 2711.740 ;
      LAYER met1 ;
        RECT 300.070 1604.460 1395.190 2695.780 ;
      LAYER met1 ;
        RECT 1407.670 2145.980 1407.990 2146.040 ;
        RECT 1835.470 2145.980 1835.790 2146.040 ;
        RECT 1407.670 2145.840 1835.790 2145.980 ;
        RECT 1407.670 2145.780 1407.990 2145.840 ;
        RECT 1835.470 2145.780 1835.790 2145.840 ;
        RECT 1407.670 2139.180 1407.990 2139.240 ;
        RECT 1842.370 2139.180 1842.690 2139.240 ;
        RECT 1407.670 2139.040 1842.690 2139.180 ;
        RECT 1407.670 2138.980 1407.990 2139.040 ;
        RECT 1842.370 2138.980 1842.690 2139.040 ;
        RECT 1408.130 2132.720 1408.450 2132.780 ;
        RECT 1849.270 2132.720 1849.590 2132.780 ;
        RECT 1408.130 2132.580 1849.590 2132.720 ;
        RECT 1408.130 2132.520 1408.450 2132.580 ;
        RECT 1849.270 2132.520 1849.590 2132.580 ;
        RECT 1407.670 2132.380 1407.990 2132.440 ;
        RECT 1856.170 2132.380 1856.490 2132.440 ;
        RECT 1407.670 2132.240 1856.490 2132.380 ;
        RECT 1407.670 2132.180 1407.990 2132.240 ;
        RECT 1856.170 2132.180 1856.490 2132.240 ;
        RECT 1407.670 2125.580 1407.990 2125.640 ;
        RECT 1863.070 2125.580 1863.390 2125.640 ;
        RECT 1407.670 2125.440 1863.390 2125.580 ;
        RECT 1407.670 2125.380 1407.990 2125.440 ;
        RECT 1863.070 2125.380 1863.390 2125.440 ;
        RECT 1407.670 2118.440 1407.990 2118.500 ;
        RECT 1869.970 2118.440 1870.290 2118.500 ;
        RECT 1407.670 2118.300 1870.290 2118.440 ;
        RECT 1407.670 2118.240 1407.990 2118.300 ;
        RECT 1869.970 2118.240 1870.290 2118.300 ;
        RECT 1408.130 2111.980 1408.450 2112.040 ;
        RECT 1870.430 2111.980 1870.750 2112.040 ;
        RECT 1408.130 2111.840 1870.750 2111.980 ;
        RECT 1408.130 2111.780 1408.450 2111.840 ;
        RECT 1870.430 2111.780 1870.750 2111.840 ;
        RECT 1407.670 2111.640 1407.990 2111.700 ;
        RECT 1876.870 2111.640 1877.190 2111.700 ;
        RECT 1407.670 2111.500 1877.190 2111.640 ;
        RECT 1407.670 2111.440 1407.990 2111.500 ;
        RECT 1876.870 2111.440 1877.190 2111.500 ;
        RECT 1407.670 2104.840 1407.990 2104.900 ;
        RECT 1883.770 2104.840 1884.090 2104.900 ;
        RECT 1407.670 2104.700 1884.090 2104.840 ;
        RECT 1407.670 2104.640 1407.990 2104.700 ;
        RECT 1883.770 2104.640 1884.090 2104.700 ;
        RECT 1407.670 2097.700 1407.990 2097.760 ;
        RECT 1890.670 2097.700 1890.990 2097.760 ;
        RECT 1407.670 2097.560 1890.990 2097.700 ;
        RECT 1407.670 2097.500 1407.990 2097.560 ;
        RECT 1890.670 2097.500 1890.990 2097.560 ;
        RECT 1408.130 2091.240 1408.450 2091.300 ;
        RECT 1897.570 2091.240 1897.890 2091.300 ;
        RECT 1408.130 2091.100 1897.890 2091.240 ;
        RECT 1408.130 2091.040 1408.450 2091.100 ;
        RECT 1897.570 2091.040 1897.890 2091.100 ;
        RECT 1407.670 2090.900 1407.990 2090.960 ;
        RECT 1904.470 2090.900 1904.790 2090.960 ;
        RECT 1407.670 2090.760 1904.790 2090.900 ;
        RECT 1407.670 2090.700 1407.990 2090.760 ;
        RECT 1904.470 2090.700 1904.790 2090.760 ;
        RECT 1414.110 2084.100 1414.430 2084.160 ;
        RECT 1911.370 2084.100 1911.690 2084.160 ;
        RECT 1414.110 2083.960 1911.690 2084.100 ;
        RECT 1414.110 2083.900 1414.430 2083.960 ;
        RECT 1911.370 2083.900 1911.690 2083.960 ;
        RECT 1411.350 2077.300 1411.670 2077.360 ;
        RECT 1911.830 2077.300 1912.150 2077.360 ;
        RECT 1411.350 2077.160 1912.150 2077.300 ;
        RECT 1411.350 2077.100 1411.670 2077.160 ;
        RECT 1911.830 2077.100 1912.150 2077.160 ;
        RECT 1408.590 2070.500 1408.910 2070.560 ;
        RECT 1919.190 2070.500 1919.510 2070.560 ;
        RECT 1408.590 2070.360 1919.510 2070.500 ;
        RECT 1408.590 2070.300 1408.910 2070.360 ;
        RECT 1919.190 2070.300 1919.510 2070.360 ;
        RECT 1410.430 2070.160 1410.750 2070.220 ;
        RECT 1925.170 2070.160 1925.490 2070.220 ;
        RECT 1410.430 2070.020 1925.490 2070.160 ;
        RECT 1410.430 2069.960 1410.750 2070.020 ;
        RECT 1925.170 2069.960 1925.490 2070.020 ;
        RECT 1917.810 2069.480 1918.130 2069.540 ;
        RECT 1965.650 2069.480 1965.970 2069.540 ;
        RECT 1917.810 2069.340 1965.970 2069.480 ;
        RECT 1917.810 2069.280 1918.130 2069.340 ;
        RECT 1965.650 2069.280 1965.970 2069.340 ;
        RECT 1629.390 2069.140 1629.710 2069.200 ;
        RECT 1675.850 2069.140 1676.170 2069.200 ;
        RECT 1629.390 2069.000 1676.170 2069.140 ;
        RECT 1629.390 2068.940 1629.710 2069.000 ;
        RECT 1675.850 2068.940 1676.170 2069.000 ;
        RECT 1725.990 2069.140 1726.310 2069.200 ;
        RECT 1772.450 2069.140 1772.770 2069.200 ;
        RECT 1725.990 2069.000 1772.770 2069.140 ;
        RECT 1725.990 2068.940 1726.310 2069.000 ;
        RECT 1772.450 2068.940 1772.770 2069.000 ;
        RECT 1890.210 2069.140 1890.530 2069.200 ;
        RECT 1936.670 2069.140 1936.990 2069.200 ;
        RECT 1980.370 2069.140 1980.690 2069.200 ;
        RECT 1890.210 2069.000 1980.690 2069.140 ;
        RECT 1890.210 2068.940 1890.530 2069.000 ;
        RECT 1936.670 2068.940 1936.990 2069.000 ;
        RECT 1980.370 2068.940 1980.690 2069.000 ;
        RECT 1628.930 2068.800 1629.250 2068.860 ;
        RECT 1676.310 2068.800 1676.630 2068.860 ;
        RECT 1628.930 2068.660 1676.630 2068.800 ;
        RECT 1628.930 2068.600 1629.250 2068.660 ;
        RECT 1676.310 2068.600 1676.630 2068.660 ;
        RECT 1725.530 2068.800 1725.850 2068.860 ;
        RECT 1772.910 2068.800 1773.230 2068.860 ;
        RECT 1725.530 2068.660 1773.230 2068.800 ;
        RECT 1725.530 2068.600 1725.850 2068.660 ;
        RECT 1772.910 2068.600 1773.230 2068.660 ;
        RECT 1848.810 2068.800 1849.130 2068.860 ;
        RECT 1893.890 2068.800 1894.210 2068.860 ;
        RECT 1941.730 2068.800 1942.050 2068.860 ;
        RECT 1987.270 2068.800 1987.590 2068.860 ;
        RECT 1848.810 2068.660 1987.590 2068.800 ;
        RECT 1848.810 2068.600 1849.130 2068.660 ;
        RECT 1893.890 2068.600 1894.210 2068.660 ;
        RECT 1941.730 2068.600 1942.050 2068.660 ;
        RECT 1987.270 2068.600 1987.590 2068.660 ;
        RECT 1413.190 2068.460 1413.510 2068.520 ;
        RECT 1841.450 2068.460 1841.770 2068.520 ;
        RECT 1890.210 2068.460 1890.530 2068.520 ;
        RECT 1413.190 2068.320 1890.530 2068.460 ;
        RECT 1413.190 2068.260 1413.510 2068.320 ;
        RECT 1841.450 2068.260 1841.770 2068.320 ;
        RECT 1890.210 2068.260 1890.530 2068.320 ;
        RECT 1930.230 2068.460 1930.550 2068.520 ;
        RECT 1973.470 2068.460 1973.790 2068.520 ;
        RECT 1930.230 2068.320 1973.790 2068.460 ;
        RECT 1930.230 2068.260 1930.550 2068.320 ;
        RECT 1973.470 2068.260 1973.790 2068.320 ;
        RECT 1407.670 2068.120 1407.990 2068.180 ;
        RECT 1843.750 2068.120 1844.070 2068.180 ;
        RECT 1407.670 2067.980 1844.070 2068.120 ;
        RECT 1407.670 2067.920 1407.990 2067.980 ;
        RECT 1843.750 2067.920 1844.070 2067.980 ;
        RECT 1844.210 2068.120 1844.530 2068.180 ;
        RECT 1849.270 2068.120 1849.590 2068.180 ;
        RECT 1898.030 2068.120 1898.350 2068.180 ;
        RECT 1948.170 2068.120 1948.490 2068.180 ;
        RECT 1844.210 2067.980 1948.490 2068.120 ;
        RECT 1844.210 2067.920 1844.530 2067.980 ;
        RECT 1849.270 2067.920 1849.590 2067.980 ;
        RECT 1898.030 2067.920 1898.350 2067.980 ;
        RECT 1948.170 2067.920 1948.490 2067.980 ;
        RECT 1591.210 2067.780 1591.530 2067.840 ;
        RECT 2028.670 2067.780 2028.990 2067.840 ;
        RECT 1591.210 2067.640 2028.990 2067.780 ;
        RECT 1591.210 2067.580 1591.530 2067.640 ;
        RECT 2028.670 2067.580 2028.990 2067.640 ;
        RECT 1409.050 2067.440 1409.370 2067.500 ;
        RECT 1844.210 2067.440 1844.530 2067.500 ;
        RECT 1409.050 2067.300 1844.530 2067.440 ;
        RECT 1409.050 2067.240 1409.370 2067.300 ;
        RECT 1844.210 2067.240 1844.530 2067.300 ;
        RECT 1844.670 2067.440 1844.990 2067.500 ;
        RECT 1864.910 2067.440 1865.230 2067.500 ;
        RECT 1911.370 2067.440 1911.690 2067.500 ;
        RECT 1844.670 2067.300 1911.690 2067.440 ;
        RECT 1844.670 2067.240 1844.990 2067.300 ;
        RECT 1864.910 2067.240 1865.230 2067.300 ;
        RECT 1911.370 2067.240 1911.690 2067.300 ;
        RECT 1924.710 2067.440 1925.030 2067.500 ;
        RECT 1969.790 2067.440 1970.110 2067.500 ;
        RECT 1924.710 2067.300 1970.110 2067.440 ;
        RECT 1924.710 2067.240 1925.030 2067.300 ;
        RECT 1969.790 2067.240 1970.110 2067.300 ;
        RECT 1973.470 2067.440 1973.790 2067.500 ;
        RECT 1976.690 2067.440 1977.010 2067.500 ;
        RECT 2021.770 2067.440 2022.090 2067.500 ;
        RECT 1973.470 2067.300 2022.090 2067.440 ;
        RECT 1973.470 2067.240 1973.790 2067.300 ;
        RECT 1976.690 2067.240 1977.010 2067.300 ;
        RECT 2021.770 2067.240 2022.090 2067.300 ;
        RECT 1435.730 2067.100 1436.050 2067.160 ;
        RECT 1482.650 2067.100 1482.970 2067.160 ;
        RECT 1435.730 2066.960 1482.970 2067.100 ;
        RECT 1435.730 2066.900 1436.050 2066.960 ;
        RECT 1482.650 2066.900 1482.970 2066.960 ;
        RECT 1532.330 2067.100 1532.650 2067.160 ;
        RECT 1579.250 2067.100 1579.570 2067.160 ;
        RECT 1532.330 2066.960 1579.570 2067.100 ;
        RECT 1532.330 2066.900 1532.650 2066.960 ;
        RECT 1579.250 2066.900 1579.570 2066.960 ;
        RECT 1590.750 2067.100 1591.070 2067.160 ;
        RECT 2035.570 2067.100 2035.890 2067.160 ;
        RECT 1590.750 2066.960 2035.890 2067.100 ;
        RECT 1590.750 2066.900 1591.070 2066.960 ;
        RECT 2035.570 2066.900 2035.890 2066.960 ;
        RECT 1410.890 2066.760 1411.210 2066.820 ;
        RECT 1859.850 2066.760 1860.170 2066.820 ;
        RECT 1907.690 2066.760 1908.010 2066.820 ;
        RECT 1954.610 2066.760 1954.930 2066.820 ;
        RECT 1959.210 2066.760 1959.530 2066.820 ;
        RECT 1410.890 2066.620 1959.530 2066.760 ;
        RECT 1410.890 2066.560 1411.210 2066.620 ;
        RECT 1859.850 2066.560 1860.170 2066.620 ;
        RECT 1907.690 2066.560 1908.010 2066.620 ;
        RECT 1954.610 2066.560 1954.930 2066.620 ;
        RECT 1959.210 2066.560 1959.530 2066.620 ;
        RECT 1965.650 2066.760 1965.970 2066.820 ;
        RECT 2007.970 2066.760 2008.290 2066.820 ;
        RECT 1965.650 2066.620 2008.290 2066.760 ;
        RECT 1965.650 2066.560 1965.970 2066.620 ;
        RECT 2007.970 2066.560 2008.290 2066.620 ;
        RECT 1414.110 2066.420 1414.430 2066.480 ;
        RECT 1932.070 2066.420 1932.390 2066.480 ;
        RECT 1414.110 2066.280 1932.390 2066.420 ;
        RECT 1414.110 2066.220 1414.430 2066.280 ;
        RECT 1932.070 2066.220 1932.390 2066.280 ;
        RECT 1969.790 2066.420 1970.110 2066.480 ;
        RECT 2015.790 2066.420 2016.110 2066.480 ;
        RECT 1969.790 2066.280 2016.110 2066.420 ;
        RECT 1969.790 2066.220 1970.110 2066.280 ;
        RECT 2015.790 2066.220 2016.110 2066.280 ;
        RECT 1435.270 2066.080 1435.590 2066.140 ;
        RECT 1483.110 2066.080 1483.430 2066.140 ;
        RECT 1435.270 2065.940 1483.430 2066.080 ;
        RECT 1435.270 2065.880 1435.590 2065.940 ;
        RECT 1483.110 2065.880 1483.430 2065.940 ;
        RECT 1531.870 2066.080 1532.190 2066.140 ;
        RECT 1579.710 2066.080 1580.030 2066.140 ;
        RECT 1531.870 2065.940 1580.030 2066.080 ;
        RECT 1531.870 2065.880 1532.190 2065.940 ;
        RECT 1579.710 2065.880 1580.030 2065.940 ;
        RECT 1590.290 2066.080 1590.610 2066.140 ;
        RECT 2042.470 2066.080 2042.790 2066.140 ;
        RECT 1590.290 2065.940 2042.790 2066.080 ;
        RECT 1590.290 2065.880 1590.610 2065.940 ;
        RECT 2042.470 2065.880 2042.790 2065.940 ;
        RECT 1411.810 2065.740 1412.130 2065.800 ;
        RECT 1844.670 2065.740 1844.990 2065.800 ;
        RECT 1911.370 2065.740 1911.690 2065.800 ;
        RECT 1958.750 2065.740 1959.070 2065.800 ;
        RECT 1411.810 2065.600 1844.990 2065.740 ;
        RECT 1411.810 2065.540 1412.130 2065.600 ;
        RECT 1844.670 2065.540 1844.990 2065.600 ;
        RECT 1845.220 2065.600 1846.740 2065.740 ;
        RECT 1409.970 2065.400 1410.290 2065.460 ;
        RECT 1435.730 2065.400 1436.050 2065.460 ;
        RECT 1409.970 2065.260 1436.050 2065.400 ;
        RECT 1409.970 2065.200 1410.290 2065.260 ;
        RECT 1435.730 2065.200 1436.050 2065.260 ;
        RECT 1482.650 2065.400 1482.970 2065.460 ;
        RECT 1532.330 2065.400 1532.650 2065.460 ;
        RECT 1482.650 2065.260 1532.650 2065.400 ;
        RECT 1482.650 2065.200 1482.970 2065.260 ;
        RECT 1532.330 2065.200 1532.650 2065.260 ;
        RECT 1579.250 2065.400 1579.570 2065.460 ;
        RECT 1629.390 2065.400 1629.710 2065.460 ;
        RECT 1579.250 2065.260 1629.710 2065.400 ;
        RECT 1579.250 2065.200 1579.570 2065.260 ;
        RECT 1629.390 2065.200 1629.710 2065.260 ;
        RECT 1675.850 2065.400 1676.170 2065.460 ;
        RECT 1725.990 2065.400 1726.310 2065.460 ;
        RECT 1675.850 2065.260 1726.310 2065.400 ;
        RECT 1675.850 2065.200 1676.170 2065.260 ;
        RECT 1725.990 2065.200 1726.310 2065.260 ;
        RECT 1772.450 2065.400 1772.770 2065.460 ;
        RECT 1844.210 2065.400 1844.530 2065.460 ;
        RECT 1772.450 2065.260 1844.530 2065.400 ;
        RECT 1772.450 2065.200 1772.770 2065.260 ;
        RECT 1844.210 2065.200 1844.530 2065.260 ;
        RECT 1412.270 2065.060 1412.590 2065.120 ;
        RECT 1435.270 2065.060 1435.590 2065.120 ;
        RECT 1412.270 2064.920 1435.590 2065.060 ;
        RECT 1412.270 2064.860 1412.590 2064.920 ;
        RECT 1435.270 2064.860 1435.590 2064.920 ;
        RECT 1483.110 2065.060 1483.430 2065.120 ;
        RECT 1531.870 2065.060 1532.190 2065.120 ;
        RECT 1483.110 2064.920 1532.190 2065.060 ;
        RECT 1483.110 2064.860 1483.430 2064.920 ;
        RECT 1531.870 2064.860 1532.190 2064.920 ;
        RECT 1579.710 2065.060 1580.030 2065.120 ;
        RECT 1628.930 2065.060 1629.250 2065.120 ;
        RECT 1579.710 2064.920 1629.250 2065.060 ;
        RECT 1579.710 2064.860 1580.030 2064.920 ;
        RECT 1628.930 2064.860 1629.250 2064.920 ;
        RECT 1676.310 2065.060 1676.630 2065.120 ;
        RECT 1725.530 2065.060 1725.850 2065.120 ;
        RECT 1676.310 2064.920 1725.850 2065.060 ;
        RECT 1676.310 2064.860 1676.630 2064.920 ;
        RECT 1725.530 2064.860 1725.850 2064.920 ;
        RECT 1772.910 2065.060 1773.230 2065.120 ;
        RECT 1845.220 2065.060 1845.360 2065.600 ;
        RECT 1846.600 2065.400 1846.740 2065.600 ;
        RECT 1911.370 2065.600 1959.070 2065.740 ;
        RECT 1911.370 2065.540 1911.690 2065.600 ;
        RECT 1958.750 2065.540 1959.070 2065.600 ;
        RECT 1959.210 2065.740 1959.530 2065.800 ;
        RECT 1994.170 2065.740 1994.490 2065.800 ;
        RECT 1959.210 2065.600 1994.490 2065.740 ;
        RECT 1959.210 2065.540 1959.530 2065.600 ;
        RECT 1994.170 2065.540 1994.490 2065.600 ;
        RECT 1877.330 2065.400 1877.650 2065.460 ;
        RECT 1958.840 2065.400 1958.980 2065.540 ;
        RECT 2001.070 2065.400 2001.390 2065.460 ;
        RECT 1846.600 2065.260 1918.040 2065.400 ;
        RECT 1958.840 2065.260 2001.390 2065.400 ;
        RECT 1877.330 2065.200 1877.650 2065.260 ;
        RECT 1772.910 2064.920 1845.360 2065.060 ;
        RECT 1846.510 2065.060 1846.830 2065.120 ;
        RECT 1871.810 2065.060 1872.130 2065.120 ;
        RECT 1917.350 2065.060 1917.670 2065.120 ;
        RECT 1846.510 2064.920 1917.670 2065.060 ;
        RECT 1917.900 2065.060 1918.040 2065.260 ;
        RECT 2001.070 2065.200 2001.390 2065.260 ;
        RECT 1924.710 2065.060 1925.030 2065.120 ;
        RECT 1917.900 2064.920 1925.030 2065.060 ;
        RECT 1772.910 2064.860 1773.230 2064.920 ;
        RECT 1846.510 2064.860 1846.830 2064.920 ;
        RECT 1871.810 2064.860 1872.130 2064.920 ;
        RECT 1917.350 2064.860 1917.670 2064.920 ;
        RECT 1924.710 2064.860 1925.030 2064.920 ;
        RECT 1411.350 2064.720 1411.670 2064.780 ;
        RECT 1882.850 2064.720 1883.170 2064.780 ;
        RECT 1930.230 2064.720 1930.550 2064.780 ;
        RECT 1411.350 2064.580 1930.550 2064.720 ;
        RECT 1411.350 2064.520 1411.670 2064.580 ;
        RECT 1882.850 2064.520 1883.170 2064.580 ;
        RECT 1930.230 2064.520 1930.550 2064.580 ;
        RECT 1948.170 2064.720 1948.490 2064.780 ;
        RECT 1987.270 2064.720 1987.590 2064.780 ;
        RECT 1948.170 2064.580 1987.590 2064.720 ;
        RECT 1948.170 2064.520 1948.490 2064.580 ;
        RECT 1987.270 2064.520 1987.590 2064.580 ;
        RECT 1413.650 2064.380 1413.970 2064.440 ;
        RECT 1966.570 2064.380 1966.890 2064.440 ;
        RECT 1413.650 2064.240 1966.890 2064.380 ;
        RECT 1413.650 2064.180 1413.970 2064.240 ;
        RECT 1966.570 2064.180 1966.890 2064.240 ;
        RECT 1410.430 2064.040 1410.750 2064.100 ;
        RECT 1973.470 2064.040 1973.790 2064.100 ;
        RECT 1410.430 2063.900 1973.790 2064.040 ;
        RECT 1410.430 2063.840 1410.750 2063.900 ;
        RECT 1973.470 2063.840 1973.790 2063.900 ;
        RECT 1407.670 2063.500 1407.990 2063.760 ;
        RECT 1408.130 2063.700 1408.450 2063.760 ;
        RECT 1980.370 2063.700 1980.690 2063.760 ;
        RECT 1408.130 2063.560 1980.690 2063.700 ;
        RECT 1408.130 2063.500 1408.450 2063.560 ;
        RECT 1980.370 2063.500 1980.690 2063.560 ;
        RECT 1407.760 2063.360 1407.900 2063.500 ;
        RECT 2028.670 2063.360 2028.990 2063.420 ;
        RECT 1407.760 2063.220 2028.990 2063.360 ;
        RECT 2028.670 2063.160 2028.990 2063.220 ;
        RECT 1407.670 2062.820 1407.990 2063.080 ;
        RECT 1407.760 2061.720 1407.900 2062.820 ;
        RECT 1409.050 2062.480 1409.370 2062.740 ;
        RECT 1409.140 2062.340 1409.280 2062.480 ;
        RECT 1413.650 2062.340 1413.970 2062.400 ;
        RECT 1409.140 2062.200 1413.970 2062.340 ;
        RECT 1413.650 2062.140 1413.970 2062.200 ;
        RECT 1409.050 2062.000 1409.370 2062.060 ;
        RECT 1410.430 2062.000 1410.750 2062.060 ;
        RECT 1409.050 2061.860 1410.750 2062.000 ;
        RECT 1409.050 2061.800 1409.370 2061.860 ;
        RECT 1410.430 2061.800 1410.750 2061.860 ;
        RECT 1420.550 2062.000 1420.870 2062.060 ;
        RECT 1718.630 2062.000 1718.950 2062.060 ;
        RECT 1420.550 2061.860 1718.950 2062.000 ;
        RECT 1420.550 2061.800 1420.870 2061.860 ;
        RECT 1718.630 2061.800 1718.950 2061.860 ;
        RECT 1407.670 2061.460 1407.990 2061.720 ;
        RECT 1420.090 2061.660 1420.410 2061.720 ;
        RECT 1718.170 2061.660 1718.490 2061.720 ;
        RECT 1420.090 2061.520 1718.490 2061.660 ;
        RECT 1420.090 2061.460 1420.410 2061.520 ;
        RECT 1718.170 2061.460 1718.490 2061.520 ;
        RECT 1421.010 2061.320 1421.330 2061.380 ;
        RECT 1725.070 2061.320 1725.390 2061.380 ;
        RECT 1421.010 2061.180 1725.390 2061.320 ;
        RECT 1421.010 2061.120 1421.330 2061.180 ;
        RECT 1725.070 2061.120 1725.390 2061.180 ;
        RECT 1417.330 2060.980 1417.650 2061.040 ;
        RECT 1731.970 2060.980 1732.290 2061.040 ;
        RECT 1417.330 2060.840 1732.290 2060.980 ;
        RECT 1417.330 2060.780 1417.650 2060.840 ;
        RECT 1731.970 2060.780 1732.290 2060.840 ;
        RECT 1416.870 2060.640 1417.190 2060.700 ;
        RECT 1738.870 2060.640 1739.190 2060.700 ;
        RECT 1416.870 2060.500 1739.190 2060.640 ;
        RECT 1416.870 2060.440 1417.190 2060.500 ;
        RECT 1738.870 2060.440 1739.190 2060.500 ;
        RECT 1414.570 2060.300 1414.890 2060.360 ;
        RECT 1745.770 2060.300 1746.090 2060.360 ;
        RECT 1414.570 2060.160 1746.090 2060.300 ;
        RECT 1414.570 2060.100 1414.890 2060.160 ;
        RECT 1745.770 2060.100 1746.090 2060.160 ;
        RECT 1409.510 2059.960 1409.830 2060.020 ;
        RECT 1753.130 2059.960 1753.450 2060.020 ;
        RECT 1409.510 2059.820 1753.450 2059.960 ;
        RECT 1409.510 2059.760 1409.830 2059.820 ;
        RECT 1753.130 2059.760 1753.450 2059.820 ;
        RECT 1528.190 2059.620 1528.510 2059.680 ;
        RECT 2097.670 2059.620 2097.990 2059.680 ;
        RECT 1528.190 2059.480 2097.990 2059.620 ;
        RECT 1528.190 2059.420 1528.510 2059.480 ;
        RECT 2097.670 2059.420 2097.990 2059.480 ;
        RECT 1555.790 2059.280 1556.110 2059.340 ;
        RECT 1987.270 2059.280 1987.590 2059.340 ;
        RECT 1555.790 2059.140 1987.590 2059.280 ;
        RECT 1555.790 2059.080 1556.110 2059.140 ;
        RECT 1987.270 2059.080 1987.590 2059.140 ;
        RECT 1410.430 2058.940 1410.750 2059.000 ;
        RECT 1940.350 2058.940 1940.670 2059.000 ;
        RECT 1410.430 2058.800 1940.670 2058.940 ;
        RECT 1410.430 2058.740 1410.750 2058.800 ;
        RECT 1940.350 2058.740 1940.670 2058.800 ;
        RECT 1415.030 2058.600 1415.350 2058.660 ;
        RECT 1955.070 2058.600 1955.390 2058.660 ;
        RECT 1415.030 2058.460 1955.390 2058.600 ;
        RECT 1415.030 2058.400 1415.350 2058.460 ;
        RECT 1955.070 2058.400 1955.390 2058.460 ;
        RECT 1425.150 2058.260 1425.470 2058.320 ;
        RECT 1995.550 2058.260 1995.870 2058.320 ;
        RECT 1425.150 2058.120 1995.870 2058.260 ;
        RECT 1425.150 2058.060 1425.470 2058.120 ;
        RECT 1995.550 2058.060 1995.870 2058.120 ;
        RECT 1410.430 2057.920 1410.750 2057.980 ;
        RECT 1990.030 2057.920 1990.350 2057.980 ;
        RECT 1410.430 2057.780 1990.350 2057.920 ;
        RECT 1410.430 2057.720 1410.750 2057.780 ;
        RECT 1990.030 2057.720 1990.350 2057.780 ;
        RECT 1415.490 2057.580 1415.810 2057.640 ;
        RECT 2004.750 2057.580 2005.070 2057.640 ;
        RECT 1415.490 2057.440 2005.070 2057.580 ;
        RECT 1415.490 2057.380 1415.810 2057.440 ;
        RECT 2004.750 2057.380 2005.070 2057.440 ;
        RECT 1416.410 2057.240 1416.730 2057.300 ;
        RECT 2008.430 2057.240 2008.750 2057.300 ;
        RECT 1416.410 2057.100 2008.750 2057.240 ;
        RECT 1416.410 2057.040 1416.730 2057.100 ;
        RECT 2008.430 2057.040 2008.750 2057.100 ;
        RECT 1412.270 2056.900 1412.590 2056.960 ;
        RECT 1414.110 2056.900 1414.430 2056.960 ;
        RECT 1412.270 2056.760 1414.430 2056.900 ;
        RECT 1412.270 2056.700 1412.590 2056.760 ;
        RECT 1414.110 2056.700 1414.430 2056.760 ;
        RECT 1424.690 2056.900 1425.010 2056.960 ;
        RECT 2021.770 2056.900 2022.090 2056.960 ;
        RECT 1424.690 2056.760 2022.090 2056.900 ;
        RECT 1424.690 2056.700 1425.010 2056.760 ;
        RECT 2021.770 2056.700 2022.090 2056.760 ;
        RECT 1409.510 2056.560 1409.830 2056.620 ;
        RECT 1409.140 2056.420 1409.830 2056.560 ;
        RECT 1409.140 2050.780 1409.280 2056.420 ;
        RECT 1409.510 2056.360 1409.830 2056.420 ;
        RECT 1415.950 2056.560 1416.270 2056.620 ;
        RECT 2016.250 2056.560 2016.570 2056.620 ;
        RECT 1415.950 2056.420 2016.570 2056.560 ;
        RECT 1415.950 2056.360 1416.270 2056.420 ;
        RECT 2016.250 2056.360 2016.570 2056.420 ;
        RECT 1414.110 2056.220 1414.430 2056.280 ;
        RECT 1946.330 2056.220 1946.650 2056.280 ;
        RECT 1414.110 2056.080 1946.650 2056.220 ;
        RECT 1414.110 2056.020 1414.430 2056.080 ;
        RECT 1946.330 2056.020 1946.650 2056.080 ;
        RECT 1409.510 2055.880 1409.830 2055.940 ;
        RECT 1948.630 2055.880 1948.950 2055.940 ;
        RECT 1409.510 2055.740 1948.950 2055.880 ;
        RECT 1409.510 2055.680 1409.830 2055.740 ;
        RECT 1948.630 2055.680 1948.950 2055.740 ;
        RECT 1493.690 2053.840 1494.010 2053.900 ;
        RECT 1711.270 2053.840 1711.590 2053.900 ;
        RECT 1493.690 2053.700 1711.590 2053.840 ;
        RECT 1493.690 2053.640 1494.010 2053.700 ;
        RECT 1711.270 2053.640 1711.590 2053.700 ;
        RECT 1419.630 2053.500 1419.950 2053.560 ;
        RECT 1704.370 2053.500 1704.690 2053.560 ;
        RECT 1419.630 2053.360 1704.690 2053.500 ;
        RECT 1419.630 2053.300 1419.950 2053.360 ;
        RECT 1704.370 2053.300 1704.690 2053.360 ;
        RECT 1414.570 2053.160 1414.890 2053.220 ;
        RECT 1961.510 2053.160 1961.830 2053.220 ;
        RECT 1414.570 2053.020 1961.830 2053.160 ;
        RECT 1414.570 2052.960 1414.890 2053.020 ;
        RECT 1961.510 2052.960 1961.830 2053.020 ;
        RECT 1419.170 2052.820 1419.490 2052.880 ;
        RECT 2049.830 2052.820 2050.150 2052.880 ;
        RECT 1419.170 2052.680 2050.150 2052.820 ;
        RECT 1419.170 2052.620 1419.490 2052.680 ;
        RECT 2049.830 2052.620 2050.150 2052.680 ;
        RECT 1409.510 2050.780 1409.830 2050.840 ;
        RECT 1409.140 2050.640 1409.830 2050.780 ;
        RECT 1409.510 2050.580 1409.830 2050.640 ;
        RECT 1410.430 2039.360 1410.750 2039.620 ;
        RECT 1410.890 2039.560 1411.210 2039.620 ;
        RECT 1413.190 2039.560 1413.510 2039.620 ;
        RECT 1410.890 2039.420 1413.510 2039.560 ;
        RECT 1410.890 2039.360 1411.210 2039.420 ;
        RECT 1413.190 2039.360 1413.510 2039.420 ;
        RECT 1408.130 2039.220 1408.450 2039.280 ;
        RECT 1408.130 2039.080 1410.200 2039.220 ;
        RECT 1408.130 2039.020 1408.450 2039.080 ;
        RECT 1410.060 2038.600 1410.200 2039.080 ;
        RECT 1408.130 2038.540 1408.450 2038.600 ;
        RECT 1409.510 2038.540 1409.830 2038.600 ;
        RECT 1408.130 2038.400 1409.830 2038.540 ;
        RECT 1408.130 2038.340 1408.450 2038.400 ;
        RECT 1409.510 2038.340 1409.830 2038.400 ;
        RECT 1409.970 2038.340 1410.290 2038.600 ;
        RECT 1410.520 2038.200 1410.660 2039.360 ;
        RECT 1409.600 2038.060 1410.660 2038.200 ;
        RECT 1409.600 2037.920 1409.740 2038.060 ;
        RECT 1409.510 2037.660 1409.830 2037.920 ;
        RECT 1409.970 2037.860 1410.290 2037.920 ;
        RECT 1413.650 2037.860 1413.970 2037.920 ;
        RECT 1409.970 2037.720 1413.970 2037.860 ;
        RECT 1409.970 2037.660 1410.290 2037.720 ;
        RECT 1413.650 2037.660 1413.970 2037.720 ;
        RECT 1414.110 2021.540 1414.430 2021.600 ;
        RECT 1555.790 2021.540 1556.110 2021.600 ;
        RECT 1414.110 2021.400 1556.110 2021.540 ;
        RECT 1414.110 2021.340 1414.430 2021.400 ;
        RECT 1555.790 2021.340 1556.110 2021.400 ;
        RECT 1411.350 2014.200 1411.670 2014.460 ;
        RECT 1411.440 2013.440 1411.580 2014.200 ;
        RECT 1411.350 2013.180 1411.670 2013.440 ;
        RECT 1410.890 2013.040 1411.210 2013.100 ;
        RECT 1425.150 2013.040 1425.470 2013.100 ;
        RECT 1410.890 2012.900 1425.470 2013.040 ;
        RECT 1410.890 2012.840 1411.210 2012.900 ;
        RECT 1425.150 2012.840 1425.470 2012.900 ;
        RECT 1408.130 2005.900 1408.450 2005.960 ;
        RECT 1415.490 2005.900 1415.810 2005.960 ;
        RECT 1408.130 2005.760 1415.810 2005.900 ;
        RECT 1408.130 2005.700 1408.450 2005.760 ;
        RECT 1415.490 2005.700 1415.810 2005.760 ;
        RECT 1408.130 2000.800 1408.450 2000.860 ;
        RECT 1416.410 2000.800 1416.730 2000.860 ;
        RECT 1408.130 2000.660 1416.730 2000.800 ;
        RECT 1408.130 2000.600 1408.450 2000.660 ;
        RECT 1416.410 2000.600 1416.730 2000.660 ;
        RECT 1408.130 1997.740 1408.450 1997.800 ;
        RECT 1415.950 1997.740 1416.270 1997.800 ;
        RECT 1408.130 1997.600 1416.270 1997.740 ;
        RECT 1408.130 1997.540 1408.450 1997.600 ;
        RECT 1415.950 1997.540 1416.270 1997.600 ;
        RECT 1410.890 1990.940 1411.210 1991.000 ;
        RECT 1424.690 1990.940 1425.010 1991.000 ;
        RECT 1410.890 1990.800 1425.010 1990.940 ;
        RECT 1410.890 1990.740 1411.210 1990.800 ;
        RECT 1424.690 1990.740 1425.010 1990.800 ;
        RECT 1408.130 1972.920 1408.450 1972.980 ;
        RECT 1418.710 1972.920 1419.030 1972.980 ;
        RECT 1408.130 1972.780 1419.030 1972.920 ;
        RECT 1408.130 1972.720 1408.450 1972.780 ;
        RECT 1418.710 1972.720 1419.030 1972.780 ;
        RECT 1410.890 1966.460 1411.210 1966.520 ;
        RECT 1412.730 1966.460 1413.050 1966.520 ;
        RECT 1410.890 1966.320 1413.050 1966.460 ;
        RECT 1410.890 1966.260 1411.210 1966.320 ;
        RECT 1412.730 1966.260 1413.050 1966.320 ;
        RECT 1409.050 1966.120 1409.370 1966.180 ;
        RECT 1411.810 1966.120 1412.130 1966.180 ;
        RECT 1409.050 1965.980 1412.130 1966.120 ;
        RECT 1409.050 1965.920 1409.370 1965.980 ;
        RECT 1411.810 1965.920 1412.130 1965.980 ;
        RECT 1408.130 1965.780 1408.450 1965.840 ;
        RECT 1417.790 1965.780 1418.110 1965.840 ;
        RECT 1408.130 1965.640 1418.110 1965.780 ;
        RECT 1408.130 1965.580 1408.450 1965.640 ;
        RECT 1417.790 1965.580 1418.110 1965.640 ;
        RECT 1408.130 1962.040 1408.450 1962.100 ;
        RECT 1418.250 1962.040 1418.570 1962.100 ;
        RECT 1408.130 1961.900 1418.570 1962.040 ;
        RECT 1408.130 1961.840 1408.450 1961.900 ;
        RECT 1418.250 1961.840 1418.570 1961.900 ;
        RECT 1552.110 1949.120 1552.430 1949.180 ;
        RECT 1690.110 1949.120 1690.430 1949.180 ;
        RECT 1552.110 1948.980 1690.430 1949.120 ;
        RECT 1552.110 1948.920 1552.430 1948.980 ;
        RECT 1690.110 1948.920 1690.430 1948.980 ;
        RECT 1408.130 1940.960 1408.450 1941.020 ;
        RECT 1416.870 1940.960 1417.190 1941.020 ;
        RECT 1408.130 1940.820 1417.190 1940.960 ;
        RECT 1408.130 1940.760 1408.450 1940.820 ;
        RECT 1416.870 1940.760 1417.190 1940.820 ;
        RECT 1408.130 1935.180 1408.450 1935.240 ;
        RECT 1417.330 1935.180 1417.650 1935.240 ;
        RECT 1408.130 1935.040 1417.650 1935.180 ;
        RECT 1408.130 1934.980 1408.450 1935.040 ;
        RECT 1417.330 1934.980 1417.650 1935.040 ;
        RECT 1408.590 1930.420 1408.910 1930.480 ;
        RECT 1421.010 1930.420 1421.330 1930.480 ;
        RECT 1408.590 1930.280 1421.330 1930.420 ;
        RECT 1408.590 1930.220 1408.910 1930.280 ;
        RECT 1421.010 1930.220 1421.330 1930.280 ;
        RECT 1408.130 1928.040 1408.450 1928.100 ;
        RECT 1420.550 1928.040 1420.870 1928.100 ;
        RECT 1408.130 1927.900 1420.870 1928.040 ;
        RECT 1408.130 1927.840 1408.450 1927.900 ;
        RECT 1420.550 1927.840 1420.870 1927.900 ;
        RECT 1408.130 1924.640 1408.450 1924.700 ;
        RECT 1420.090 1924.640 1420.410 1924.700 ;
        RECT 1408.130 1924.500 1420.410 1924.640 ;
        RECT 1408.130 1924.440 1408.450 1924.500 ;
        RECT 1420.090 1924.440 1420.410 1924.500 ;
        RECT 1408.590 1919.200 1408.910 1919.260 ;
        RECT 1408.590 1919.060 1412.500 1919.200 ;
        RECT 1408.590 1919.000 1408.910 1919.060 ;
        RECT 1412.360 1918.920 1412.500 1919.060 ;
        RECT 1409.050 1918.860 1409.370 1918.920 ;
        RECT 1411.810 1918.860 1412.130 1918.920 ;
        RECT 1409.050 1918.720 1412.130 1918.860 ;
        RECT 1409.050 1918.660 1409.370 1918.720 ;
        RECT 1411.810 1918.660 1412.130 1918.720 ;
        RECT 1412.270 1918.660 1412.590 1918.920 ;
        RECT 1410.890 1918.520 1411.210 1918.580 ;
        RECT 1412.730 1918.520 1413.050 1918.580 ;
        RECT 1410.890 1918.380 1413.050 1918.520 ;
        RECT 1410.890 1918.320 1411.210 1918.380 ;
        RECT 1412.730 1918.320 1413.050 1918.380 ;
        RECT 1414.110 1918.180 1414.430 1918.240 ;
        RECT 1493.690 1918.180 1494.010 1918.240 ;
        RECT 1414.110 1918.040 1494.010 1918.180 ;
        RECT 1414.110 1917.980 1414.430 1918.040 ;
        RECT 1493.690 1917.980 1494.010 1918.040 ;
        RECT 1408.590 1911.040 1408.910 1911.100 ;
        RECT 1697.470 1911.040 1697.790 1911.100 ;
        RECT 1408.590 1910.900 1697.790 1911.040 ;
        RECT 1408.590 1910.840 1408.910 1910.900 ;
        RECT 1697.470 1910.840 1697.790 1910.900 ;
        RECT 1408.130 1910.020 1408.450 1910.080 ;
        RECT 1419.630 1910.020 1419.950 1910.080 ;
        RECT 1408.130 1909.880 1419.950 1910.020 ;
        RECT 1408.130 1909.820 1408.450 1909.880 ;
        RECT 1419.630 1909.820 1419.950 1909.880 ;
        RECT 1414.110 1904.240 1414.430 1904.300 ;
        RECT 1690.570 1904.240 1690.890 1904.300 ;
        RECT 1414.110 1904.100 1690.890 1904.240 ;
        RECT 1414.110 1904.040 1414.430 1904.100 ;
        RECT 1690.570 1904.040 1690.890 1904.100 ;
        RECT 1414.110 1897.440 1414.430 1897.500 ;
        RECT 1684.130 1897.440 1684.450 1897.500 ;
        RECT 1414.110 1897.300 1684.450 1897.440 ;
        RECT 1414.110 1897.240 1414.430 1897.300 ;
        RECT 1684.130 1897.240 1684.450 1897.300 ;
        RECT 1414.110 1890.640 1414.430 1890.700 ;
        RECT 1683.670 1890.640 1683.990 1890.700 ;
        RECT 1414.110 1890.500 1683.990 1890.640 ;
        RECT 1414.110 1890.440 1414.430 1890.500 ;
        RECT 1683.670 1890.440 1683.990 1890.500 ;
        RECT 1410.890 1890.300 1411.210 1890.360 ;
        RECT 1676.770 1890.300 1677.090 1890.360 ;
        RECT 1410.890 1890.160 1677.090 1890.300 ;
        RECT 1410.890 1890.100 1411.210 1890.160 ;
        RECT 1676.770 1890.100 1677.090 1890.160 ;
        RECT 1414.110 1883.500 1414.430 1883.560 ;
        RECT 1669.870 1883.500 1670.190 1883.560 ;
        RECT 1414.110 1883.360 1670.190 1883.500 ;
        RECT 1414.110 1883.300 1414.430 1883.360 ;
        RECT 1669.870 1883.300 1670.190 1883.360 ;
        RECT 1414.110 1876.700 1414.430 1876.760 ;
        RECT 1662.970 1876.700 1663.290 1876.760 ;
        RECT 1414.110 1876.560 1663.290 1876.700 ;
        RECT 1414.110 1876.500 1414.430 1876.560 ;
        RECT 1662.970 1876.500 1663.290 1876.560 ;
        RECT 1409.510 1869.900 1409.830 1869.960 ;
        RECT 1412.730 1869.900 1413.050 1869.960 ;
        RECT 1409.510 1869.760 1413.050 1869.900 ;
        RECT 1409.510 1869.700 1409.830 1869.760 ;
        RECT 1412.730 1869.700 1413.050 1869.760 ;
        RECT 1414.110 1869.900 1414.430 1869.960 ;
        RECT 1656.070 1869.900 1656.390 1869.960 ;
        RECT 1414.110 1869.760 1656.390 1869.900 ;
        RECT 1414.110 1869.700 1414.430 1869.760 ;
        RECT 1656.070 1869.700 1656.390 1869.760 ;
        RECT 1410.890 1869.560 1411.210 1869.620 ;
        RECT 1649.630 1869.560 1649.950 1869.620 ;
        RECT 1410.890 1869.420 1649.950 1869.560 ;
        RECT 1410.890 1869.360 1411.210 1869.420 ;
        RECT 1649.630 1869.360 1649.950 1869.420 ;
        RECT 1409.050 1869.220 1409.370 1869.280 ;
        RECT 1411.810 1869.220 1412.130 1869.280 ;
        RECT 1409.050 1869.080 1412.130 1869.220 ;
        RECT 1409.050 1869.020 1409.370 1869.080 ;
        RECT 1411.810 1869.020 1412.130 1869.080 ;
        RECT 1412.270 1869.020 1412.590 1869.280 ;
        RECT 1408.590 1868.880 1408.910 1868.940 ;
        RECT 1412.360 1868.880 1412.500 1869.020 ;
        RECT 1408.590 1868.740 1412.500 1868.880 ;
        RECT 1408.590 1868.680 1408.910 1868.740 ;
        RECT 1414.110 1862.760 1414.430 1862.820 ;
        RECT 1649.170 1862.760 1649.490 1862.820 ;
        RECT 1414.110 1862.620 1649.490 1862.760 ;
        RECT 1414.110 1862.560 1414.430 1862.620 ;
        RECT 1649.170 1862.560 1649.490 1862.620 ;
        RECT 1414.110 1855.960 1414.430 1856.020 ;
        RECT 1642.270 1855.960 1642.590 1856.020 ;
        RECT 1414.110 1855.820 1642.590 1855.960 ;
        RECT 1414.110 1855.760 1414.430 1855.820 ;
        RECT 1642.270 1855.760 1642.590 1855.820 ;
        RECT 1410.890 1855.620 1411.210 1855.680 ;
        RECT 1635.370 1855.620 1635.690 1855.680 ;
        RECT 1410.890 1855.480 1635.690 1855.620 ;
        RECT 1410.890 1855.420 1411.210 1855.480 ;
        RECT 1635.370 1855.420 1635.690 1855.480 ;
        RECT 1414.110 1849.160 1414.430 1849.220 ;
        RECT 1628.470 1849.160 1628.790 1849.220 ;
        RECT 1414.110 1849.020 1628.790 1849.160 ;
        RECT 1414.110 1848.960 1414.430 1849.020 ;
        RECT 1628.470 1848.960 1628.790 1849.020 ;
        RECT 1414.110 1842.360 1414.430 1842.420 ;
        RECT 1621.570 1842.360 1621.890 1842.420 ;
        RECT 1414.110 1842.220 1621.890 1842.360 ;
        RECT 1414.110 1842.160 1414.430 1842.220 ;
        RECT 1621.570 1842.160 1621.890 1842.220 ;
        RECT 1414.110 1835.220 1414.430 1835.280 ;
        RECT 1614.670 1835.220 1614.990 1835.280 ;
        RECT 1414.110 1835.080 1614.990 1835.220 ;
        RECT 1414.110 1835.020 1414.430 1835.080 ;
        RECT 1614.670 1835.020 1614.990 1835.080 ;
        RECT 1410.890 1834.880 1411.210 1834.940 ;
        RECT 1607.770 1834.880 1608.090 1834.940 ;
        RECT 1410.890 1834.740 1608.090 1834.880 ;
        RECT 1410.890 1834.680 1411.210 1834.740 ;
        RECT 1607.770 1834.680 1608.090 1834.740 ;
        RECT 1414.110 1828.420 1414.430 1828.480 ;
        RECT 1652.390 1828.420 1652.710 1828.480 ;
        RECT 1414.110 1828.280 1652.710 1828.420 ;
        RECT 1414.110 1828.220 1414.430 1828.280 ;
        RECT 1652.390 1828.220 1652.710 1828.280 ;
        RECT 1408.590 1822.640 1408.910 1822.700 ;
        RECT 1408.590 1822.500 1412.500 1822.640 ;
        RECT 1408.590 1822.440 1408.910 1822.500 ;
        RECT 1412.360 1822.360 1412.500 1822.500 ;
        RECT 1409.050 1822.300 1409.370 1822.360 ;
        RECT 1411.810 1822.300 1412.130 1822.360 ;
        RECT 1409.050 1822.160 1412.130 1822.300 ;
        RECT 1409.050 1822.100 1409.370 1822.160 ;
        RECT 1411.810 1822.100 1412.130 1822.160 ;
        RECT 1412.270 1822.100 1412.590 1822.360 ;
        RECT 1409.510 1821.960 1409.830 1822.020 ;
        RECT 1412.730 1821.960 1413.050 1822.020 ;
        RECT 1409.510 1821.820 1413.050 1821.960 ;
        RECT 1409.510 1821.760 1409.830 1821.820 ;
        RECT 1412.730 1821.760 1413.050 1821.820 ;
        RECT 1414.110 1821.620 1414.430 1821.680 ;
        RECT 1646.410 1821.620 1646.730 1821.680 ;
        RECT 1414.110 1821.480 1646.730 1821.620 ;
        RECT 1414.110 1821.420 1414.430 1821.480 ;
        RECT 1646.410 1821.420 1646.730 1821.480 ;
        RECT 1410.890 1814.820 1411.210 1814.880 ;
        RECT 1413.650 1814.820 1413.970 1814.880 ;
        RECT 1410.890 1814.680 1413.970 1814.820 ;
        RECT 1410.890 1814.620 1411.210 1814.680 ;
        RECT 1413.650 1814.620 1413.970 1814.680 ;
        RECT 1414.110 1814.480 1414.430 1814.540 ;
        RECT 1645.490 1814.480 1645.810 1814.540 ;
        RECT 1414.110 1814.340 1645.810 1814.480 ;
        RECT 1414.110 1814.280 1414.430 1814.340 ;
        RECT 1645.490 1814.280 1645.810 1814.340 ;
        RECT 1413.650 1814.140 1413.970 1814.200 ;
        RECT 1638.590 1814.140 1638.910 1814.200 ;
        RECT 1413.650 1814.000 1638.910 1814.140 ;
        RECT 1413.650 1813.940 1413.970 1814.000 ;
        RECT 1638.590 1813.940 1638.910 1814.000 ;
        RECT 1408.590 1807.680 1408.910 1807.740 ;
        RECT 1631.690 1807.680 1632.010 1807.740 ;
        RECT 1408.590 1807.540 1632.010 1807.680 ;
        RECT 1408.590 1807.480 1408.910 1807.540 ;
        RECT 1631.690 1807.480 1632.010 1807.540 ;
        RECT 1414.110 1800.880 1414.430 1800.940 ;
        RECT 1624.790 1800.880 1625.110 1800.940 ;
        RECT 1414.110 1800.740 1625.110 1800.880 ;
        RECT 1414.110 1800.680 1414.430 1800.740 ;
        RECT 1624.790 1800.680 1625.110 1800.740 ;
        RECT 1413.650 1800.540 1413.970 1800.600 ;
        RECT 1617.890 1800.540 1618.210 1800.600 ;
        RECT 1413.650 1800.400 1618.210 1800.540 ;
        RECT 1413.650 1800.340 1413.970 1800.400 ;
        RECT 1617.890 1800.340 1618.210 1800.400 ;
        RECT 1409.510 1793.740 1409.830 1793.800 ;
        RECT 1610.990 1793.740 1611.310 1793.800 ;
        RECT 1409.510 1793.600 1611.310 1793.740 ;
        RECT 1409.510 1793.540 1409.830 1793.600 ;
        RECT 1610.990 1793.540 1611.310 1793.600 ;
        RECT 1410.430 1773.000 1410.750 1773.060 ;
        RECT 1412.270 1773.000 1412.590 1773.060 ;
        RECT 1410.430 1772.860 1412.590 1773.000 ;
        RECT 1410.430 1772.800 1410.750 1772.860 ;
        RECT 1412.270 1772.800 1412.590 1772.860 ;
        RECT 1414.110 1745.460 1414.430 1745.520 ;
        RECT 1486.790 1745.460 1487.110 1745.520 ;
        RECT 1414.110 1745.320 1487.110 1745.460 ;
        RECT 1414.110 1745.260 1414.430 1745.320 ;
        RECT 1486.790 1745.260 1487.110 1745.320 ;
        RECT 1414.110 1738.660 1414.430 1738.720 ;
        RECT 1472.990 1738.660 1473.310 1738.720 ;
        RECT 1414.110 1738.520 1473.310 1738.660 ;
        RECT 1414.110 1738.460 1414.430 1738.520 ;
        RECT 1472.990 1738.460 1473.310 1738.520 ;
        RECT 1411.350 1738.320 1411.670 1738.380 ;
        RECT 1459.190 1738.320 1459.510 1738.380 ;
        RECT 1411.350 1738.180 1459.510 1738.320 ;
        RECT 1411.350 1738.120 1411.670 1738.180 ;
        RECT 1459.190 1738.120 1459.510 1738.180 ;
        RECT 1410.430 1731.860 1410.750 1731.920 ;
        RECT 1452.290 1731.860 1452.610 1731.920 ;
        RECT 1410.430 1731.720 1452.610 1731.860 ;
        RECT 1410.430 1731.660 1410.750 1731.720 ;
        RECT 1452.290 1731.660 1452.610 1731.720 ;
        RECT 1414.110 1722.680 1414.430 1722.740 ;
        RECT 1438.490 1722.680 1438.810 1722.740 ;
        RECT 1414.110 1722.540 1438.810 1722.680 ;
        RECT 1414.110 1722.480 1414.430 1722.540 ;
        RECT 1438.490 1722.480 1438.810 1722.540 ;
        RECT 1412.730 1717.920 1413.050 1717.980 ;
        RECT 1507.490 1717.920 1507.810 1717.980 ;
        RECT 1412.730 1717.780 1507.810 1717.920 ;
        RECT 1412.730 1717.720 1413.050 1717.780 ;
        RECT 1507.490 1717.720 1507.810 1717.780 ;
        RECT 1413.650 1717.580 1413.970 1717.640 ;
        RECT 1431.590 1717.580 1431.910 1717.640 ;
        RECT 1413.650 1717.440 1431.910 1717.580 ;
        RECT 1413.650 1717.380 1413.970 1717.440 ;
        RECT 1431.590 1717.380 1431.910 1717.440 ;
        RECT 1414.110 1711.120 1414.430 1711.180 ;
        RECT 1580.170 1711.120 1580.490 1711.180 ;
        RECT 1414.110 1710.980 1580.490 1711.120 ;
        RECT 1414.110 1710.920 1414.430 1710.980 ;
        RECT 1580.170 1710.920 1580.490 1710.980 ;
        RECT 1410.890 1669.640 1411.210 1669.700 ;
        RECT 1535.090 1669.640 1535.410 1669.700 ;
        RECT 1410.890 1669.500 1535.410 1669.640 ;
        RECT 1410.890 1669.440 1411.210 1669.500 ;
        RECT 1535.090 1669.440 1535.410 1669.500 ;
        RECT 1408.130 1667.940 1408.450 1668.000 ;
        RECT 1419.170 1667.940 1419.490 1668.000 ;
        RECT 1408.130 1667.800 1419.490 1667.940 ;
        RECT 1408.130 1667.740 1408.450 1667.800 ;
        RECT 1419.170 1667.740 1419.490 1667.800 ;
        RECT 1409.970 1659.100 1410.290 1659.160 ;
        RECT 1413.650 1659.100 1413.970 1659.160 ;
        RECT 1409.970 1658.960 1413.970 1659.100 ;
        RECT 1409.970 1658.900 1410.290 1658.960 ;
        RECT 1413.650 1658.900 1413.970 1658.960 ;
        RECT 1408.130 1656.040 1408.450 1656.100 ;
        RECT 1601.330 1656.040 1601.650 1656.100 ;
        RECT 1408.130 1655.900 1601.650 1656.040 ;
        RECT 1408.130 1655.840 1408.450 1655.900 ;
        RECT 1601.330 1655.840 1601.650 1655.900 ;
        RECT 1408.130 1648.900 1408.450 1648.960 ;
        RECT 1593.970 1648.900 1594.290 1648.960 ;
        RECT 1408.130 1648.760 1594.290 1648.900 ;
        RECT 1408.130 1648.700 1408.450 1648.760 ;
        RECT 1593.970 1648.700 1594.290 1648.760 ;
        RECT 1407.670 1648.560 1407.990 1648.620 ;
        RECT 1487.250 1648.560 1487.570 1648.620 ;
        RECT 1407.670 1648.420 1487.570 1648.560 ;
        RECT 1407.670 1648.360 1407.990 1648.420 ;
        RECT 1487.250 1648.360 1487.570 1648.420 ;
        RECT 1407.670 1642.100 1407.990 1642.160 ;
        RECT 1514.390 1642.100 1514.710 1642.160 ;
        RECT 1407.670 1641.960 1514.710 1642.100 ;
        RECT 1407.670 1641.900 1407.990 1641.960 ;
        RECT 1514.390 1641.900 1514.710 1641.960 ;
        RECT 1407.670 1635.300 1407.990 1635.360 ;
        RECT 1591.210 1635.300 1591.530 1635.360 ;
        RECT 1407.670 1635.160 1591.530 1635.300 ;
        RECT 1407.670 1635.100 1407.990 1635.160 ;
        RECT 1591.210 1635.100 1591.530 1635.160 ;
        RECT 1410.430 1632.240 1410.750 1632.300 ;
        RECT 1413.650 1632.240 1413.970 1632.300 ;
        RECT 1410.430 1632.100 1413.970 1632.240 ;
        RECT 1410.430 1632.040 1410.750 1632.100 ;
        RECT 1413.650 1632.040 1413.970 1632.100 ;
        RECT 1409.510 1631.900 1409.830 1631.960 ;
        RECT 1410.890 1631.900 1411.210 1631.960 ;
        RECT 1409.510 1631.760 1411.210 1631.900 ;
        RECT 1409.510 1631.700 1409.830 1631.760 ;
        RECT 1410.890 1631.700 1411.210 1631.760 ;
        RECT 1411.350 1631.900 1411.670 1631.960 ;
        RECT 1413.190 1631.900 1413.510 1631.960 ;
        RECT 1411.350 1631.760 1413.510 1631.900 ;
        RECT 1411.350 1631.700 1411.670 1631.760 ;
        RECT 1413.190 1631.700 1413.510 1631.760 ;
        RECT 1409.050 1631.560 1409.370 1631.620 ;
        RECT 1413.650 1631.560 1413.970 1631.620 ;
        RECT 1409.050 1631.420 1413.970 1631.560 ;
        RECT 1409.050 1631.360 1409.370 1631.420 ;
        RECT 1413.650 1631.360 1413.970 1631.420 ;
        RECT 1407.670 1628.160 1407.990 1628.220 ;
        RECT 1590.750 1628.160 1591.070 1628.220 ;
        RECT 1407.670 1628.020 1591.070 1628.160 ;
        RECT 1407.670 1627.960 1407.990 1628.020 ;
        RECT 1590.750 1627.960 1591.070 1628.020 ;
        RECT 1407.670 1621.360 1407.990 1621.420 ;
        RECT 1590.290 1621.360 1590.610 1621.420 ;
        RECT 1407.670 1621.220 1590.610 1621.360 ;
        RECT 1407.670 1621.160 1407.990 1621.220 ;
        RECT 1590.290 1621.160 1590.610 1621.220 ;
        RECT 1407.670 1614.560 1407.990 1614.620 ;
        RECT 1528.190 1614.560 1528.510 1614.620 ;
        RECT 1407.670 1614.420 1528.510 1614.560 ;
        RECT 1407.670 1614.360 1407.990 1614.420 ;
        RECT 1528.190 1614.360 1528.510 1614.420 ;
        RECT 1421.470 1611.160 1421.790 1611.220 ;
        RECT 1427.910 1611.160 1428.230 1611.220 ;
        RECT 1688.730 1611.160 1689.050 1611.220 ;
        RECT 1421.470 1611.020 1689.050 1611.160 ;
        RECT 1421.470 1610.960 1421.790 1611.020 ;
        RECT 1427.910 1610.960 1428.230 1611.020 ;
        RECT 1688.730 1610.960 1689.050 1611.020 ;
        RECT 1414.110 1607.760 1414.430 1607.820 ;
        RECT 1421.470 1607.760 1421.790 1607.820 ;
        RECT 1414.110 1607.620 1421.790 1607.760 ;
        RECT 1414.110 1607.560 1414.430 1607.620 ;
        RECT 1421.470 1607.560 1421.790 1607.620 ;
        RECT 1414.110 1605.040 1414.430 1605.100 ;
        RECT 1686.890 1605.040 1687.210 1605.100 ;
        RECT 1690.110 1605.040 1690.430 1605.100 ;
        RECT 1414.110 1604.900 1690.430 1605.040 ;
      LAYER met1 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met1 ;
        RECT 1414.110 1604.840 1414.430 1604.900 ;
        RECT 1686.890 1604.840 1687.210 1604.900 ;
        RECT 1690.110 1604.840 1690.430 1604.900 ;
        RECT 1410.890 1604.700 1411.210 1604.760 ;
        RECT 2097.670 1604.700 2097.990 1604.760 ;
        RECT 1410.890 1604.560 2097.990 1604.700 ;
        RECT 1410.890 1604.500 1411.210 1604.560 ;
        RECT 2097.670 1604.500 2097.990 1604.560 ;
        RECT 1412.730 1604.360 1413.050 1604.420 ;
        RECT 2099.050 1604.360 2099.370 1604.420 ;
        RECT 1412.730 1604.220 2099.370 1604.360 ;
        RECT 1412.730 1604.160 1413.050 1604.220 ;
        RECT 2099.050 1604.160 2099.370 1604.220 ;
        RECT 1411.810 1603.000 1412.130 1603.060 ;
        RECT 2098.590 1603.000 2098.910 1603.060 ;
        RECT 1411.810 1602.860 2098.910 1603.000 ;
        RECT 1411.810 1602.800 1412.130 1602.860 ;
        RECT 2098.590 1602.800 2098.910 1602.860 ;
        RECT 1409.970 1602.660 1410.290 1602.720 ;
        RECT 2098.130 1602.660 2098.450 1602.720 ;
        RECT 1409.970 1602.520 2098.450 1602.660 ;
        RECT 1409.970 1602.460 1410.290 1602.520 ;
        RECT 2098.130 1602.460 2098.450 1602.520 ;
        RECT 1412.270 1602.320 1412.590 1602.380 ;
        RECT 2082.030 1602.320 2082.350 1602.380 ;
        RECT 1412.270 1602.180 2082.350 1602.320 ;
        RECT 1412.270 1602.120 1412.590 1602.180 ;
        RECT 2082.030 1602.120 2082.350 1602.180 ;
        RECT 1411.350 1601.980 1411.670 1602.040 ;
        RECT 2100.890 1601.980 2101.210 1602.040 ;
        RECT 1411.350 1601.840 2101.210 1601.980 ;
        RECT 1411.350 1601.780 1411.670 1601.840 ;
        RECT 2100.890 1601.780 2101.210 1601.840 ;
        RECT 1413.650 1601.640 1413.970 1601.700 ;
        RECT 2099.510 1601.640 2099.830 1601.700 ;
        RECT 1413.650 1601.500 2099.830 1601.640 ;
        RECT 1413.650 1601.440 1413.970 1601.500 ;
        RECT 2099.510 1601.440 2099.830 1601.500 ;
        RECT 1410.430 1601.300 1410.750 1601.360 ;
        RECT 2099.970 1601.300 2100.290 1601.360 ;
        RECT 1410.430 1601.160 2100.290 1601.300 ;
        RECT 1410.430 1601.100 1410.750 1601.160 ;
        RECT 2099.970 1601.100 2100.290 1601.160 ;
        RECT 1690.110 1593.820 1690.430 1593.880 ;
        RECT 1720.010 1593.820 1720.330 1593.880 ;
        RECT 1690.110 1593.680 1720.330 1593.820 ;
        RECT 1690.110 1593.620 1690.430 1593.680 ;
        RECT 1720.010 1593.620 1720.330 1593.680 ;
        RECT 1720.010 1590.420 1720.330 1590.480 ;
        RECT 1738.870 1590.420 1739.190 1590.480 ;
        RECT 1720.010 1590.280 1739.190 1590.420 ;
        RECT 1720.010 1590.220 1720.330 1590.280 ;
        RECT 1738.870 1590.220 1739.190 1590.280 ;
      LAYER via ;
        RECT 1317.540 3266.760 1317.800 3267.020 ;
        RECT 1890.700 3266.760 1890.960 3267.020 ;
        RECT 646.400 3263.700 646.660 3263.960 ;
        RECT 668.480 3263.700 668.740 3263.960 ;
        RECT 697.000 3264.040 697.260 3264.300 ;
        RECT 1890.700 3264.040 1890.960 3264.300 ;
        RECT 1917.380 3264.040 1917.640 3264.300 ;
        RECT 1939.000 3264.040 1939.260 3264.300 ;
        RECT 1293.160 3263.700 1293.420 3263.960 ;
        RECT 1317.540 3263.700 1317.800 3263.960 ;
        RECT 986.800 3254.520 987.060 3254.780 ;
        RECT 1034.640 3254.520 1034.900 3254.780 ;
        RECT 976.220 3253.840 976.480 3254.100 ;
        RECT 986.800 3253.840 987.060 3254.100 ;
        RECT 1035.100 3252.820 1035.360 3253.080 ;
        RECT 688.260 3252.140 688.520 3252.400 ;
        RECT 737.940 3252.140 738.200 3252.400 ;
        RECT 738.400 3251.800 738.660 3252.060 ;
        RECT 786.240 3251.800 786.500 3252.060 ;
        RECT 786.700 3251.800 786.960 3252.060 ;
        RECT 820.740 3251.460 821.000 3251.720 ;
        RECT 821.200 3251.460 821.460 3251.720 ;
        RECT 976.220 3251.800 976.480 3252.060 ;
        RECT 1186.900 3252.480 1187.160 3252.740 ;
        RECT 1187.820 3251.800 1188.080 3252.060 ;
        RECT 1331.800 3252.140 1332.060 3252.400 ;
        RECT 1427.940 3251.460 1428.200 3251.720 ;
        RECT 1932.100 3251.460 1932.360 3251.720 ;
        RECT 1400.340 3250.440 1400.600 3250.700 ;
        RECT 1427.940 3250.780 1428.200 3251.040 ;
        RECT 1331.800 3250.100 1332.060 3250.360 ;
        RECT 1352.500 3250.100 1352.760 3250.360 ;
        RECT 1486.820 3229.360 1487.080 3229.620 ;
        RECT 1535.580 3229.360 1535.840 3229.620 ;
        RECT 1473.020 3222.220 1473.280 3222.480 ;
        RECT 1535.580 3222.220 1535.840 3222.480 ;
        RECT 1459.220 3215.420 1459.480 3215.680 ;
        RECT 1535.580 3215.420 1535.840 3215.680 ;
        RECT 1452.320 3208.620 1452.580 3208.880 ;
        RECT 1538.340 3208.620 1538.600 3208.880 ;
        RECT 1438.520 3201.480 1438.780 3201.740 ;
        RECT 1538.340 3201.480 1538.600 3201.740 ;
        RECT 1431.620 3194.680 1431.880 3194.940 ;
        RECT 1533.280 3194.680 1533.540 3194.940 ;
        RECT 1507.520 3187.880 1507.780 3188.140 ;
        RECT 1534.200 3187.880 1534.460 3188.140 ;
        RECT 1352.040 2946.480 1352.300 2946.740 ;
        RECT 1548.920 2946.480 1549.180 2946.740 ;
        RECT 284.380 2804.360 284.640 2804.620 ;
        RECT 944.940 2804.360 945.200 2804.620 ;
        RECT 1528.220 2804.360 1528.480 2804.620 ;
        RECT 1548.920 2800.960 1549.180 2801.220 ;
        RECT 1552.140 2800.960 1552.400 2801.220 ;
        RECT 1945.900 2800.960 1946.160 2801.220 ;
        RECT 310.140 2794.160 310.400 2794.420 ;
        RECT 986.800 2794.160 987.060 2794.420 ;
        RECT 1076.500 2794.160 1076.760 2794.420 ;
        RECT 1122.500 2794.160 1122.760 2794.420 ;
        RECT 1677.260 2794.160 1677.520 2794.420 ;
        RECT 1724.180 2794.160 1724.440 2794.420 ;
        RECT 337.280 2793.820 337.540 2794.080 ;
        RECT 1007.500 2793.820 1007.760 2794.080 ;
        RECT 1642.300 2793.820 1642.560 2794.080 ;
        RECT 1690.140 2793.820 1690.400 2794.080 ;
        RECT 386.960 2793.480 387.220 2793.740 ;
        RECT 432.040 2793.480 432.300 2793.740 ;
        RECT 478.960 2793.480 479.220 2793.740 ;
        RECT 527.720 2793.480 527.980 2793.740 ;
        RECT 627.540 2793.480 627.800 2793.740 ;
        RECT 1042.000 2793.480 1042.260 2793.740 ;
        RECT 1048.440 2793.480 1048.700 2793.740 ;
        RECT 1117.900 2793.480 1118.160 2793.740 ;
        RECT 1159.300 2793.480 1159.560 2793.740 ;
        RECT 1642.760 2793.480 1643.020 2793.740 ;
        RECT 1689.680 2793.480 1689.940 2793.740 ;
        RECT 380.060 2793.140 380.320 2793.400 ;
        RECT 421.460 2793.140 421.720 2793.400 ;
        RECT 466.540 2793.140 466.800 2793.400 ;
        RECT 489.080 2793.140 489.340 2793.400 ;
        RECT 665.720 2793.140 665.980 2793.400 ;
        RECT 1122.500 2793.140 1122.760 2793.400 ;
        RECT 1166.200 2793.140 1166.460 2793.400 ;
        RECT 1724.180 2793.140 1724.440 2793.400 ;
        RECT 1766.500 2793.140 1766.760 2793.400 ;
        RECT 426.060 2792.800 426.320 2793.060 ;
        RECT 474.360 2792.800 474.620 2793.060 ;
        RECT 519.440 2792.800 519.700 2793.060 ;
        RECT 520.820 2792.800 521.080 2793.060 ;
        RECT 524.040 2792.800 524.300 2793.060 ;
        RECT 686.880 2792.800 687.140 2793.060 ;
        RECT 1088.920 2792.800 1089.180 2793.060 ;
        RECT 1129.400 2792.800 1129.660 2793.060 ;
        RECT 1174.480 2792.800 1174.740 2793.060 ;
        RECT 1682.320 2792.800 1682.580 2793.060 ;
        RECT 1728.780 2792.800 1729.040 2793.060 ;
        RECT 1773.400 2792.800 1773.660 2793.060 ;
        RECT 398.000 2792.460 398.260 2792.720 ;
        RECT 444.460 2792.460 444.720 2792.720 ;
        RECT 490.460 2792.460 490.720 2792.720 ;
        RECT 497.820 2792.460 498.080 2792.720 ;
        RECT 541.520 2792.460 541.780 2792.720 ;
        RECT 1048.440 2792.460 1048.700 2792.720 ;
        RECT 1089.840 2792.460 1090.100 2792.720 ;
        RECT 392.480 2792.120 392.740 2792.380 ;
        RECT 439.400 2792.120 439.660 2792.380 ;
        RECT 484.940 2792.120 485.200 2792.380 ;
        RECT 534.620 2792.120 534.880 2792.380 ;
        RECT 542.440 2792.120 542.700 2792.380 ;
        RECT 720.920 2792.120 721.180 2792.380 ;
        RECT 1069.600 2792.120 1069.860 2792.380 ;
        RECT 1117.900 2792.460 1118.160 2792.720 ;
        RECT 1652.420 2792.460 1652.680 2792.720 ;
        RECT 1699.340 2792.460 1699.600 2792.720 ;
        RECT 1747.640 2792.460 1747.900 2792.720 ;
        RECT 1788.580 2792.460 1788.840 2792.720 ;
        RECT 403.980 2791.780 404.240 2792.040 ;
        RECT 449.060 2791.780 449.320 2792.040 ;
        RECT 497.820 2791.780 498.080 2792.040 ;
        RECT 363.040 2791.440 363.300 2791.700 ;
        RECT 409.500 2791.440 409.760 2791.700 ;
        RECT 455.500 2791.440 455.760 2791.700 ;
        RECT 462.400 2791.440 462.660 2791.700 ;
        RECT 490.000 2791.440 490.260 2791.700 ;
        RECT 490.460 2791.440 490.720 2791.700 ;
        RECT 502.880 2791.780 503.140 2792.040 ;
        RECT 509.780 2791.780 510.040 2792.040 ;
        RECT 700.220 2791.780 700.480 2792.040 ;
        RECT 1042.920 2791.780 1043.180 2792.040 ;
        RECT 1053.040 2791.780 1053.300 2792.040 ;
        RECT 501.960 2791.440 502.220 2791.700 ;
        RECT 700.680 2791.440 700.940 2791.700 ;
        RECT 1055.800 2791.440 1056.060 2791.700 ;
        RECT 1059.020 2791.440 1059.280 2791.700 ;
        RECT 1075.580 2791.440 1075.840 2791.700 ;
        RECT 1089.840 2791.780 1090.100 2792.040 ;
        RECT 1135.840 2792.120 1136.100 2792.380 ;
        RECT 1159.300 2792.120 1159.560 2792.380 ;
        RECT 1688.760 2792.120 1689.020 2792.380 ;
        RECT 1734.300 2792.120 1734.560 2792.380 ;
        RECT 1780.300 2792.120 1780.560 2792.380 ;
        RECT 1100.420 2791.440 1100.680 2791.700 ;
        RECT 1104.100 2791.440 1104.360 2791.700 ;
        RECT 1105.480 2791.440 1105.740 2791.700 ;
        RECT 1147.800 2791.780 1148.060 2792.040 ;
        RECT 1193.800 2791.780 1194.060 2792.040 ;
        RECT 1646.440 2791.780 1646.700 2792.040 ;
        RECT 1695.200 2791.780 1695.460 2792.040 ;
        RECT 1741.200 2791.780 1741.460 2792.040 ;
        RECT 1787.200 2791.780 1787.460 2792.040 ;
        RECT 1107.780 2791.440 1108.040 2791.700 ;
        RECT 1152.400 2791.440 1152.660 2791.700 ;
        RECT 1663.460 2791.440 1663.720 2791.700 ;
        RECT 1712.680 2791.440 1712.940 2791.700 ;
        RECT 1740.740 2791.440 1741.000 2791.700 ;
        RECT 406.280 2791.100 406.540 2791.360 ;
        RECT 727.820 2791.100 728.080 2791.360 ;
        RECT 384.200 2790.760 384.460 2791.020 ;
        RECT 707.120 2790.760 707.380 2791.020 ;
        RECT 1034.640 2790.760 1034.900 2791.020 ;
        RECT 1076.500 2790.760 1076.760 2791.020 ;
        RECT 1111.920 2791.100 1112.180 2791.360 ;
        RECT 1159.300 2791.100 1159.560 2791.360 ;
        RECT 1656.560 2791.100 1656.820 2791.360 ;
        RECT 1658.860 2791.100 1659.120 2791.360 ;
        RECT 1706.240 2791.100 1706.500 2791.360 ;
        RECT 1752.700 2791.100 1752.960 2791.360 ;
        RECT 369.020 2790.420 369.280 2790.680 ;
        RECT 414.100 2790.420 414.360 2790.680 ;
        RECT 419.160 2790.420 419.420 2790.680 ;
        RECT 762.320 2790.420 762.580 2790.680 ;
        RECT 397.080 2790.080 397.340 2790.340 ;
        RECT 741.620 2790.080 741.880 2790.340 ;
        RECT 371.320 2789.740 371.580 2790.000 ;
        RECT 679.520 2789.740 679.780 2790.000 ;
        RECT 1017.620 2789.740 1017.880 2790.000 ;
        RECT 1065.460 2789.740 1065.720 2790.000 ;
        RECT 1094.900 2790.080 1095.160 2790.340 ;
        RECT 1140.900 2790.760 1141.160 2791.020 ;
        RECT 1186.900 2790.760 1187.160 2791.020 ;
        RECT 1670.360 2790.760 1670.620 2791.020 ;
        RECT 1718.200 2790.760 1718.460 2791.020 ;
        RECT 1759.600 2790.760 1759.860 2791.020 ;
        RECT 1418.740 2790.420 1419.000 2790.680 ;
        RECT 1773.400 2790.420 1773.660 2790.680 ;
        RECT 1631.720 2789.740 1631.980 2790.000 ;
        RECT 1677.260 2789.740 1677.520 2790.000 ;
        RECT 414.100 2789.400 414.360 2789.660 ;
        RECT 462.400 2789.400 462.660 2789.660 ;
        RECT 468.840 2789.400 469.100 2789.660 ;
        RECT 636.280 2789.400 636.540 2789.660 ;
        RECT 648.240 2789.400 648.500 2789.660 ;
        RECT 1042.920 2789.400 1043.180 2789.660 ;
        RECT 1514.420 2789.400 1514.680 2789.660 ;
        RECT 1587.100 2789.400 1587.360 2789.660 ;
        RECT 1617.920 2789.400 1618.180 2789.660 ;
        RECT 1663.460 2789.400 1663.720 2789.660 ;
        RECT 399.840 2789.060 400.100 2789.320 ;
        RECT 514.380 2789.060 514.640 2789.320 ;
        RECT 606.840 2789.060 607.100 2789.320 ;
        RECT 1030.500 2789.060 1030.760 2789.320 ;
        RECT 1034.640 2789.060 1034.900 2789.320 ;
        RECT 1045.220 2789.060 1045.480 2789.320 ;
        RECT 1094.900 2789.060 1095.160 2789.320 ;
        RECT 1487.280 2789.060 1487.540 2789.320 ;
        RECT 1600.900 2789.060 1601.160 2789.320 ;
        RECT 1611.020 2789.060 1611.280 2789.320 ;
        RECT 1656.560 2789.060 1656.820 2789.320 ;
        RECT 330.840 2788.720 331.100 2788.980 ;
        RECT 1001.060 2788.720 1001.320 2788.980 ;
        RECT 1010.720 2788.720 1010.980 2788.980 ;
        RECT 1055.800 2788.720 1056.060 2788.980 ;
        RECT 1624.820 2788.720 1625.080 2788.980 ;
        RECT 1670.360 2788.720 1670.620 2788.980 ;
        RECT 375.000 2788.380 375.260 2788.640 ;
        RECT 421.000 2788.380 421.260 2788.640 ;
        RECT 466.540 2788.380 466.800 2788.640 ;
        RECT 499.200 2788.380 499.460 2788.640 ;
        RECT 537.380 2788.380 537.640 2788.640 ;
        RECT 707.580 2788.380 707.840 2788.640 ;
        RECT 1024.520 2788.380 1024.780 2788.640 ;
        RECT 1069.600 2788.380 1069.860 2788.640 ;
        RECT 1418.280 2788.380 1418.540 2788.640 ;
        RECT 1759.600 2788.380 1759.860 2788.640 ;
        RECT 317.040 2788.040 317.300 2788.300 ;
        RECT 993.700 2788.040 993.960 2788.300 ;
        RECT 1038.320 2788.040 1038.580 2788.300 ;
        RECT 1088.920 2788.040 1089.180 2788.300 ;
        RECT 1417.820 2788.040 1418.080 2788.300 ;
        RECT 1766.500 2788.040 1766.760 2788.300 ;
        RECT 455.500 2787.700 455.760 2787.960 ;
        RECT 500.120 2787.700 500.380 2787.960 ;
        RECT 499.200 2787.360 499.460 2787.620 ;
        RECT 513.920 2787.700 514.180 2787.960 ;
        RECT 502.880 2787.360 503.140 2787.620 ;
        RECT 538.760 2787.700 539.020 2787.960 ;
        RECT 542.440 2787.700 542.700 2787.960 ;
        RECT 636.280 2787.700 636.540 2787.960 ;
        RECT 658.820 2787.700 659.080 2787.960 ;
        RECT 1638.620 2787.700 1638.880 2787.960 ;
        RECT 1682.320 2787.700 1682.580 2787.960 ;
        RECT 387.880 2728.540 388.140 2728.800 ;
        RECT 944.020 2728.540 944.280 2728.800 ;
        RECT 288.060 2725.140 288.320 2725.400 ;
        RECT 564.060 2725.140 564.320 2725.400 ;
        RECT 574.640 2725.140 574.900 2725.400 ;
        RECT 1010.720 2725.140 1010.980 2725.400 ;
        RECT 448.140 2724.800 448.400 2725.060 ;
        RECT 886.060 2724.800 886.320 2725.060 ;
        RECT 461.940 2724.460 462.200 2724.720 ;
        RECT 906.760 2724.460 907.020 2724.720 ;
        RECT 481.260 2724.120 481.520 2724.380 ;
        RECT 941.720 2724.120 941.980 2724.380 ;
        RECT 455.040 2723.780 455.300 2724.040 ;
        RECT 896.180 2723.780 896.440 2724.040 ;
        RECT 482.640 2723.440 482.900 2723.700 ;
        RECT 948.160 2723.440 948.420 2723.700 ;
        RECT 470.680 2723.100 470.940 2723.360 ;
        RECT 942.180 2723.100 942.440 2723.360 ;
        RECT 449.980 2722.760 450.240 2723.020 ;
        RECT 943.100 2722.760 943.360 2723.020 ;
        RECT 285.300 2722.420 285.560 2722.680 ;
        RECT 512.540 2722.420 512.800 2722.680 ;
        RECT 517.140 2722.420 517.400 2722.680 ;
        RECT 1010.260 2722.420 1010.520 2722.680 ;
        RECT 287.140 2722.080 287.400 2722.340 ;
        RECT 543.360 2722.080 543.620 2722.340 ;
        RECT 551.640 2722.080 551.900 2722.340 ;
        RECT 1060.860 2722.080 1061.120 2722.340 ;
        RECT 408.580 2721.740 408.840 2722.000 ;
        RECT 979.900 2721.740 980.160 2722.000 ;
        RECT 434.340 2721.400 434.600 2721.660 ;
        RECT 865.360 2721.400 865.620 2721.660 ;
        RECT 441.240 2721.060 441.500 2721.320 ;
        RECT 875.480 2721.060 875.740 2721.320 ;
        RECT 433.880 2720.720 434.140 2720.980 ;
        RECT 854.780 2720.720 855.040 2720.980 ;
        RECT 427.440 2720.380 427.700 2720.640 ;
        RECT 844.200 2720.380 844.460 2720.640 ;
        RECT 365.340 2720.040 365.600 2720.300 ;
        RECT 740.700 2720.040 740.960 2720.300 ;
        RECT 514.380 2719.700 514.640 2719.960 ;
        RECT 802.800 2719.700 803.060 2719.960 ;
        RECT 287.600 2719.360 287.860 2719.620 ;
        RECT 553.940 2719.360 554.200 2719.620 ;
        RECT 286.680 2719.020 286.940 2719.280 ;
        RECT 533.240 2719.020 533.500 2719.280 ;
        RECT 286.220 2718.680 286.480 2718.940 ;
        RECT 522.660 2718.680 522.920 2718.940 ;
        RECT 358.440 2718.340 358.700 2718.600 ;
        RECT 377.300 2718.340 377.560 2718.600 ;
        RECT 379.140 2718.340 379.400 2718.600 ;
        RECT 761.400 2718.340 761.660 2718.600 ;
        RECT 762.320 2718.340 762.580 2718.600 ;
        RECT 834.080 2718.340 834.340 2718.600 ;
        RECT 1034.640 2718.340 1034.900 2718.600 ;
        RECT 1102.260 2718.340 1102.520 2718.600 ;
        RECT 1145.040 2718.340 1145.300 2718.600 ;
        RECT 1300.980 2718.340 1301.240 2718.600 ;
        RECT 392.940 2718.000 393.200 2718.260 ;
        RECT 782.100 2718.000 782.360 2718.260 ;
        RECT 1027.740 2718.000 1028.000 2718.260 ;
        RECT 1093.520 2718.000 1093.780 2718.260 ;
        RECT 1138.140 2718.000 1138.400 2718.260 ;
        RECT 1290.400 2718.000 1290.660 2718.260 ;
        RECT 305.080 2717.660 305.340 2717.920 ;
        RECT 310.140 2717.660 310.400 2717.920 ;
        RECT 351.080 2717.660 351.340 2717.920 ;
        RECT 356.600 2717.660 356.860 2717.920 ;
        RECT 413.640 2717.660 413.900 2717.920 ;
        RECT 823.500 2717.660 823.760 2717.920 ;
        RECT 1041.540 2717.660 1041.800 2717.920 ;
        RECT 1114.220 2717.660 1114.480 2717.920 ;
        RECT 1151.940 2717.660 1152.200 2717.920 ;
        RECT 1311.100 2717.660 1311.360 2717.920 ;
        RECT 636.740 2717.320 637.000 2717.580 ;
        RECT 1045.220 2717.320 1045.480 2717.580 ;
        RECT 1048.440 2717.320 1048.700 2717.580 ;
        RECT 1122.500 2717.320 1122.760 2717.580 ;
        RECT 1158.840 2717.320 1159.100 2717.580 ;
        RECT 1321.680 2717.320 1321.940 2717.580 ;
        RECT 616.040 2716.980 616.300 2717.240 ;
        RECT 1038.320 2716.980 1038.580 2717.240 ;
        RECT 1055.340 2716.980 1055.600 2717.240 ;
        RECT 1134.920 2716.980 1135.180 2717.240 ;
        RECT 1165.740 2716.980 1166.000 2717.240 ;
        RECT 1332.260 2716.980 1332.520 2717.240 ;
        RECT 595.340 2716.640 595.600 2716.900 ;
        RECT 1024.520 2716.640 1024.780 2716.900 ;
        RECT 1062.240 2716.640 1062.500 2716.900 ;
        RECT 1155.620 2716.640 1155.880 2716.900 ;
        RECT 1165.280 2716.640 1165.540 2716.900 ;
        RECT 1342.380 2716.640 1342.640 2716.900 ;
        RECT 585.220 2716.300 585.480 2716.560 ;
        RECT 1017.620 2716.300 1017.880 2716.560 ;
        RECT 1076.040 2716.300 1076.300 2716.560 ;
        RECT 1176.320 2716.300 1176.580 2716.560 ;
        RECT 1179.540 2716.300 1179.800 2716.560 ;
        RECT 1363.080 2716.300 1363.340 2716.560 ;
        RECT 468.380 2715.960 468.640 2716.220 ;
        RECT 916.880 2715.960 917.140 2716.220 ;
        RECT 1054.880 2715.960 1055.140 2716.220 ;
        RECT 1145.500 2715.960 1145.760 2716.220 ;
        RECT 1172.640 2715.960 1172.900 2716.220 ;
        RECT 1352.960 2715.960 1353.220 2716.220 ;
        RECT 284.840 2715.620 285.100 2715.880 ;
        RECT 398.460 2715.620 398.720 2715.880 ;
        RECT 475.740 2715.620 476.000 2715.880 ;
        RECT 937.580 2715.620 937.840 2715.880 ;
        RECT 1020.840 2715.620 1021.100 2715.880 ;
        RECT 1081.100 2715.620 1081.360 2715.880 ;
        RECT 1082.940 2715.620 1083.200 2715.880 ;
        RECT 1186.900 2715.620 1187.160 2715.880 ;
        RECT 1193.340 2715.620 1193.600 2715.880 ;
        RECT 1383.780 2715.620 1384.040 2715.880 ;
        RECT 337.740 2715.280 338.000 2715.540 ;
        RECT 491.840 2715.280 492.100 2715.540 ;
        RECT 496.440 2715.280 496.700 2715.540 ;
        RECT 968.860 2715.280 969.120 2715.540 ;
        RECT 1069.140 2715.280 1069.400 2715.540 ;
        RECT 1166.200 2715.280 1166.460 2715.540 ;
        RECT 1186.440 2715.280 1186.700 2715.540 ;
        RECT 1373.660 2715.280 1373.920 2715.540 ;
        RECT 285.760 2714.940 286.020 2715.200 ;
        RECT 501.960 2714.940 502.220 2715.200 ;
        RECT 510.240 2714.940 510.500 2715.200 ;
        RECT 989.560 2714.940 989.820 2715.200 ;
        RECT 1013.940 2714.940 1014.200 2715.200 ;
        RECT 1072.820 2714.940 1073.080 2715.200 ;
        RECT 1089.380 2714.940 1089.640 2715.200 ;
        RECT 1197.020 2714.940 1197.280 2715.200 ;
        RECT 1200.240 2714.940 1200.500 2715.200 ;
        RECT 1394.360 2714.940 1394.620 2715.200 ;
        RECT 520.820 2714.600 521.080 2714.860 ;
        RECT 688.720 2714.600 688.980 2714.860 ;
        RECT 351.540 2714.260 351.800 2714.520 ;
        RECT 367.180 2714.260 367.440 2714.520 ;
        RECT 527.720 2714.260 527.980 2714.520 ;
        RECT 699.300 2714.260 699.560 2714.520 ;
        RECT 500.120 2713.920 500.380 2714.180 ;
        RECT 657.440 2713.920 657.700 2714.180 ;
        RECT 665.720 2713.920 665.980 2714.180 ;
        RECT 513.920 2713.580 514.180 2713.840 ;
        RECT 678.600 2713.580 678.860 2713.840 ;
        RECT 686.880 2713.920 687.140 2714.180 ;
        RECT 1020.840 2714.600 1021.100 2714.860 ;
        RECT 1131.240 2714.600 1131.500 2714.860 ;
        RECT 1280.280 2714.600 1280.540 2714.860 ;
        RECT 700.220 2714.260 700.480 2714.520 ;
        RECT 1000.140 2714.260 1000.400 2714.520 ;
        RECT 1130.780 2714.260 1131.040 2714.520 ;
        RECT 1269.700 2714.260 1269.960 2714.520 ;
        RECT 958.740 2713.920 959.000 2714.180 ;
        RECT 1117.440 2713.920 1117.700 2714.180 ;
        RECT 1249.000 2713.920 1249.260 2714.180 ;
        RECT 700.680 2713.580 700.940 2713.840 ;
        RECT 979.440 2713.580 979.700 2713.840 ;
        RECT 1124.340 2713.580 1124.600 2713.840 ;
        RECT 1259.580 2713.580 1259.840 2713.840 ;
        RECT 658.820 2713.240 659.080 2713.500 ;
        RECT 927.460 2713.240 927.720 2713.500 ;
        RECT 1110.540 2713.240 1110.800 2713.500 ;
        RECT 1238.880 2713.240 1239.140 2713.500 ;
        RECT 541.520 2712.900 541.780 2713.160 ;
        RECT 730.120 2712.900 730.380 2713.160 ;
        RECT 325.780 2712.560 326.040 2712.820 ;
        RECT 330.840 2712.560 331.100 2712.820 ;
        RECT 542.440 2712.560 542.700 2712.820 ;
        RECT 720.000 2712.560 720.260 2712.820 ;
        RECT 727.820 2712.560 728.080 2712.820 ;
        RECT 813.380 2712.900 813.640 2713.160 ;
        RECT 1103.640 2712.900 1103.900 2713.160 ;
        RECT 1228.300 2712.900 1228.560 2713.160 ;
        RECT 741.620 2712.560 741.880 2712.820 ;
        RECT 792.680 2712.560 792.940 2712.820 ;
        RECT 1089.840 2712.560 1090.100 2712.820 ;
        RECT 1207.600 2712.560 1207.860 2712.820 ;
        RECT 534.620 2712.220 534.880 2712.480 ;
        RECT 709.420 2712.220 709.680 2712.480 ;
        RECT 507.020 2711.880 507.280 2712.140 ;
        RECT 668.020 2711.880 668.280 2712.140 ;
        RECT 679.520 2711.880 679.780 2712.140 ;
        RECT 707.120 2711.880 707.380 2712.140 ;
        RECT 771.980 2712.220 772.240 2712.480 ;
        RECT 1096.740 2712.220 1097.000 2712.480 ;
        RECT 1217.720 2712.220 1217.980 2712.480 ;
        RECT 750.820 2711.880 751.080 2712.140 ;
        RECT 1407.700 2145.780 1407.960 2146.040 ;
        RECT 1835.500 2145.780 1835.760 2146.040 ;
        RECT 1407.700 2138.980 1407.960 2139.240 ;
        RECT 1842.400 2138.980 1842.660 2139.240 ;
        RECT 1408.160 2132.520 1408.420 2132.780 ;
        RECT 1849.300 2132.520 1849.560 2132.780 ;
        RECT 1407.700 2132.180 1407.960 2132.440 ;
        RECT 1856.200 2132.180 1856.460 2132.440 ;
        RECT 1407.700 2125.380 1407.960 2125.640 ;
        RECT 1863.100 2125.380 1863.360 2125.640 ;
        RECT 1407.700 2118.240 1407.960 2118.500 ;
        RECT 1870.000 2118.240 1870.260 2118.500 ;
        RECT 1408.160 2111.780 1408.420 2112.040 ;
        RECT 1870.460 2111.780 1870.720 2112.040 ;
        RECT 1407.700 2111.440 1407.960 2111.700 ;
        RECT 1876.900 2111.440 1877.160 2111.700 ;
        RECT 1407.700 2104.640 1407.960 2104.900 ;
        RECT 1883.800 2104.640 1884.060 2104.900 ;
        RECT 1407.700 2097.500 1407.960 2097.760 ;
        RECT 1890.700 2097.500 1890.960 2097.760 ;
        RECT 1408.160 2091.040 1408.420 2091.300 ;
        RECT 1897.600 2091.040 1897.860 2091.300 ;
        RECT 1407.700 2090.700 1407.960 2090.960 ;
        RECT 1904.500 2090.700 1904.760 2090.960 ;
        RECT 1414.140 2083.900 1414.400 2084.160 ;
        RECT 1911.400 2083.900 1911.660 2084.160 ;
        RECT 1411.380 2077.100 1411.640 2077.360 ;
        RECT 1911.860 2077.100 1912.120 2077.360 ;
        RECT 1408.620 2070.300 1408.880 2070.560 ;
        RECT 1919.220 2070.300 1919.480 2070.560 ;
        RECT 1410.460 2069.960 1410.720 2070.220 ;
        RECT 1925.200 2069.960 1925.460 2070.220 ;
        RECT 1917.840 2069.280 1918.100 2069.540 ;
        RECT 1965.680 2069.280 1965.940 2069.540 ;
        RECT 1629.420 2068.940 1629.680 2069.200 ;
        RECT 1675.880 2068.940 1676.140 2069.200 ;
        RECT 1726.020 2068.940 1726.280 2069.200 ;
        RECT 1772.480 2068.940 1772.740 2069.200 ;
        RECT 1890.240 2068.940 1890.500 2069.200 ;
        RECT 1936.700 2068.940 1936.960 2069.200 ;
        RECT 1980.400 2068.940 1980.660 2069.200 ;
        RECT 1628.960 2068.600 1629.220 2068.860 ;
        RECT 1676.340 2068.600 1676.600 2068.860 ;
        RECT 1725.560 2068.600 1725.820 2068.860 ;
        RECT 1772.940 2068.600 1773.200 2068.860 ;
        RECT 1848.840 2068.600 1849.100 2068.860 ;
        RECT 1893.920 2068.600 1894.180 2068.860 ;
        RECT 1941.760 2068.600 1942.020 2068.860 ;
        RECT 1987.300 2068.600 1987.560 2068.860 ;
        RECT 1413.220 2068.260 1413.480 2068.520 ;
        RECT 1841.480 2068.260 1841.740 2068.520 ;
        RECT 1890.240 2068.260 1890.500 2068.520 ;
        RECT 1930.260 2068.260 1930.520 2068.520 ;
        RECT 1973.500 2068.260 1973.760 2068.520 ;
        RECT 1407.700 2067.920 1407.960 2068.180 ;
        RECT 1843.780 2067.920 1844.040 2068.180 ;
        RECT 1844.240 2067.920 1844.500 2068.180 ;
        RECT 1849.300 2067.920 1849.560 2068.180 ;
        RECT 1898.060 2067.920 1898.320 2068.180 ;
        RECT 1948.200 2067.920 1948.460 2068.180 ;
        RECT 1591.240 2067.580 1591.500 2067.840 ;
        RECT 2028.700 2067.580 2028.960 2067.840 ;
        RECT 1409.080 2067.240 1409.340 2067.500 ;
        RECT 1844.240 2067.240 1844.500 2067.500 ;
        RECT 1844.700 2067.240 1844.960 2067.500 ;
        RECT 1864.940 2067.240 1865.200 2067.500 ;
        RECT 1911.400 2067.240 1911.660 2067.500 ;
        RECT 1924.740 2067.240 1925.000 2067.500 ;
        RECT 1969.820 2067.240 1970.080 2067.500 ;
        RECT 1973.500 2067.240 1973.760 2067.500 ;
        RECT 1976.720 2067.240 1976.980 2067.500 ;
        RECT 2021.800 2067.240 2022.060 2067.500 ;
        RECT 1435.760 2066.900 1436.020 2067.160 ;
        RECT 1482.680 2066.900 1482.940 2067.160 ;
        RECT 1532.360 2066.900 1532.620 2067.160 ;
        RECT 1579.280 2066.900 1579.540 2067.160 ;
        RECT 1590.780 2066.900 1591.040 2067.160 ;
        RECT 2035.600 2066.900 2035.860 2067.160 ;
        RECT 1410.920 2066.560 1411.180 2066.820 ;
        RECT 1859.880 2066.560 1860.140 2066.820 ;
        RECT 1907.720 2066.560 1907.980 2066.820 ;
        RECT 1954.640 2066.560 1954.900 2066.820 ;
        RECT 1959.240 2066.560 1959.500 2066.820 ;
        RECT 1965.680 2066.560 1965.940 2066.820 ;
        RECT 2008.000 2066.560 2008.260 2066.820 ;
        RECT 1414.140 2066.220 1414.400 2066.480 ;
        RECT 1932.100 2066.220 1932.360 2066.480 ;
        RECT 1969.820 2066.220 1970.080 2066.480 ;
        RECT 2015.820 2066.220 2016.080 2066.480 ;
        RECT 1435.300 2065.880 1435.560 2066.140 ;
        RECT 1483.140 2065.880 1483.400 2066.140 ;
        RECT 1531.900 2065.880 1532.160 2066.140 ;
        RECT 1579.740 2065.880 1580.000 2066.140 ;
        RECT 1590.320 2065.880 1590.580 2066.140 ;
        RECT 2042.500 2065.880 2042.760 2066.140 ;
        RECT 1411.840 2065.540 1412.100 2065.800 ;
        RECT 1844.700 2065.540 1844.960 2065.800 ;
        RECT 1410.000 2065.200 1410.260 2065.460 ;
        RECT 1435.760 2065.200 1436.020 2065.460 ;
        RECT 1482.680 2065.200 1482.940 2065.460 ;
        RECT 1532.360 2065.200 1532.620 2065.460 ;
        RECT 1579.280 2065.200 1579.540 2065.460 ;
        RECT 1629.420 2065.200 1629.680 2065.460 ;
        RECT 1675.880 2065.200 1676.140 2065.460 ;
        RECT 1726.020 2065.200 1726.280 2065.460 ;
        RECT 1772.480 2065.200 1772.740 2065.460 ;
        RECT 1844.240 2065.200 1844.500 2065.460 ;
        RECT 1412.300 2064.860 1412.560 2065.120 ;
        RECT 1435.300 2064.860 1435.560 2065.120 ;
        RECT 1483.140 2064.860 1483.400 2065.120 ;
        RECT 1531.900 2064.860 1532.160 2065.120 ;
        RECT 1579.740 2064.860 1580.000 2065.120 ;
        RECT 1628.960 2064.860 1629.220 2065.120 ;
        RECT 1676.340 2064.860 1676.600 2065.120 ;
        RECT 1725.560 2064.860 1725.820 2065.120 ;
        RECT 1772.940 2064.860 1773.200 2065.120 ;
        RECT 1911.400 2065.540 1911.660 2065.800 ;
        RECT 1958.780 2065.540 1959.040 2065.800 ;
        RECT 1959.240 2065.540 1959.500 2065.800 ;
        RECT 1994.200 2065.540 1994.460 2065.800 ;
        RECT 1877.360 2065.200 1877.620 2065.460 ;
        RECT 1846.540 2064.860 1846.800 2065.120 ;
        RECT 1871.840 2064.860 1872.100 2065.120 ;
        RECT 1917.380 2064.860 1917.640 2065.120 ;
        RECT 2001.100 2065.200 2001.360 2065.460 ;
        RECT 1924.740 2064.860 1925.000 2065.120 ;
        RECT 1411.380 2064.520 1411.640 2064.780 ;
        RECT 1882.880 2064.520 1883.140 2064.780 ;
        RECT 1930.260 2064.520 1930.520 2064.780 ;
        RECT 1948.200 2064.520 1948.460 2064.780 ;
        RECT 1987.300 2064.520 1987.560 2064.780 ;
        RECT 1413.680 2064.180 1413.940 2064.440 ;
        RECT 1966.600 2064.180 1966.860 2064.440 ;
        RECT 1410.460 2063.840 1410.720 2064.100 ;
        RECT 1973.500 2063.840 1973.760 2064.100 ;
        RECT 1407.700 2063.500 1407.960 2063.760 ;
        RECT 1408.160 2063.500 1408.420 2063.760 ;
        RECT 1980.400 2063.500 1980.660 2063.760 ;
        RECT 2028.700 2063.160 2028.960 2063.420 ;
        RECT 1407.700 2062.820 1407.960 2063.080 ;
        RECT 1409.080 2062.480 1409.340 2062.740 ;
        RECT 1413.680 2062.140 1413.940 2062.400 ;
        RECT 1409.080 2061.800 1409.340 2062.060 ;
        RECT 1410.460 2061.800 1410.720 2062.060 ;
        RECT 1420.580 2061.800 1420.840 2062.060 ;
        RECT 1718.660 2061.800 1718.920 2062.060 ;
        RECT 1407.700 2061.460 1407.960 2061.720 ;
        RECT 1420.120 2061.460 1420.380 2061.720 ;
        RECT 1718.200 2061.460 1718.460 2061.720 ;
        RECT 1421.040 2061.120 1421.300 2061.380 ;
        RECT 1725.100 2061.120 1725.360 2061.380 ;
        RECT 1417.360 2060.780 1417.620 2061.040 ;
        RECT 1732.000 2060.780 1732.260 2061.040 ;
        RECT 1416.900 2060.440 1417.160 2060.700 ;
        RECT 1738.900 2060.440 1739.160 2060.700 ;
        RECT 1414.600 2060.100 1414.860 2060.360 ;
        RECT 1745.800 2060.100 1746.060 2060.360 ;
        RECT 1409.540 2059.760 1409.800 2060.020 ;
        RECT 1753.160 2059.760 1753.420 2060.020 ;
        RECT 1528.220 2059.420 1528.480 2059.680 ;
        RECT 2097.700 2059.420 2097.960 2059.680 ;
        RECT 1555.820 2059.080 1556.080 2059.340 ;
        RECT 1987.300 2059.080 1987.560 2059.340 ;
        RECT 1410.460 2058.740 1410.720 2059.000 ;
        RECT 1940.380 2058.740 1940.640 2059.000 ;
        RECT 1415.060 2058.400 1415.320 2058.660 ;
        RECT 1955.100 2058.400 1955.360 2058.660 ;
        RECT 1425.180 2058.060 1425.440 2058.320 ;
        RECT 1995.580 2058.060 1995.840 2058.320 ;
        RECT 1410.460 2057.720 1410.720 2057.980 ;
        RECT 1990.060 2057.720 1990.320 2057.980 ;
        RECT 1415.520 2057.380 1415.780 2057.640 ;
        RECT 2004.780 2057.380 2005.040 2057.640 ;
        RECT 1416.440 2057.040 1416.700 2057.300 ;
        RECT 2008.460 2057.040 2008.720 2057.300 ;
        RECT 1412.300 2056.700 1412.560 2056.960 ;
        RECT 1414.140 2056.700 1414.400 2056.960 ;
        RECT 1424.720 2056.700 1424.980 2056.960 ;
        RECT 2021.800 2056.700 2022.060 2056.960 ;
        RECT 1409.540 2056.360 1409.800 2056.620 ;
        RECT 1415.980 2056.360 1416.240 2056.620 ;
        RECT 2016.280 2056.360 2016.540 2056.620 ;
        RECT 1414.140 2056.020 1414.400 2056.280 ;
        RECT 1946.360 2056.020 1946.620 2056.280 ;
        RECT 1409.540 2055.680 1409.800 2055.940 ;
        RECT 1948.660 2055.680 1948.920 2055.940 ;
        RECT 1493.720 2053.640 1493.980 2053.900 ;
        RECT 1711.300 2053.640 1711.560 2053.900 ;
        RECT 1419.660 2053.300 1419.920 2053.560 ;
        RECT 1704.400 2053.300 1704.660 2053.560 ;
        RECT 1414.600 2052.960 1414.860 2053.220 ;
        RECT 1961.540 2052.960 1961.800 2053.220 ;
        RECT 1419.200 2052.620 1419.460 2052.880 ;
        RECT 2049.860 2052.620 2050.120 2052.880 ;
        RECT 1409.540 2050.580 1409.800 2050.840 ;
        RECT 1410.460 2039.360 1410.720 2039.620 ;
        RECT 1410.920 2039.360 1411.180 2039.620 ;
        RECT 1413.220 2039.360 1413.480 2039.620 ;
        RECT 1408.160 2039.020 1408.420 2039.280 ;
        RECT 1408.160 2038.340 1408.420 2038.600 ;
        RECT 1409.540 2038.340 1409.800 2038.600 ;
        RECT 1410.000 2038.340 1410.260 2038.600 ;
        RECT 1409.540 2037.660 1409.800 2037.920 ;
        RECT 1410.000 2037.660 1410.260 2037.920 ;
        RECT 1413.680 2037.660 1413.940 2037.920 ;
        RECT 1414.140 2021.340 1414.400 2021.600 ;
        RECT 1555.820 2021.340 1556.080 2021.600 ;
        RECT 1411.380 2014.200 1411.640 2014.460 ;
        RECT 1411.380 2013.180 1411.640 2013.440 ;
        RECT 1410.920 2012.840 1411.180 2013.100 ;
        RECT 1425.180 2012.840 1425.440 2013.100 ;
        RECT 1408.160 2005.700 1408.420 2005.960 ;
        RECT 1415.520 2005.700 1415.780 2005.960 ;
        RECT 1408.160 2000.600 1408.420 2000.860 ;
        RECT 1416.440 2000.600 1416.700 2000.860 ;
        RECT 1408.160 1997.540 1408.420 1997.800 ;
        RECT 1415.980 1997.540 1416.240 1997.800 ;
        RECT 1410.920 1990.740 1411.180 1991.000 ;
        RECT 1424.720 1990.740 1424.980 1991.000 ;
        RECT 1408.160 1972.720 1408.420 1972.980 ;
        RECT 1418.740 1972.720 1419.000 1972.980 ;
        RECT 1410.920 1966.260 1411.180 1966.520 ;
        RECT 1412.760 1966.260 1413.020 1966.520 ;
        RECT 1409.080 1965.920 1409.340 1966.180 ;
        RECT 1411.840 1965.920 1412.100 1966.180 ;
        RECT 1408.160 1965.580 1408.420 1965.840 ;
        RECT 1417.820 1965.580 1418.080 1965.840 ;
        RECT 1408.160 1961.840 1408.420 1962.100 ;
        RECT 1418.280 1961.840 1418.540 1962.100 ;
        RECT 1552.140 1948.920 1552.400 1949.180 ;
        RECT 1690.140 1948.920 1690.400 1949.180 ;
        RECT 1408.160 1940.760 1408.420 1941.020 ;
        RECT 1416.900 1940.760 1417.160 1941.020 ;
        RECT 1408.160 1934.980 1408.420 1935.240 ;
        RECT 1417.360 1934.980 1417.620 1935.240 ;
        RECT 1408.620 1930.220 1408.880 1930.480 ;
        RECT 1421.040 1930.220 1421.300 1930.480 ;
        RECT 1408.160 1927.840 1408.420 1928.100 ;
        RECT 1420.580 1927.840 1420.840 1928.100 ;
        RECT 1408.160 1924.440 1408.420 1924.700 ;
        RECT 1420.120 1924.440 1420.380 1924.700 ;
        RECT 1408.620 1919.000 1408.880 1919.260 ;
        RECT 1409.080 1918.660 1409.340 1918.920 ;
        RECT 1411.840 1918.660 1412.100 1918.920 ;
        RECT 1412.300 1918.660 1412.560 1918.920 ;
        RECT 1410.920 1918.320 1411.180 1918.580 ;
        RECT 1412.760 1918.320 1413.020 1918.580 ;
        RECT 1414.140 1917.980 1414.400 1918.240 ;
        RECT 1493.720 1917.980 1493.980 1918.240 ;
        RECT 1408.620 1910.840 1408.880 1911.100 ;
        RECT 1697.500 1910.840 1697.760 1911.100 ;
        RECT 1408.160 1909.820 1408.420 1910.080 ;
        RECT 1419.660 1909.820 1419.920 1910.080 ;
        RECT 1414.140 1904.040 1414.400 1904.300 ;
        RECT 1690.600 1904.040 1690.860 1904.300 ;
        RECT 1414.140 1897.240 1414.400 1897.500 ;
        RECT 1684.160 1897.240 1684.420 1897.500 ;
        RECT 1414.140 1890.440 1414.400 1890.700 ;
        RECT 1683.700 1890.440 1683.960 1890.700 ;
        RECT 1410.920 1890.100 1411.180 1890.360 ;
        RECT 1676.800 1890.100 1677.060 1890.360 ;
        RECT 1414.140 1883.300 1414.400 1883.560 ;
        RECT 1669.900 1883.300 1670.160 1883.560 ;
        RECT 1414.140 1876.500 1414.400 1876.760 ;
        RECT 1663.000 1876.500 1663.260 1876.760 ;
        RECT 1409.540 1869.700 1409.800 1869.960 ;
        RECT 1412.760 1869.700 1413.020 1869.960 ;
        RECT 1414.140 1869.700 1414.400 1869.960 ;
        RECT 1656.100 1869.700 1656.360 1869.960 ;
        RECT 1410.920 1869.360 1411.180 1869.620 ;
        RECT 1649.660 1869.360 1649.920 1869.620 ;
        RECT 1409.080 1869.020 1409.340 1869.280 ;
        RECT 1411.840 1869.020 1412.100 1869.280 ;
        RECT 1412.300 1869.020 1412.560 1869.280 ;
        RECT 1408.620 1868.680 1408.880 1868.940 ;
        RECT 1414.140 1862.560 1414.400 1862.820 ;
        RECT 1649.200 1862.560 1649.460 1862.820 ;
        RECT 1414.140 1855.760 1414.400 1856.020 ;
        RECT 1642.300 1855.760 1642.560 1856.020 ;
        RECT 1410.920 1855.420 1411.180 1855.680 ;
        RECT 1635.400 1855.420 1635.660 1855.680 ;
        RECT 1414.140 1848.960 1414.400 1849.220 ;
        RECT 1628.500 1848.960 1628.760 1849.220 ;
        RECT 1414.140 1842.160 1414.400 1842.420 ;
        RECT 1621.600 1842.160 1621.860 1842.420 ;
        RECT 1414.140 1835.020 1414.400 1835.280 ;
        RECT 1614.700 1835.020 1614.960 1835.280 ;
        RECT 1410.920 1834.680 1411.180 1834.940 ;
        RECT 1607.800 1834.680 1608.060 1834.940 ;
        RECT 1414.140 1828.220 1414.400 1828.480 ;
        RECT 1652.420 1828.220 1652.680 1828.480 ;
        RECT 1408.620 1822.440 1408.880 1822.700 ;
        RECT 1409.080 1822.100 1409.340 1822.360 ;
        RECT 1411.840 1822.100 1412.100 1822.360 ;
        RECT 1412.300 1822.100 1412.560 1822.360 ;
        RECT 1409.540 1821.760 1409.800 1822.020 ;
        RECT 1412.760 1821.760 1413.020 1822.020 ;
        RECT 1414.140 1821.420 1414.400 1821.680 ;
        RECT 1646.440 1821.420 1646.700 1821.680 ;
        RECT 1410.920 1814.620 1411.180 1814.880 ;
        RECT 1413.680 1814.620 1413.940 1814.880 ;
        RECT 1414.140 1814.280 1414.400 1814.540 ;
        RECT 1645.520 1814.280 1645.780 1814.540 ;
        RECT 1413.680 1813.940 1413.940 1814.200 ;
        RECT 1638.620 1813.940 1638.880 1814.200 ;
        RECT 1408.620 1807.480 1408.880 1807.740 ;
        RECT 1631.720 1807.480 1631.980 1807.740 ;
        RECT 1414.140 1800.680 1414.400 1800.940 ;
        RECT 1624.820 1800.680 1625.080 1800.940 ;
        RECT 1413.680 1800.340 1413.940 1800.600 ;
        RECT 1617.920 1800.340 1618.180 1800.600 ;
        RECT 1409.540 1793.540 1409.800 1793.800 ;
        RECT 1611.020 1793.540 1611.280 1793.800 ;
        RECT 1410.460 1772.800 1410.720 1773.060 ;
        RECT 1412.300 1772.800 1412.560 1773.060 ;
        RECT 1414.140 1745.260 1414.400 1745.520 ;
        RECT 1486.820 1745.260 1487.080 1745.520 ;
        RECT 1414.140 1738.460 1414.400 1738.720 ;
        RECT 1473.020 1738.460 1473.280 1738.720 ;
        RECT 1411.380 1738.120 1411.640 1738.380 ;
        RECT 1459.220 1738.120 1459.480 1738.380 ;
        RECT 1410.460 1731.660 1410.720 1731.920 ;
        RECT 1452.320 1731.660 1452.580 1731.920 ;
        RECT 1414.140 1722.480 1414.400 1722.740 ;
        RECT 1438.520 1722.480 1438.780 1722.740 ;
        RECT 1412.760 1717.720 1413.020 1717.980 ;
        RECT 1507.520 1717.720 1507.780 1717.980 ;
        RECT 1413.680 1717.380 1413.940 1717.640 ;
        RECT 1431.620 1717.380 1431.880 1717.640 ;
        RECT 1414.140 1710.920 1414.400 1711.180 ;
        RECT 1580.200 1710.920 1580.460 1711.180 ;
        RECT 1410.920 1669.440 1411.180 1669.700 ;
        RECT 1535.120 1669.440 1535.380 1669.700 ;
        RECT 1408.160 1667.740 1408.420 1668.000 ;
        RECT 1419.200 1667.740 1419.460 1668.000 ;
        RECT 1410.000 1658.900 1410.260 1659.160 ;
        RECT 1413.680 1658.900 1413.940 1659.160 ;
        RECT 1408.160 1655.840 1408.420 1656.100 ;
        RECT 1601.360 1655.840 1601.620 1656.100 ;
        RECT 1408.160 1648.700 1408.420 1648.960 ;
        RECT 1594.000 1648.700 1594.260 1648.960 ;
        RECT 1407.700 1648.360 1407.960 1648.620 ;
        RECT 1487.280 1648.360 1487.540 1648.620 ;
        RECT 1407.700 1641.900 1407.960 1642.160 ;
        RECT 1514.420 1641.900 1514.680 1642.160 ;
        RECT 1407.700 1635.100 1407.960 1635.360 ;
        RECT 1591.240 1635.100 1591.500 1635.360 ;
        RECT 1410.460 1632.040 1410.720 1632.300 ;
        RECT 1413.680 1632.040 1413.940 1632.300 ;
        RECT 1409.540 1631.700 1409.800 1631.960 ;
        RECT 1410.920 1631.700 1411.180 1631.960 ;
        RECT 1411.380 1631.700 1411.640 1631.960 ;
        RECT 1413.220 1631.700 1413.480 1631.960 ;
        RECT 1409.080 1631.360 1409.340 1631.620 ;
        RECT 1413.680 1631.360 1413.940 1631.620 ;
        RECT 1407.700 1627.960 1407.960 1628.220 ;
        RECT 1590.780 1627.960 1591.040 1628.220 ;
        RECT 1407.700 1621.160 1407.960 1621.420 ;
        RECT 1590.320 1621.160 1590.580 1621.420 ;
        RECT 1407.700 1614.360 1407.960 1614.620 ;
        RECT 1528.220 1614.360 1528.480 1614.620 ;
        RECT 1421.500 1610.960 1421.760 1611.220 ;
        RECT 1427.940 1610.960 1428.200 1611.220 ;
        RECT 1688.760 1610.960 1689.020 1611.220 ;
        RECT 1414.140 1607.560 1414.400 1607.820 ;
        RECT 1421.500 1607.560 1421.760 1607.820 ;
        RECT 1414.140 1604.840 1414.400 1605.100 ;
        RECT 1686.920 1604.840 1687.180 1605.100 ;
        RECT 1690.140 1604.840 1690.400 1605.100 ;
        RECT 1410.920 1604.500 1411.180 1604.760 ;
        RECT 2097.700 1604.500 2097.960 1604.760 ;
        RECT 1412.760 1604.160 1413.020 1604.420 ;
        RECT 2099.080 1604.160 2099.340 1604.420 ;
        RECT 1411.840 1602.800 1412.100 1603.060 ;
        RECT 2098.620 1602.800 2098.880 1603.060 ;
        RECT 1410.000 1602.460 1410.260 1602.720 ;
        RECT 2098.160 1602.460 2098.420 1602.720 ;
        RECT 1412.300 1602.120 1412.560 1602.380 ;
        RECT 2082.060 1602.120 2082.320 1602.380 ;
        RECT 1411.380 1601.780 1411.640 1602.040 ;
        RECT 2100.920 1601.780 2101.180 1602.040 ;
        RECT 1413.680 1601.440 1413.940 1601.700 ;
        RECT 2099.540 1601.440 2099.800 1601.700 ;
        RECT 1410.460 1601.100 1410.720 1601.360 ;
        RECT 2100.000 1601.100 2100.260 1601.360 ;
        RECT 1690.140 1593.620 1690.400 1593.880 ;
        RECT 1720.040 1593.620 1720.300 1593.880 ;
        RECT 1720.040 1590.220 1720.300 1590.480 ;
        RECT 1738.900 1590.220 1739.160 1590.480 ;
      LAYER met2 ;
        RECT 1317.540 3266.730 1317.800 3267.050 ;
        RECT 1890.700 3266.730 1890.960 3267.050 ;
        RECT 646.390 3264.155 646.670 3264.525 ;
        RECT 668.470 3264.155 668.750 3264.525 ;
        RECT 646.460 3263.990 646.600 3264.155 ;
        RECT 668.540 3263.990 668.680 3264.155 ;
        RECT 697.000 3264.010 697.260 3264.330 ;
        RECT 1293.150 3264.155 1293.430 3264.525 ;
        RECT 646.400 3263.670 646.660 3263.990 ;
        RECT 668.480 3263.670 668.740 3263.990 ;
        RECT 688.260 3252.110 688.520 3252.430 ;
        RECT 288.050 3230.155 288.330 3230.525 ;
        RECT 287.590 3224.715 287.870 3225.085 ;
        RECT 287.130 3215.875 287.410 3216.245 ;
        RECT 286.670 3209.755 286.950 3210.125 ;
        RECT 286.210 3201.595 286.490 3201.965 ;
        RECT 285.290 3196.155 285.570 3196.525 ;
        RECT 284.830 2898.315 285.110 2898.685 ;
        RECT 284.370 2891.515 284.650 2891.885 ;
        RECT 284.440 2804.650 284.580 2891.515 ;
        RECT 284.380 2804.330 284.640 2804.650 ;
        RECT 284.900 2715.910 285.040 2898.315 ;
        RECT 285.360 2722.710 285.500 3196.155 ;
        RECT 285.750 3187.995 286.030 3188.365 ;
        RECT 285.300 2722.390 285.560 2722.710 ;
        RECT 284.840 2715.590 285.100 2715.910 ;
        RECT 285.820 2715.230 285.960 3187.995 ;
        RECT 286.280 2718.970 286.420 3201.595 ;
        RECT 286.740 2719.310 286.880 3209.755 ;
        RECT 287.200 2722.370 287.340 3215.875 ;
        RECT 287.140 2722.050 287.400 2722.370 ;
        RECT 287.660 2719.650 287.800 3224.715 ;
        RECT 288.120 2725.430 288.260 3230.155 ;
      LAYER met2 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met2 ;
        RECT 688.320 3248.600 688.460 3252.110 ;
        RECT 688.250 3248.230 688.530 3248.600 ;
        RECT 697.060 2948.325 697.200 3264.010 ;
        RECT 1293.220 3263.990 1293.360 3264.155 ;
        RECT 1317.600 3263.990 1317.740 3266.730 ;
        RECT 1890.760 3264.525 1890.900 3266.730 ;
        RECT 1890.690 3264.155 1890.970 3264.525 ;
        RECT 1917.370 3264.155 1917.650 3264.525 ;
        RECT 1890.700 3264.010 1890.960 3264.155 ;
        RECT 1917.380 3264.010 1917.640 3264.155 ;
        RECT 1939.000 3264.010 1939.260 3264.330 ;
        RECT 1293.160 3263.670 1293.420 3263.990 ;
        RECT 1317.540 3263.670 1317.800 3263.990 ;
        RECT 1890.760 3263.855 1890.900 3264.010 ;
        RECT 1317.600 3258.405 1317.740 3263.670 ;
        RECT 1317.530 3258.035 1317.810 3258.405 ;
        RECT 986.800 3254.490 987.060 3254.810 ;
        RECT 1034.640 3254.490 1034.900 3254.810 ;
        RECT 986.860 3254.130 987.000 3254.490 ;
        RECT 976.220 3253.810 976.480 3254.130 ;
        RECT 986.800 3253.810 987.060 3254.130 ;
        RECT 1034.700 3254.040 1034.840 3254.490 ;
        RECT 1034.700 3253.900 1035.300 3254.040 ;
        RECT 737.940 3252.170 738.200 3252.430 ;
        RECT 737.940 3252.110 738.600 3252.170 ;
        RECT 738.000 3252.090 738.600 3252.110 ;
        RECT 786.300 3252.090 786.900 3252.170 ;
        RECT 976.280 3252.090 976.420 3253.810 ;
        RECT 1035.160 3253.110 1035.300 3253.900 ;
        RECT 1035.100 3252.790 1035.360 3253.110 ;
        RECT 1186.890 3252.595 1187.170 3252.965 ;
        RECT 1187.810 3252.595 1188.090 3252.965 ;
        RECT 1186.900 3252.450 1187.160 3252.595 ;
        RECT 1187.880 3252.090 1188.020 3252.595 ;
        RECT 1331.800 3252.110 1332.060 3252.430 ;
        RECT 738.000 3252.030 738.660 3252.090 ;
        RECT 738.400 3251.770 738.660 3252.030 ;
        RECT 786.240 3252.030 786.960 3252.090 ;
        RECT 786.240 3251.770 786.500 3252.030 ;
        RECT 786.700 3251.770 786.960 3252.030 ;
        RECT 976.220 3251.770 976.480 3252.090 ;
        RECT 1187.820 3251.770 1188.080 3252.090 ;
        RECT 820.740 3251.490 821.000 3251.750 ;
        RECT 821.200 3251.490 821.460 3251.750 ;
        RECT 820.740 3251.430 821.460 3251.490 ;
        RECT 820.800 3251.350 821.400 3251.430 ;
        RECT 941.710 3230.155 941.990 3230.525 ;
        RECT 941.250 3187.995 941.530 3188.365 ;
        RECT 696.990 2947.955 697.270 2948.325 ;
        RECT 310.140 2794.130 310.400 2794.450 ;
        RECT 337.730 2794.275 338.010 2794.645 ;
        RECT 344.630 2794.275 344.910 2794.645 ;
        RECT 351.530 2794.275 351.810 2794.645 ;
        RECT 358.430 2794.275 358.710 2794.645 ;
        RECT 363.030 2794.275 363.310 2794.645 ;
        RECT 365.330 2794.275 365.610 2794.645 ;
        RECT 369.010 2794.275 369.290 2794.645 ;
        RECT 371.310 2794.275 371.590 2794.645 ;
        RECT 374.990 2794.275 375.270 2794.645 ;
        RECT 380.050 2794.275 380.330 2794.645 ;
        RECT 384.190 2794.275 384.470 2794.645 ;
        RECT 386.950 2794.275 387.230 2794.645 ;
        RECT 392.470 2794.275 392.750 2794.645 ;
        RECT 397.070 2794.275 397.350 2794.645 ;
        RECT 399.830 2794.275 400.110 2794.645 ;
        RECT 403.970 2794.275 404.250 2794.645 ;
        RECT 406.270 2794.275 406.550 2794.645 ;
        RECT 409.490 2794.275 409.770 2794.645 ;
        RECT 413.630 2794.275 413.910 2794.645 ;
        RECT 419.150 2794.275 419.430 2794.645 ;
        RECT 420.990 2794.275 421.270 2794.645 ;
        RECT 427.430 2794.275 427.710 2794.645 ;
        RECT 432.030 2794.275 432.310 2794.645 ;
        RECT 434.330 2794.275 434.610 2794.645 ;
        RECT 439.390 2794.275 439.670 2794.645 ;
        RECT 441.230 2794.275 441.510 2794.645 ;
        RECT 444.450 2794.275 444.730 2794.645 ;
        RECT 448.130 2794.275 448.410 2794.645 ;
        RECT 449.050 2794.275 449.330 2794.645 ;
        RECT 455.030 2794.275 455.310 2794.645 ;
        RECT 462.390 2794.275 462.670 2794.645 ;
        RECT 468.370 2794.275 468.650 2794.645 ;
        RECT 474.350 2794.275 474.630 2794.645 ;
        RECT 475.730 2794.275 476.010 2794.645 ;
        RECT 478.950 2794.275 479.230 2794.645 ;
        RECT 482.630 2794.275 482.910 2794.645 ;
        RECT 484.930 2794.275 485.210 2794.645 ;
        RECT 489.070 2794.275 489.350 2794.645 ;
        RECT 490.450 2794.275 490.730 2794.645 ;
        RECT 496.430 2794.275 496.710 2794.645 ;
        RECT 497.810 2794.275 498.090 2794.645 ;
        RECT 501.950 2794.275 502.230 2794.645 ;
        RECT 510.230 2794.275 510.510 2794.645 ;
        RECT 517.130 2794.275 517.410 2794.645 ;
        RECT 524.030 2794.275 524.310 2794.645 ;
        RECT 527.710 2794.275 527.990 2794.645 ;
        RECT 530.930 2794.275 531.210 2794.645 ;
        RECT 537.370 2794.275 537.650 2794.645 ;
        RECT 542.430 2794.275 542.710 2794.645 ;
        RECT 551.630 2794.275 551.910 2794.645 ;
        RECT 288.060 2725.110 288.320 2725.430 ;
        RECT 287.600 2719.330 287.860 2719.650 ;
        RECT 286.680 2718.990 286.940 2719.310 ;
        RECT 286.220 2718.650 286.480 2718.970 ;
        RECT 310.200 2717.950 310.340 2794.130 ;
        RECT 337.280 2793.790 337.540 2794.110 ;
        RECT 330.840 2788.690 331.100 2789.010 ;
        RECT 317.040 2788.010 317.300 2788.330 ;
        RECT 305.080 2717.630 305.340 2717.950 ;
        RECT 310.140 2717.630 310.400 2717.950 ;
        RECT 285.760 2714.910 286.020 2715.230 ;
        RECT 305.140 2700.000 305.280 2717.630 ;
        RECT 317.100 2700.010 317.240 2788.010 ;
        RECT 330.900 2712.850 331.040 2788.690 ;
        RECT 325.780 2712.530 326.040 2712.850 ;
        RECT 330.840 2712.530 331.100 2712.850 ;
        RECT 315.330 2700.000 317.240 2700.010 ;
        RECT 305.140 2699.940 305.430 2700.000 ;
        RECT 305.150 2696.000 305.430 2699.940 ;
        RECT 315.270 2699.870 317.240 2700.000 ;
        RECT 325.840 2700.000 325.980 2712.530 ;
        RECT 337.340 2700.010 337.480 2793.790 ;
        RECT 337.800 2715.570 337.940 2794.275 ;
        RECT 337.740 2715.250 338.000 2715.570 ;
        RECT 344.700 2712.250 344.840 2794.275 ;
        RECT 351.070 2792.915 351.350 2793.285 ;
        RECT 351.140 2717.950 351.280 2792.915 ;
        RECT 351.080 2717.630 351.340 2717.950 ;
        RECT 351.600 2714.550 351.740 2794.275 ;
        RECT 358.500 2718.630 358.640 2794.275 ;
        RECT 363.100 2791.730 363.240 2794.275 ;
        RECT 363.040 2791.410 363.300 2791.730 ;
        RECT 365.400 2720.330 365.540 2794.275 ;
        RECT 369.080 2790.710 369.220 2794.275 ;
        RECT 369.020 2790.390 369.280 2790.710 ;
        RECT 371.380 2790.030 371.520 2794.275 ;
        RECT 371.320 2789.710 371.580 2790.030 ;
        RECT 375.060 2788.670 375.200 2794.275 ;
        RECT 380.120 2793.430 380.260 2794.275 ;
        RECT 380.060 2793.110 380.320 2793.430 ;
        RECT 379.130 2790.875 379.410 2791.245 ;
        RECT 384.260 2791.050 384.400 2794.275 ;
        RECT 387.020 2793.770 387.160 2794.275 ;
        RECT 386.960 2793.450 387.220 2793.770 ;
        RECT 392.540 2792.410 392.680 2794.275 ;
        RECT 392.480 2792.090 392.740 2792.410 ;
        RECT 392.930 2791.555 393.210 2791.925 ;
        RECT 375.000 2788.350 375.260 2788.670 ;
        RECT 365.340 2720.010 365.600 2720.330 ;
        RECT 379.200 2718.630 379.340 2790.875 ;
        RECT 384.200 2790.730 384.460 2791.050 ;
        RECT 387.880 2728.510 388.140 2728.830 ;
        RECT 358.440 2718.310 358.700 2718.630 ;
        RECT 377.300 2718.310 377.560 2718.630 ;
        RECT 379.140 2718.310 379.400 2718.630 ;
        RECT 356.600 2717.630 356.860 2717.950 ;
        RECT 351.540 2714.230 351.800 2714.550 ;
        RECT 344.700 2712.110 345.300 2712.250 ;
        RECT 336.030 2700.000 337.480 2700.010 ;
        RECT 325.840 2699.940 326.130 2700.000 ;
        RECT 315.270 2696.000 315.550 2699.870 ;
        RECT 325.850 2696.000 326.130 2699.940 ;
        RECT 335.970 2699.870 337.480 2700.000 ;
        RECT 345.160 2700.010 345.300 2712.110 ;
        RECT 345.160 2700.000 346.610 2700.010 ;
        RECT 356.660 2700.000 356.800 2717.630 ;
        RECT 367.180 2714.230 367.440 2714.550 ;
        RECT 367.240 2700.000 367.380 2714.230 ;
        RECT 377.360 2700.000 377.500 2718.310 ;
        RECT 387.940 2700.000 388.080 2728.510 ;
        RECT 393.000 2718.290 393.140 2791.555 ;
        RECT 397.140 2790.370 397.280 2794.275 ;
        RECT 397.990 2792.915 398.270 2793.285 ;
        RECT 398.060 2792.750 398.200 2792.915 ;
        RECT 398.000 2792.430 398.260 2792.750 ;
        RECT 397.080 2790.050 397.340 2790.370 ;
        RECT 399.900 2789.350 400.040 2794.275 ;
        RECT 404.040 2792.070 404.180 2794.275 ;
        RECT 403.980 2791.750 404.240 2792.070 ;
        RECT 406.340 2791.390 406.480 2794.275 ;
        RECT 409.560 2791.730 409.700 2794.275 ;
        RECT 409.500 2791.410 409.760 2791.730 ;
        RECT 406.280 2791.070 406.540 2791.390 ;
        RECT 399.840 2789.030 400.100 2789.350 ;
        RECT 408.580 2721.710 408.840 2722.030 ;
        RECT 392.940 2717.970 393.200 2718.290 ;
        RECT 398.460 2715.590 398.720 2715.910 ;
        RECT 398.520 2700.000 398.660 2715.590 ;
        RECT 408.640 2700.000 408.780 2721.710 ;
        RECT 413.700 2717.950 413.840 2794.275 ;
        RECT 414.090 2792.915 414.370 2793.285 ;
        RECT 414.160 2790.710 414.300 2792.915 ;
        RECT 419.220 2790.710 419.360 2794.275 ;
        RECT 421.060 2793.170 421.200 2794.275 ;
        RECT 421.460 2793.170 421.720 2793.430 ;
        RECT 421.060 2793.110 421.720 2793.170 ;
        RECT 421.060 2793.030 421.660 2793.110 ;
        RECT 414.100 2790.390 414.360 2790.710 ;
        RECT 419.160 2790.390 419.420 2790.710 ;
        RECT 414.160 2789.690 414.300 2790.390 ;
        RECT 414.100 2789.370 414.360 2789.690 ;
        RECT 421.060 2788.670 421.200 2793.030 ;
        RECT 426.050 2792.915 426.330 2793.285 ;
        RECT 426.060 2792.770 426.320 2792.915 ;
        RECT 421.000 2788.350 421.260 2788.670 ;
        RECT 419.150 2721.515 419.430 2721.885 ;
        RECT 413.640 2717.630 413.900 2717.950 ;
        RECT 419.220 2700.000 419.360 2721.515 ;
        RECT 427.500 2720.670 427.640 2794.275 ;
        RECT 432.100 2793.770 432.240 2794.275 ;
        RECT 432.040 2793.450 432.300 2793.770 ;
        RECT 433.870 2792.915 434.150 2793.285 ;
        RECT 429.270 2722.195 429.550 2722.565 ;
        RECT 427.440 2720.350 427.700 2720.670 ;
        RECT 429.340 2700.000 429.480 2722.195 ;
        RECT 433.940 2721.010 434.080 2792.915 ;
        RECT 434.400 2721.690 434.540 2794.275 ;
        RECT 439.460 2792.410 439.600 2794.275 ;
        RECT 439.400 2792.090 439.660 2792.410 ;
        RECT 439.850 2722.875 440.130 2723.245 ;
        RECT 434.340 2721.370 434.600 2721.690 ;
        RECT 433.880 2720.690 434.140 2721.010 ;
        RECT 439.920 2700.000 440.060 2722.875 ;
        RECT 441.300 2721.350 441.440 2794.275 ;
        RECT 444.520 2792.750 444.660 2794.275 ;
        RECT 444.460 2792.430 444.720 2792.750 ;
        RECT 448.200 2725.090 448.340 2794.275 ;
        RECT 449.120 2792.070 449.260 2794.275 ;
        RECT 449.060 2791.750 449.320 2792.070 ;
        RECT 448.140 2724.770 448.400 2725.090 ;
        RECT 455.100 2724.070 455.240 2794.275 ;
        RECT 455.490 2792.915 455.770 2793.285 ;
        RECT 455.560 2791.730 455.700 2792.915 ;
        RECT 455.500 2791.410 455.760 2791.730 ;
        RECT 461.930 2791.555 462.210 2791.925 ;
        RECT 462.460 2791.730 462.600 2794.275 ;
        RECT 466.540 2793.285 466.800 2793.430 ;
        RECT 466.530 2792.915 466.810 2793.285 ;
        RECT 455.560 2787.990 455.700 2791.410 ;
        RECT 455.500 2787.670 455.760 2787.990 ;
        RECT 462.000 2724.750 462.140 2791.555 ;
        RECT 462.400 2791.410 462.660 2791.730 ;
        RECT 462.460 2789.690 462.600 2791.410 ;
        RECT 462.400 2789.370 462.660 2789.690 ;
        RECT 466.600 2788.670 466.740 2792.915 ;
        RECT 466.540 2788.350 466.800 2788.670 ;
        RECT 461.940 2724.430 462.200 2724.750 ;
        RECT 455.040 2723.750 455.300 2724.070 ;
        RECT 460.550 2723.555 460.830 2723.925 ;
        RECT 449.980 2722.730 450.240 2723.050 ;
        RECT 441.240 2721.030 441.500 2721.350 ;
        RECT 450.040 2700.000 450.180 2722.730 ;
        RECT 460.620 2700.000 460.760 2723.555 ;
        RECT 468.440 2716.250 468.580 2794.275 ;
        RECT 468.830 2792.915 469.110 2793.285 ;
        RECT 474.420 2793.090 474.560 2794.275 ;
        RECT 468.900 2789.690 469.040 2792.915 ;
        RECT 474.360 2792.770 474.620 2793.090 ;
        RECT 468.840 2789.370 469.100 2789.690 ;
        RECT 470.680 2723.070 470.940 2723.390 ;
        RECT 468.380 2715.930 468.640 2716.250 ;
        RECT 470.740 2700.000 470.880 2723.070 ;
        RECT 475.800 2715.910 475.940 2794.275 ;
        RECT 479.020 2793.770 479.160 2794.275 ;
        RECT 478.960 2793.450 479.220 2793.770 ;
        RECT 481.260 2724.090 481.520 2724.410 ;
        RECT 475.740 2715.590 476.000 2715.910 ;
        RECT 481.320 2700.000 481.460 2724.090 ;
        RECT 482.700 2723.730 482.840 2794.275 ;
        RECT 485.000 2792.410 485.140 2794.275 ;
        RECT 489.140 2793.430 489.280 2794.275 ;
        RECT 489.080 2793.110 489.340 2793.430 ;
        RECT 490.520 2792.750 490.660 2794.275 ;
        RECT 490.460 2792.430 490.720 2792.750 ;
        RECT 484.940 2792.090 485.200 2792.410 ;
        RECT 489.990 2791.555 490.270 2791.925 ;
        RECT 490.520 2791.730 490.660 2792.430 ;
        RECT 490.000 2791.410 490.260 2791.555 ;
        RECT 490.460 2791.410 490.720 2791.730 ;
        RECT 482.640 2723.410 482.900 2723.730 ;
        RECT 496.500 2715.570 496.640 2794.275 ;
        RECT 497.880 2792.750 498.020 2794.275 ;
        RECT 500.110 2792.915 500.390 2793.285 ;
        RECT 497.820 2792.430 498.080 2792.750 ;
        RECT 497.880 2792.070 498.020 2792.430 ;
        RECT 497.820 2791.750 498.080 2792.070 ;
        RECT 499.200 2788.350 499.460 2788.670 ;
        RECT 499.260 2787.650 499.400 2788.350 ;
        RECT 500.180 2787.990 500.320 2792.915 ;
        RECT 502.020 2791.730 502.160 2794.275 ;
        RECT 509.770 2792.915 510.050 2793.285 ;
        RECT 509.840 2792.070 509.980 2792.915 ;
        RECT 502.880 2791.750 503.140 2792.070 ;
        RECT 501.960 2791.410 502.220 2791.730 ;
        RECT 500.120 2787.670 500.380 2787.990 ;
        RECT 499.200 2787.330 499.460 2787.650 ;
        RECT 491.840 2715.250 492.100 2715.570 ;
        RECT 496.440 2715.250 496.700 2715.570 ;
        RECT 491.900 2700.000 492.040 2715.250 ;
        RECT 500.180 2714.210 500.320 2787.670 ;
        RECT 502.940 2787.650 503.080 2791.750 ;
        RECT 507.010 2791.555 507.290 2791.925 ;
        RECT 509.780 2791.750 510.040 2792.070 ;
        RECT 502.880 2787.330 503.140 2787.650 ;
        RECT 501.960 2714.910 502.220 2715.230 ;
        RECT 500.120 2713.890 500.380 2714.210 ;
        RECT 502.020 2700.000 502.160 2714.910 ;
        RECT 507.080 2712.170 507.220 2791.555 ;
        RECT 510.300 2715.230 510.440 2794.275 ;
        RECT 513.910 2792.915 514.190 2793.285 ;
        RECT 513.980 2787.990 514.120 2792.915 ;
        RECT 514.380 2789.030 514.640 2789.350 ;
        RECT 513.920 2787.670 514.180 2787.990 ;
        RECT 512.540 2722.390 512.800 2722.710 ;
        RECT 510.240 2714.910 510.500 2715.230 ;
        RECT 507.020 2711.850 507.280 2712.170 ;
        RECT 512.600 2700.000 512.740 2722.390 ;
        RECT 513.980 2713.870 514.120 2787.670 ;
        RECT 514.440 2719.990 514.580 2789.030 ;
        RECT 517.200 2722.710 517.340 2794.275 ;
        RECT 519.430 2792.915 519.710 2793.285 ;
        RECT 524.100 2793.090 524.240 2794.275 ;
        RECT 527.780 2793.770 527.920 2794.275 ;
        RECT 527.720 2793.450 527.980 2793.770 ;
        RECT 519.440 2792.770 519.700 2792.915 ;
        RECT 520.820 2792.770 521.080 2793.090 ;
        RECT 524.040 2792.770 524.300 2793.090 ;
        RECT 517.140 2722.390 517.400 2722.710 ;
        RECT 514.380 2719.670 514.640 2719.990 ;
        RECT 520.880 2714.890 521.020 2792.770 ;
        RECT 522.660 2718.650 522.920 2718.970 ;
        RECT 520.820 2714.570 521.080 2714.890 ;
        RECT 513.920 2713.550 514.180 2713.870 ;
        RECT 522.720 2700.000 522.860 2718.650 ;
        RECT 527.780 2714.550 527.920 2793.450 ;
        RECT 531.000 2715.085 531.140 2794.275 ;
        RECT 534.610 2792.915 534.890 2793.285 ;
        RECT 534.680 2792.410 534.820 2792.915 ;
        RECT 534.620 2792.090 534.880 2792.410 ;
        RECT 533.240 2718.990 533.500 2719.310 ;
        RECT 530.930 2714.715 531.210 2715.085 ;
        RECT 527.720 2714.230 527.980 2714.550 ;
        RECT 533.300 2700.000 533.440 2718.990 ;
        RECT 534.680 2712.510 534.820 2792.090 ;
        RECT 537.440 2788.670 537.580 2794.275 ;
        RECT 538.750 2792.915 539.030 2793.285 ;
        RECT 541.510 2792.915 541.790 2793.285 ;
        RECT 537.380 2788.350 537.640 2788.670 ;
        RECT 538.820 2787.990 538.960 2792.915 ;
        RECT 541.580 2792.750 541.720 2792.915 ;
        RECT 541.520 2792.430 541.780 2792.750 ;
        RECT 538.760 2787.670 539.020 2787.990 ;
        RECT 541.580 2713.190 541.720 2792.430 ;
        RECT 542.500 2792.410 542.640 2794.275 ;
        RECT 542.440 2792.090 542.700 2792.410 ;
        RECT 542.440 2787.670 542.700 2787.990 ;
        RECT 541.520 2712.870 541.780 2713.190 ;
        RECT 542.500 2712.850 542.640 2787.670 ;
        RECT 551.700 2722.370 551.840 2794.275 ;
        RECT 627.540 2793.450 627.800 2793.770 ;
        RECT 606.840 2789.030 607.100 2789.350 ;
        RECT 564.060 2725.110 564.320 2725.430 ;
        RECT 574.640 2725.110 574.900 2725.430 ;
        RECT 543.360 2722.050 543.620 2722.370 ;
        RECT 551.640 2722.050 551.900 2722.370 ;
        RECT 542.440 2712.530 542.700 2712.850 ;
        RECT 534.620 2712.190 534.880 2712.510 ;
        RECT 543.420 2700.000 543.560 2722.050 ;
        RECT 553.940 2719.330 554.200 2719.650 ;
        RECT 554.000 2700.000 554.140 2719.330 ;
        RECT 564.120 2700.000 564.260 2725.110 ;
        RECT 574.700 2700.000 574.840 2725.110 ;
        RECT 595.340 2716.610 595.600 2716.930 ;
        RECT 585.220 2716.270 585.480 2716.590 ;
        RECT 585.280 2700.000 585.420 2716.270 ;
        RECT 595.400 2700.000 595.540 2716.610 ;
        RECT 606.900 2700.010 607.040 2789.030 ;
        RECT 616.040 2716.950 616.300 2717.270 ;
        RECT 606.050 2700.000 607.040 2700.010 ;
        RECT 345.160 2699.870 346.830 2700.000 ;
        RECT 356.660 2699.940 356.950 2700.000 ;
        RECT 367.240 2699.940 367.530 2700.000 ;
        RECT 377.360 2699.940 377.650 2700.000 ;
        RECT 387.940 2699.940 388.230 2700.000 ;
        RECT 398.520 2699.940 398.810 2700.000 ;
        RECT 408.640 2699.940 408.930 2700.000 ;
        RECT 419.220 2699.940 419.510 2700.000 ;
        RECT 429.340 2699.940 429.630 2700.000 ;
        RECT 439.920 2699.940 440.210 2700.000 ;
        RECT 450.040 2699.940 450.330 2700.000 ;
        RECT 460.620 2699.940 460.910 2700.000 ;
        RECT 470.740 2699.940 471.030 2700.000 ;
        RECT 481.320 2699.940 481.610 2700.000 ;
        RECT 491.900 2699.940 492.190 2700.000 ;
        RECT 502.020 2699.940 502.310 2700.000 ;
        RECT 512.600 2699.940 512.890 2700.000 ;
        RECT 522.720 2699.940 523.010 2700.000 ;
        RECT 533.300 2699.940 533.590 2700.000 ;
        RECT 543.420 2699.940 543.710 2700.000 ;
        RECT 554.000 2699.940 554.290 2700.000 ;
        RECT 564.120 2699.940 564.410 2700.000 ;
        RECT 574.700 2699.940 574.990 2700.000 ;
        RECT 585.280 2699.940 585.570 2700.000 ;
        RECT 595.400 2699.940 595.690 2700.000 ;
        RECT 335.970 2696.000 336.250 2699.870 ;
        RECT 346.550 2696.000 346.830 2699.870 ;
        RECT 356.670 2696.000 356.950 2699.940 ;
        RECT 367.250 2696.000 367.530 2699.940 ;
        RECT 377.370 2696.000 377.650 2699.940 ;
        RECT 387.950 2696.000 388.230 2699.940 ;
        RECT 398.530 2696.000 398.810 2699.940 ;
        RECT 408.650 2696.000 408.930 2699.940 ;
        RECT 419.230 2696.000 419.510 2699.940 ;
        RECT 429.350 2696.000 429.630 2699.940 ;
        RECT 439.930 2696.000 440.210 2699.940 ;
        RECT 450.050 2696.000 450.330 2699.940 ;
        RECT 460.630 2696.000 460.910 2699.940 ;
        RECT 470.750 2696.000 471.030 2699.940 ;
        RECT 481.330 2696.000 481.610 2699.940 ;
        RECT 491.910 2696.000 492.190 2699.940 ;
        RECT 502.030 2696.000 502.310 2699.940 ;
        RECT 512.610 2696.000 512.890 2699.940 ;
        RECT 522.730 2696.000 523.010 2699.940 ;
        RECT 533.310 2696.000 533.590 2699.940 ;
        RECT 543.430 2696.000 543.710 2699.940 ;
        RECT 554.010 2696.000 554.290 2699.940 ;
        RECT 564.130 2696.000 564.410 2699.940 ;
        RECT 574.710 2696.000 574.990 2699.940 ;
        RECT 585.290 2696.000 585.570 2699.940 ;
        RECT 595.410 2696.000 595.690 2699.940 ;
        RECT 605.990 2699.870 607.040 2700.000 ;
        RECT 616.100 2700.000 616.240 2716.950 ;
        RECT 627.600 2700.010 627.740 2793.450 ;
        RECT 665.720 2793.110 665.980 2793.430 ;
        RECT 636.280 2789.370 636.540 2789.690 ;
        RECT 648.240 2789.370 648.500 2789.690 ;
        RECT 636.340 2787.990 636.480 2789.370 ;
        RECT 636.280 2787.670 636.540 2787.990 ;
        RECT 636.740 2717.290 637.000 2717.610 ;
        RECT 626.750 2700.000 627.740 2700.010 ;
        RECT 616.100 2699.940 616.390 2700.000 ;
        RECT 605.990 2696.000 606.270 2699.870 ;
        RECT 616.110 2696.000 616.390 2699.940 ;
        RECT 626.690 2699.870 627.740 2700.000 ;
        RECT 636.800 2700.000 636.940 2717.290 ;
        RECT 648.300 2700.010 648.440 2789.370 ;
        RECT 658.820 2787.670 659.080 2787.990 ;
        RECT 657.440 2713.890 657.700 2714.210 ;
        RECT 647.450 2700.000 648.440 2700.010 ;
        RECT 636.800 2699.940 637.090 2700.000 ;
        RECT 626.690 2696.000 626.970 2699.870 ;
        RECT 636.810 2696.000 637.090 2699.940 ;
        RECT 647.390 2699.870 648.440 2700.000 ;
        RECT 657.500 2700.000 657.640 2713.890 ;
        RECT 658.880 2713.530 659.020 2787.670 ;
        RECT 665.780 2714.210 665.920 2793.110 ;
        RECT 686.880 2792.770 687.140 2793.090 ;
        RECT 679.520 2789.710 679.780 2790.030 ;
        RECT 665.720 2713.890 665.980 2714.210 ;
        RECT 678.600 2713.550 678.860 2713.870 ;
        RECT 658.820 2713.210 659.080 2713.530 ;
        RECT 668.020 2711.850 668.280 2712.170 ;
        RECT 668.080 2700.000 668.220 2711.850 ;
        RECT 678.660 2700.000 678.800 2713.550 ;
        RECT 679.580 2712.170 679.720 2789.710 ;
        RECT 686.940 2714.210 687.080 2792.770 ;
        RECT 720.920 2792.090 721.180 2792.410 ;
        RECT 700.220 2791.750 700.480 2792.070 ;
        RECT 688.720 2714.570 688.980 2714.890 ;
        RECT 686.880 2713.890 687.140 2714.210 ;
        RECT 679.520 2711.850 679.780 2712.170 ;
        RECT 688.780 2700.000 688.920 2714.570 ;
        RECT 700.280 2714.550 700.420 2791.750 ;
        RECT 700.680 2791.410 700.940 2791.730 ;
        RECT 699.300 2714.230 699.560 2714.550 ;
        RECT 700.220 2714.230 700.480 2714.550 ;
        RECT 699.360 2700.000 699.500 2714.230 ;
        RECT 700.740 2713.870 700.880 2791.410 ;
        RECT 707.120 2790.730 707.380 2791.050 ;
        RECT 700.680 2713.550 700.940 2713.870 ;
        RECT 707.180 2712.170 707.320 2790.730 ;
        RECT 707.580 2788.350 707.840 2788.670 ;
        RECT 707.640 2716.445 707.780 2788.350 ;
        RECT 707.570 2716.075 707.850 2716.445 ;
        RECT 720.980 2715.765 721.120 2792.090 ;
        RECT 727.820 2791.070 728.080 2791.390 ;
        RECT 720.910 2715.395 721.190 2715.765 ;
        RECT 727.880 2712.850 728.020 2791.070 ;
        RECT 762.320 2790.390 762.580 2790.710 ;
        RECT 741.620 2790.050 741.880 2790.370 ;
        RECT 740.700 2720.010 740.960 2720.330 ;
        RECT 730.120 2712.870 730.380 2713.190 ;
        RECT 720.000 2712.530 720.260 2712.850 ;
        RECT 727.820 2712.530 728.080 2712.850 ;
        RECT 709.420 2712.190 709.680 2712.510 ;
        RECT 707.120 2711.850 707.380 2712.170 ;
        RECT 709.480 2700.000 709.620 2712.190 ;
        RECT 720.060 2700.000 720.200 2712.530 ;
        RECT 730.180 2700.000 730.320 2712.870 ;
        RECT 740.760 2700.000 740.900 2720.010 ;
        RECT 741.680 2712.850 741.820 2790.050 ;
        RECT 762.380 2718.630 762.520 2790.390 ;
        RECT 886.060 2724.770 886.320 2725.090 ;
        RECT 865.360 2721.370 865.620 2721.690 ;
        RECT 854.780 2720.690 855.040 2721.010 ;
        RECT 844.200 2720.350 844.460 2720.670 ;
        RECT 802.800 2719.670 803.060 2719.990 ;
        RECT 761.400 2718.310 761.660 2718.630 ;
        RECT 762.320 2718.310 762.580 2718.630 ;
        RECT 741.620 2712.530 741.880 2712.850 ;
        RECT 750.820 2711.850 751.080 2712.170 ;
        RECT 750.880 2700.000 751.020 2711.850 ;
        RECT 761.460 2700.000 761.600 2718.310 ;
        RECT 782.100 2717.970 782.360 2718.290 ;
        RECT 771.980 2712.190 772.240 2712.510 ;
        RECT 772.040 2700.000 772.180 2712.190 ;
        RECT 782.160 2700.000 782.300 2717.970 ;
        RECT 792.680 2712.530 792.940 2712.850 ;
        RECT 792.740 2700.000 792.880 2712.530 ;
        RECT 802.860 2700.000 803.000 2719.670 ;
        RECT 834.080 2718.310 834.340 2718.630 ;
        RECT 823.500 2717.630 823.760 2717.950 ;
        RECT 813.380 2712.870 813.640 2713.190 ;
        RECT 813.440 2700.000 813.580 2712.870 ;
        RECT 823.560 2700.000 823.700 2717.630 ;
        RECT 834.140 2700.000 834.280 2718.310 ;
        RECT 844.260 2700.000 844.400 2720.350 ;
        RECT 854.840 2700.000 854.980 2720.690 ;
        RECT 865.420 2700.000 865.560 2721.370 ;
        RECT 875.480 2721.030 875.740 2721.350 ;
        RECT 875.540 2700.000 875.680 2721.030 ;
        RECT 886.120 2700.000 886.260 2724.770 ;
        RECT 906.760 2724.430 907.020 2724.750 ;
        RECT 896.180 2723.750 896.440 2724.070 ;
        RECT 896.240 2700.000 896.380 2723.750 ;
        RECT 906.820 2700.000 906.960 2724.430 ;
        RECT 941.320 2721.885 941.460 3187.995 ;
        RECT 941.780 2724.410 941.920 3230.155 ;
        RECT 942.170 3224.715 942.450 3225.085 ;
        RECT 941.720 2724.090 941.980 2724.410 ;
        RECT 942.240 2723.390 942.380 3224.715 ;
        RECT 942.630 3215.875 942.910 3216.245 ;
        RECT 942.700 2723.925 942.840 3215.875 ;
        RECT 943.090 3209.755 943.370 3210.125 ;
        RECT 942.630 2723.555 942.910 2723.925 ;
        RECT 942.180 2723.070 942.440 2723.390 ;
        RECT 943.160 2723.050 943.300 3209.755 ;
        RECT 943.550 3201.595 943.830 3201.965 ;
        RECT 943.620 2723.245 943.760 3201.595 ;
        RECT 944.470 3196.155 944.750 3196.525 ;
        RECT 944.010 2898.315 944.290 2898.685 ;
        RECT 944.080 2728.830 944.220 2898.315 ;
        RECT 944.020 2728.510 944.280 2728.830 ;
        RECT 943.100 2722.730 943.360 2723.050 ;
        RECT 943.550 2722.875 943.830 2723.245 ;
        RECT 944.540 2722.565 944.680 3196.155 ;
        RECT 944.930 2891.515 945.210 2891.885 ;
        RECT 945.000 2804.650 945.140 2891.515 ;
      LAYER met2 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met2 ;
        RECT 1331.860 3250.390 1332.000 3252.110 ;
        RECT 1427.940 3251.430 1428.200 3251.750 ;
        RECT 1932.100 3251.430 1932.360 3251.750 ;
        RECT 1428.000 3251.070 1428.140 3251.430 ;
        RECT 1427.940 3250.750 1428.200 3251.070 ;
        RECT 1400.340 3250.410 1400.600 3250.730 ;
        RECT 1331.800 3250.070 1332.060 3250.390 ;
        RECT 1352.500 3250.245 1352.760 3250.390 ;
        RECT 1400.400 3250.245 1400.540 3250.410 ;
        RECT 1331.860 3249.450 1332.000 3250.070 ;
        RECT 1352.490 3249.875 1352.770 3250.245 ;
        RECT 1400.330 3249.875 1400.610 3250.245 ;
        RECT 1332.250 3249.450 1332.530 3249.565 ;
        RECT 1331.860 3249.310 1332.530 3249.450 ;
        RECT 1332.250 3249.195 1332.530 3249.310 ;
        RECT 1345.590 2946.595 1345.870 2946.965 ;
        RECT 1352.030 2946.595 1352.310 2946.965 ;
        RECT 1345.660 2938.805 1345.800 2946.595 ;
        RECT 1352.040 2946.450 1352.300 2946.595 ;
        RECT 1345.590 2938.435 1345.870 2938.805 ;
        RECT 944.940 2804.330 945.200 2804.650 ;
        RECT 1054.870 2799.715 1055.150 2800.085 ;
        RECT 979.890 2794.275 980.170 2794.645 ;
        RECT 986.790 2794.275 987.070 2794.645 ;
        RECT 1007.490 2794.275 1007.770 2794.645 ;
        RECT 1013.930 2794.275 1014.210 2794.645 ;
        RECT 1020.830 2794.275 1021.110 2794.645 ;
        RECT 1027.730 2794.275 1028.010 2794.645 ;
        RECT 1030.490 2794.275 1030.770 2794.645 ;
        RECT 1041.990 2794.275 1042.270 2794.645 ;
        RECT 1053.030 2794.275 1053.310 2794.645 ;
        RECT 948.160 2723.410 948.420 2723.730 ;
        RECT 944.470 2722.195 944.750 2722.565 ;
        RECT 941.250 2721.515 941.530 2721.885 ;
        RECT 916.880 2715.930 917.140 2716.250 ;
        RECT 916.940 2700.000 917.080 2715.930 ;
        RECT 937.580 2715.590 937.840 2715.910 ;
        RECT 927.460 2713.210 927.720 2713.530 ;
        RECT 927.520 2700.000 927.660 2713.210 ;
        RECT 937.640 2700.000 937.780 2715.590 ;
        RECT 948.220 2700.000 948.360 2723.410 ;
        RECT 979.960 2722.030 980.100 2794.275 ;
        RECT 986.800 2794.130 987.060 2794.275 ;
        RECT 1007.560 2794.110 1007.700 2794.275 ;
        RECT 1007.500 2793.790 1007.760 2794.110 ;
        RECT 1010.710 2792.915 1010.990 2793.285 ;
        RECT 1001.050 2788.835 1001.330 2789.205 ;
        RECT 1010.780 2789.010 1010.920 2792.915 ;
        RECT 1001.060 2788.690 1001.320 2788.835 ;
        RECT 1010.720 2788.690 1010.980 2789.010 ;
        RECT 993.690 2788.155 993.970 2788.525 ;
        RECT 993.700 2788.010 993.960 2788.155 ;
        RECT 1010.780 2725.430 1010.920 2788.690 ;
        RECT 1010.720 2725.110 1010.980 2725.430 ;
        RECT 1010.260 2722.390 1010.520 2722.710 ;
        RECT 979.900 2721.710 980.160 2722.030 ;
        RECT 968.860 2715.250 969.120 2715.570 ;
        RECT 958.740 2713.890 959.000 2714.210 ;
        RECT 958.800 2700.000 958.940 2713.890 ;
        RECT 968.920 2700.000 969.060 2715.250 ;
        RECT 989.560 2714.910 989.820 2715.230 ;
        RECT 979.440 2713.550 979.700 2713.870 ;
        RECT 979.500 2700.000 979.640 2713.550 ;
        RECT 989.620 2700.000 989.760 2714.910 ;
        RECT 1000.140 2714.230 1000.400 2714.550 ;
        RECT 1000.200 2700.000 1000.340 2714.230 ;
        RECT 1010.320 2700.000 1010.460 2722.390 ;
        RECT 1014.000 2715.230 1014.140 2794.275 ;
        RECT 1017.610 2793.595 1017.890 2793.965 ;
        RECT 1017.680 2790.030 1017.820 2793.595 ;
        RECT 1017.620 2789.710 1017.880 2790.030 ;
        RECT 1017.680 2716.590 1017.820 2789.710 ;
        RECT 1017.620 2716.270 1017.880 2716.590 ;
        RECT 1020.900 2715.910 1021.040 2794.275 ;
        RECT 1024.510 2792.915 1024.790 2793.285 ;
        RECT 1024.580 2788.670 1024.720 2792.915 ;
        RECT 1024.520 2788.350 1024.780 2788.670 ;
        RECT 1024.580 2716.930 1024.720 2788.350 ;
        RECT 1027.800 2718.290 1027.940 2794.275 ;
        RECT 1030.560 2789.350 1030.700 2794.275 ;
        RECT 1042.060 2793.770 1042.200 2794.275 ;
        RECT 1042.000 2793.450 1042.260 2793.770 ;
        RECT 1048.440 2793.450 1048.700 2793.770 ;
        RECT 1045.210 2792.915 1045.490 2793.285 ;
        RECT 1042.920 2791.750 1043.180 2792.070 ;
        RECT 1034.640 2790.730 1034.900 2791.050 ;
        RECT 1034.700 2789.350 1034.840 2790.730 ;
        RECT 1042.980 2789.690 1043.120 2791.750 ;
        RECT 1042.920 2789.370 1043.180 2789.690 ;
        RECT 1045.280 2789.350 1045.420 2792.915 ;
        RECT 1048.500 2792.750 1048.640 2793.450 ;
        RECT 1048.440 2792.430 1048.700 2792.750 ;
        RECT 1053.100 2792.070 1053.240 2794.275 ;
        RECT 1053.040 2791.750 1053.300 2792.070 ;
        RECT 1030.500 2789.030 1030.760 2789.350 ;
        RECT 1034.640 2789.030 1034.900 2789.350 ;
        RECT 1045.220 2789.030 1045.480 2789.350 ;
        RECT 1038.310 2788.155 1038.590 2788.525 ;
        RECT 1038.320 2788.010 1038.580 2788.155 ;
        RECT 1034.630 2787.475 1034.910 2787.845 ;
        RECT 1034.700 2718.630 1034.840 2787.475 ;
        RECT 1034.640 2718.310 1034.900 2718.630 ;
        RECT 1027.740 2717.970 1028.000 2718.290 ;
        RECT 1038.380 2717.270 1038.520 2788.010 ;
        RECT 1041.530 2787.475 1041.810 2787.845 ;
        RECT 1041.600 2717.950 1041.740 2787.475 ;
        RECT 1041.540 2717.630 1041.800 2717.950 ;
        RECT 1045.280 2717.610 1045.420 2789.030 ;
        RECT 1048.430 2787.475 1048.710 2787.845 ;
        RECT 1048.500 2717.610 1048.640 2787.475 ;
        RECT 1045.220 2717.290 1045.480 2717.610 ;
        RECT 1048.440 2717.290 1048.700 2717.610 ;
        RECT 1038.320 2716.950 1038.580 2717.270 ;
        RECT 1024.520 2716.610 1024.780 2716.930 ;
        RECT 1041.530 2716.075 1041.810 2716.445 ;
        RECT 1054.940 2716.250 1055.080 2799.715 ;
        RECT 1100.410 2794.955 1100.690 2795.325 ;
        RECT 1059.010 2794.275 1059.290 2794.645 ;
        RECT 1065.450 2794.275 1065.730 2794.645 ;
        RECT 1069.590 2794.275 1069.870 2794.645 ;
        RECT 1076.490 2794.275 1076.770 2794.645 ;
        RECT 1089.830 2794.275 1090.110 2794.645 ;
        RECT 1094.890 2794.275 1095.170 2794.645 ;
        RECT 1059.080 2791.730 1059.220 2794.275 ;
        RECT 1055.800 2791.410 1056.060 2791.730 ;
        RECT 1059.020 2791.410 1059.280 2791.730 ;
        RECT 1055.860 2789.010 1056.000 2791.410 ;
        RECT 1065.520 2790.030 1065.660 2794.275 ;
        RECT 1069.660 2792.410 1069.800 2794.275 ;
        RECT 1076.500 2794.130 1076.760 2794.275 ;
        RECT 1069.600 2792.090 1069.860 2792.410 ;
        RECT 1065.460 2789.710 1065.720 2790.030 ;
        RECT 1055.800 2788.690 1056.060 2789.010 ;
        RECT 1069.660 2788.670 1069.800 2792.090 ;
        RECT 1075.570 2791.555 1075.850 2791.925 ;
        RECT 1075.580 2791.410 1075.840 2791.555 ;
        RECT 1076.560 2791.050 1076.700 2794.130 ;
        RECT 1088.910 2793.595 1089.190 2793.965 ;
        RECT 1088.980 2793.090 1089.120 2793.595 ;
        RECT 1088.920 2792.770 1089.180 2793.090 ;
        RECT 1076.500 2790.730 1076.760 2791.050 ;
        RECT 1055.330 2788.155 1055.610 2788.525 ;
        RECT 1069.600 2788.350 1069.860 2788.670 ;
        RECT 1088.980 2788.330 1089.120 2792.770 ;
        RECT 1089.900 2792.750 1090.040 2794.275 ;
        RECT 1089.840 2792.430 1090.100 2792.750 ;
        RECT 1089.900 2792.070 1090.040 2792.430 ;
        RECT 1089.840 2791.750 1090.100 2792.070 ;
        RECT 1094.960 2790.370 1095.100 2794.275 ;
        RECT 1100.480 2791.730 1100.620 2794.955 ;
        RECT 1111.910 2794.275 1112.190 2794.645 ;
        RECT 1117.890 2794.275 1118.170 2794.645 ;
        RECT 1122.490 2794.275 1122.770 2794.645 ;
        RECT 1129.390 2794.275 1129.670 2794.645 ;
        RECT 1135.830 2794.275 1136.110 2794.645 ;
        RECT 1140.890 2794.275 1141.170 2794.645 ;
        RECT 1147.790 2794.275 1148.070 2794.645 ;
        RECT 1100.420 2791.410 1100.680 2791.730 ;
        RECT 1104.100 2791.640 1104.360 2791.730 ;
        RECT 1105.480 2791.640 1105.740 2791.730 ;
        RECT 1104.100 2791.500 1105.740 2791.640 ;
        RECT 1107.770 2791.555 1108.050 2791.925 ;
        RECT 1104.100 2791.410 1104.360 2791.500 ;
        RECT 1105.480 2791.410 1105.740 2791.500 ;
        RECT 1107.780 2791.410 1108.040 2791.555 ;
        RECT 1111.980 2791.390 1112.120 2794.275 ;
        RECT 1117.960 2793.770 1118.100 2794.275 ;
        RECT 1122.500 2794.130 1122.760 2794.275 ;
        RECT 1117.900 2793.450 1118.160 2793.770 ;
        RECT 1117.960 2792.750 1118.100 2793.450 ;
        RECT 1122.560 2793.430 1122.700 2794.130 ;
        RECT 1122.500 2793.110 1122.760 2793.430 ;
        RECT 1129.460 2793.090 1129.600 2794.275 ;
        RECT 1129.400 2792.770 1129.660 2793.090 ;
        RECT 1117.900 2792.430 1118.160 2792.750 ;
        RECT 1135.900 2792.410 1136.040 2794.275 ;
        RECT 1135.840 2792.090 1136.100 2792.410 ;
        RECT 1111.920 2791.070 1112.180 2791.390 ;
        RECT 1140.960 2791.050 1141.100 2794.275 ;
        RECT 1147.860 2792.070 1148.000 2794.275 ;
        RECT 1159.290 2793.595 1159.570 2793.965 ;
        RECT 1166.190 2793.595 1166.470 2793.965 ;
        RECT 1159.300 2793.450 1159.560 2793.595 ;
        RECT 1166.260 2793.430 1166.400 2793.595 ;
        RECT 1166.200 2793.110 1166.460 2793.430 ;
        RECT 1174.470 2792.915 1174.750 2793.285 ;
        RECT 1186.890 2792.915 1187.170 2793.285 ;
        RECT 1174.480 2792.770 1174.740 2792.915 ;
        RECT 1159.300 2792.320 1159.560 2792.410 ;
        RECT 1159.750 2792.320 1160.030 2792.605 ;
        RECT 1159.300 2792.235 1160.030 2792.320 ;
        RECT 1159.300 2792.180 1159.960 2792.235 ;
        RECT 1159.300 2792.090 1159.560 2792.180 ;
        RECT 1147.800 2791.750 1148.060 2792.070 ;
        RECT 1152.390 2791.555 1152.670 2791.925 ;
        RECT 1159.290 2791.555 1159.570 2791.925 ;
        RECT 1152.400 2791.410 1152.660 2791.555 ;
        RECT 1159.360 2791.390 1159.500 2791.555 ;
        RECT 1159.300 2791.070 1159.560 2791.390 ;
        RECT 1186.960 2791.050 1187.100 2792.915 ;
        RECT 1193.790 2792.235 1194.070 2792.605 ;
        RECT 1193.860 2792.070 1194.000 2792.235 ;
        RECT 1193.800 2791.750 1194.060 2792.070 ;
        RECT 1140.900 2790.730 1141.160 2791.050 ;
        RECT 1186.900 2790.730 1187.160 2791.050 ;
        RECT 1418.740 2790.390 1419.000 2790.710 ;
        RECT 1094.900 2790.050 1095.160 2790.370 ;
        RECT 1094.960 2789.350 1095.100 2790.050 ;
        RECT 1094.900 2789.030 1095.160 2789.350 ;
        RECT 1055.400 2717.270 1055.540 2788.155 ;
        RECT 1088.920 2788.010 1089.180 2788.330 ;
        RECT 1089.370 2788.155 1089.650 2788.525 ;
        RECT 1130.770 2788.155 1131.050 2788.525 ;
        RECT 1165.730 2788.155 1166.010 2788.525 ;
        RECT 1418.280 2788.350 1418.540 2788.670 ;
        RECT 1062.230 2787.475 1062.510 2787.845 ;
        RECT 1069.130 2787.475 1069.410 2787.845 ;
        RECT 1076.030 2787.475 1076.310 2787.845 ;
        RECT 1082.930 2787.475 1083.210 2787.845 ;
        RECT 1060.860 2722.050 1061.120 2722.370 ;
        RECT 1055.340 2716.950 1055.600 2717.270 ;
        RECT 1020.840 2715.590 1021.100 2715.910 ;
        RECT 1013.940 2714.910 1014.200 2715.230 ;
        RECT 1020.840 2714.570 1021.100 2714.890 ;
        RECT 1030.950 2714.715 1031.230 2715.085 ;
        RECT 1020.900 2700.000 1021.040 2714.570 ;
        RECT 1031.020 2700.000 1031.160 2714.715 ;
        RECT 1041.600 2700.000 1041.740 2716.075 ;
        RECT 1054.880 2715.930 1055.140 2716.250 ;
        RECT 1052.110 2715.395 1052.390 2715.765 ;
        RECT 1052.180 2700.000 1052.320 2715.395 ;
        RECT 1060.920 2700.010 1061.060 2722.050 ;
        RECT 1062.300 2716.930 1062.440 2787.475 ;
        RECT 1062.240 2716.610 1062.500 2716.930 ;
        RECT 1069.200 2715.570 1069.340 2787.475 ;
        RECT 1076.100 2716.590 1076.240 2787.475 ;
        RECT 1076.040 2716.270 1076.300 2716.590 ;
        RECT 1083.000 2715.910 1083.140 2787.475 ;
        RECT 1081.100 2715.590 1081.360 2715.910 ;
        RECT 1082.940 2715.590 1083.200 2715.910 ;
        RECT 1069.140 2715.250 1069.400 2715.570 ;
        RECT 1072.820 2714.910 1073.080 2715.230 ;
        RECT 1060.920 2700.000 1062.370 2700.010 ;
        RECT 1072.880 2700.000 1073.020 2714.910 ;
        RECT 1081.160 2700.010 1081.300 2715.590 ;
        RECT 1089.440 2715.230 1089.580 2788.155 ;
        RECT 1089.830 2787.475 1090.110 2787.845 ;
        RECT 1096.730 2787.475 1097.010 2787.845 ;
        RECT 1103.630 2787.475 1103.910 2787.845 ;
        RECT 1110.530 2787.475 1110.810 2787.845 ;
        RECT 1117.430 2787.475 1117.710 2787.845 ;
        RECT 1124.330 2787.475 1124.610 2787.845 ;
        RECT 1089.380 2714.910 1089.640 2715.230 ;
        RECT 1089.900 2712.850 1090.040 2787.475 ;
        RECT 1093.520 2717.970 1093.780 2718.290 ;
        RECT 1089.840 2712.530 1090.100 2712.850 ;
        RECT 1081.160 2700.000 1083.070 2700.010 ;
        RECT 1093.580 2700.000 1093.720 2717.970 ;
        RECT 1096.800 2712.510 1096.940 2787.475 ;
        RECT 1102.260 2718.310 1102.520 2718.630 ;
        RECT 1096.740 2712.190 1097.000 2712.510 ;
        RECT 1102.320 2700.010 1102.460 2718.310 ;
        RECT 1103.700 2713.190 1103.840 2787.475 ;
        RECT 1110.600 2713.530 1110.740 2787.475 ;
        RECT 1114.220 2717.630 1114.480 2717.950 ;
        RECT 1110.540 2713.210 1110.800 2713.530 ;
        RECT 1103.640 2712.870 1103.900 2713.190 ;
        RECT 1102.320 2700.000 1103.770 2700.010 ;
        RECT 1114.280 2700.000 1114.420 2717.630 ;
        RECT 1117.500 2714.210 1117.640 2787.475 ;
        RECT 1122.500 2717.290 1122.760 2717.610 ;
        RECT 1117.440 2713.890 1117.700 2714.210 ;
        RECT 1122.560 2700.010 1122.700 2717.290 ;
        RECT 1124.400 2713.870 1124.540 2787.475 ;
        RECT 1130.840 2714.550 1130.980 2788.155 ;
        RECT 1131.230 2787.475 1131.510 2787.845 ;
        RECT 1138.130 2787.475 1138.410 2787.845 ;
        RECT 1145.030 2787.475 1145.310 2787.845 ;
        RECT 1151.930 2787.475 1152.210 2787.845 ;
        RECT 1158.830 2787.475 1159.110 2787.845 ;
        RECT 1165.270 2787.475 1165.550 2787.845 ;
        RECT 1131.300 2714.890 1131.440 2787.475 ;
        RECT 1138.200 2718.290 1138.340 2787.475 ;
        RECT 1145.100 2718.630 1145.240 2787.475 ;
        RECT 1145.040 2718.310 1145.300 2718.630 ;
        RECT 1138.140 2717.970 1138.400 2718.290 ;
        RECT 1152.000 2717.950 1152.140 2787.475 ;
        RECT 1151.940 2717.630 1152.200 2717.950 ;
        RECT 1158.900 2717.610 1159.040 2787.475 ;
        RECT 1158.840 2717.290 1159.100 2717.610 ;
        RECT 1134.920 2716.950 1135.180 2717.270 ;
        RECT 1131.240 2714.570 1131.500 2714.890 ;
        RECT 1130.780 2714.230 1131.040 2714.550 ;
        RECT 1124.340 2713.550 1124.600 2713.870 ;
        RECT 1122.560 2700.000 1124.470 2700.010 ;
        RECT 1134.980 2700.000 1135.120 2716.950 ;
        RECT 1165.340 2716.930 1165.480 2787.475 ;
        RECT 1165.800 2717.270 1165.940 2788.155 ;
        RECT 1417.820 2788.010 1418.080 2788.330 ;
        RECT 1172.630 2787.475 1172.910 2787.845 ;
        RECT 1179.530 2787.475 1179.810 2787.845 ;
        RECT 1186.430 2787.475 1186.710 2787.845 ;
        RECT 1193.330 2787.475 1193.610 2787.845 ;
        RECT 1200.230 2787.475 1200.510 2787.845 ;
        RECT 1165.740 2716.950 1166.000 2717.270 ;
        RECT 1155.620 2716.610 1155.880 2716.930 ;
        RECT 1165.280 2716.610 1165.540 2716.930 ;
        RECT 1145.500 2715.930 1145.760 2716.250 ;
        RECT 1145.560 2700.000 1145.700 2715.930 ;
        RECT 1155.680 2700.000 1155.820 2716.610 ;
        RECT 1172.700 2716.250 1172.840 2787.475 ;
        RECT 1179.600 2716.590 1179.740 2787.475 ;
        RECT 1176.320 2716.270 1176.580 2716.590 ;
        RECT 1179.540 2716.270 1179.800 2716.590 ;
        RECT 1172.640 2715.930 1172.900 2716.250 ;
        RECT 1166.200 2715.250 1166.460 2715.570 ;
        RECT 1166.260 2700.000 1166.400 2715.250 ;
        RECT 1176.380 2700.000 1176.520 2716.270 ;
        RECT 1186.500 2715.570 1186.640 2787.475 ;
        RECT 1193.400 2715.910 1193.540 2787.475 ;
        RECT 1186.900 2715.590 1187.160 2715.910 ;
        RECT 1193.340 2715.590 1193.600 2715.910 ;
        RECT 1186.440 2715.250 1186.700 2715.570 ;
        RECT 1186.960 2700.000 1187.100 2715.590 ;
        RECT 1200.300 2715.230 1200.440 2787.475 ;
        RECT 1300.980 2718.310 1301.240 2718.630 ;
        RECT 1290.400 2717.970 1290.660 2718.290 ;
        RECT 1197.020 2714.910 1197.280 2715.230 ;
        RECT 1200.240 2714.910 1200.500 2715.230 ;
        RECT 1197.080 2700.000 1197.220 2714.910 ;
        RECT 1280.280 2714.570 1280.540 2714.890 ;
        RECT 1269.700 2714.230 1269.960 2714.550 ;
        RECT 1249.000 2713.890 1249.260 2714.210 ;
        RECT 1238.880 2713.210 1239.140 2713.530 ;
        RECT 1228.300 2712.870 1228.560 2713.190 ;
        RECT 1207.600 2712.530 1207.860 2712.850 ;
        RECT 1207.660 2700.000 1207.800 2712.530 ;
        RECT 1217.720 2712.190 1217.980 2712.510 ;
        RECT 1217.780 2700.000 1217.920 2712.190 ;
        RECT 1228.360 2700.000 1228.500 2712.870 ;
        RECT 1238.940 2700.000 1239.080 2713.210 ;
        RECT 1249.060 2700.000 1249.200 2713.890 ;
        RECT 1259.580 2713.550 1259.840 2713.870 ;
        RECT 1259.640 2700.000 1259.780 2713.550 ;
        RECT 1269.760 2700.000 1269.900 2714.230 ;
        RECT 1280.340 2700.000 1280.480 2714.570 ;
        RECT 1290.460 2700.000 1290.600 2717.970 ;
        RECT 1301.040 2700.000 1301.180 2718.310 ;
        RECT 1311.100 2717.630 1311.360 2717.950 ;
        RECT 1311.160 2700.000 1311.300 2717.630 ;
        RECT 1321.680 2717.290 1321.940 2717.610 ;
        RECT 1321.740 2700.000 1321.880 2717.290 ;
        RECT 1332.260 2716.950 1332.520 2717.270 ;
        RECT 1332.320 2700.000 1332.460 2716.950 ;
        RECT 1342.380 2716.610 1342.640 2716.930 ;
        RECT 1342.440 2700.000 1342.580 2716.610 ;
        RECT 1363.080 2716.270 1363.340 2716.590 ;
        RECT 1352.960 2715.930 1353.220 2716.250 ;
        RECT 1353.020 2700.000 1353.160 2715.930 ;
        RECT 1363.140 2700.000 1363.280 2716.270 ;
        RECT 1383.780 2715.590 1384.040 2715.910 ;
        RECT 1373.660 2715.250 1373.920 2715.570 ;
        RECT 1373.720 2700.000 1373.860 2715.250 ;
        RECT 1383.840 2700.000 1383.980 2715.590 ;
        RECT 1394.360 2714.910 1394.620 2715.230 ;
        RECT 1394.420 2700.000 1394.560 2714.910 ;
        RECT 657.500 2699.940 657.790 2700.000 ;
        RECT 668.080 2699.940 668.370 2700.000 ;
        RECT 678.660 2699.940 678.950 2700.000 ;
        RECT 688.780 2699.940 689.070 2700.000 ;
        RECT 699.360 2699.940 699.650 2700.000 ;
        RECT 709.480 2699.940 709.770 2700.000 ;
        RECT 720.060 2699.940 720.350 2700.000 ;
        RECT 730.180 2699.940 730.470 2700.000 ;
        RECT 740.760 2699.940 741.050 2700.000 ;
        RECT 750.880 2699.940 751.170 2700.000 ;
        RECT 761.460 2699.940 761.750 2700.000 ;
        RECT 772.040 2699.940 772.330 2700.000 ;
        RECT 782.160 2699.940 782.450 2700.000 ;
        RECT 792.740 2699.940 793.030 2700.000 ;
        RECT 802.860 2699.940 803.150 2700.000 ;
        RECT 813.440 2699.940 813.730 2700.000 ;
        RECT 823.560 2699.940 823.850 2700.000 ;
        RECT 834.140 2699.940 834.430 2700.000 ;
        RECT 844.260 2699.940 844.550 2700.000 ;
        RECT 854.840 2699.940 855.130 2700.000 ;
        RECT 865.420 2699.940 865.710 2700.000 ;
        RECT 875.540 2699.940 875.830 2700.000 ;
        RECT 886.120 2699.940 886.410 2700.000 ;
        RECT 896.240 2699.940 896.530 2700.000 ;
        RECT 906.820 2699.940 907.110 2700.000 ;
        RECT 916.940 2699.940 917.230 2700.000 ;
        RECT 927.520 2699.940 927.810 2700.000 ;
        RECT 937.640 2699.940 937.930 2700.000 ;
        RECT 948.220 2699.940 948.510 2700.000 ;
        RECT 958.800 2699.940 959.090 2700.000 ;
        RECT 968.920 2699.940 969.210 2700.000 ;
        RECT 979.500 2699.940 979.790 2700.000 ;
        RECT 989.620 2699.940 989.910 2700.000 ;
        RECT 1000.200 2699.940 1000.490 2700.000 ;
        RECT 1010.320 2699.940 1010.610 2700.000 ;
        RECT 1020.900 2699.940 1021.190 2700.000 ;
        RECT 1031.020 2699.940 1031.310 2700.000 ;
        RECT 1041.600 2699.940 1041.890 2700.000 ;
        RECT 1052.180 2699.940 1052.470 2700.000 ;
        RECT 647.390 2696.000 647.670 2699.870 ;
        RECT 657.510 2696.000 657.790 2699.940 ;
        RECT 668.090 2696.000 668.370 2699.940 ;
        RECT 678.670 2696.000 678.950 2699.940 ;
        RECT 688.790 2696.000 689.070 2699.940 ;
        RECT 699.370 2696.000 699.650 2699.940 ;
        RECT 709.490 2696.000 709.770 2699.940 ;
        RECT 720.070 2696.000 720.350 2699.940 ;
        RECT 730.190 2696.000 730.470 2699.940 ;
        RECT 740.770 2696.000 741.050 2699.940 ;
        RECT 750.890 2696.000 751.170 2699.940 ;
        RECT 761.470 2696.000 761.750 2699.940 ;
        RECT 772.050 2696.000 772.330 2699.940 ;
        RECT 782.170 2696.000 782.450 2699.940 ;
        RECT 792.750 2696.000 793.030 2699.940 ;
        RECT 802.870 2696.000 803.150 2699.940 ;
        RECT 813.450 2696.000 813.730 2699.940 ;
        RECT 823.570 2696.000 823.850 2699.940 ;
        RECT 834.150 2696.000 834.430 2699.940 ;
        RECT 844.270 2696.000 844.550 2699.940 ;
        RECT 854.850 2696.000 855.130 2699.940 ;
        RECT 865.430 2696.000 865.710 2699.940 ;
        RECT 875.550 2696.000 875.830 2699.940 ;
        RECT 886.130 2696.000 886.410 2699.940 ;
        RECT 896.250 2696.000 896.530 2699.940 ;
        RECT 906.830 2696.000 907.110 2699.940 ;
        RECT 916.950 2696.000 917.230 2699.940 ;
        RECT 927.530 2696.000 927.810 2699.940 ;
        RECT 937.650 2696.000 937.930 2699.940 ;
        RECT 948.230 2696.000 948.510 2699.940 ;
        RECT 958.810 2696.000 959.090 2699.940 ;
        RECT 968.930 2696.000 969.210 2699.940 ;
        RECT 979.510 2696.000 979.790 2699.940 ;
        RECT 989.630 2696.000 989.910 2699.940 ;
        RECT 1000.210 2696.000 1000.490 2699.940 ;
        RECT 1010.330 2696.000 1010.610 2699.940 ;
        RECT 1020.910 2696.000 1021.190 2699.940 ;
        RECT 1031.030 2696.000 1031.310 2699.940 ;
        RECT 1041.610 2696.000 1041.890 2699.940 ;
        RECT 1052.190 2696.000 1052.470 2699.940 ;
        RECT 1060.920 2699.870 1062.590 2700.000 ;
        RECT 1072.880 2699.940 1073.170 2700.000 ;
        RECT 1062.310 2696.000 1062.590 2699.870 ;
        RECT 1072.890 2696.000 1073.170 2699.940 ;
        RECT 1081.160 2699.870 1083.290 2700.000 ;
        RECT 1093.580 2699.940 1093.870 2700.000 ;
        RECT 1083.010 2696.000 1083.290 2699.870 ;
        RECT 1093.590 2696.000 1093.870 2699.940 ;
        RECT 1102.320 2699.870 1103.990 2700.000 ;
        RECT 1114.280 2699.940 1114.570 2700.000 ;
        RECT 1103.710 2696.000 1103.990 2699.870 ;
        RECT 1114.290 2696.000 1114.570 2699.940 ;
        RECT 1122.560 2699.870 1124.690 2700.000 ;
        RECT 1134.980 2699.940 1135.270 2700.000 ;
        RECT 1145.560 2699.940 1145.850 2700.000 ;
        RECT 1155.680 2699.940 1155.970 2700.000 ;
        RECT 1166.260 2699.940 1166.550 2700.000 ;
        RECT 1176.380 2699.940 1176.670 2700.000 ;
        RECT 1186.960 2699.940 1187.250 2700.000 ;
        RECT 1197.080 2699.940 1197.370 2700.000 ;
        RECT 1207.660 2699.940 1207.950 2700.000 ;
        RECT 1217.780 2699.940 1218.070 2700.000 ;
        RECT 1228.360 2699.940 1228.650 2700.000 ;
        RECT 1238.940 2699.940 1239.230 2700.000 ;
        RECT 1249.060 2699.940 1249.350 2700.000 ;
        RECT 1259.640 2699.940 1259.930 2700.000 ;
        RECT 1269.760 2699.940 1270.050 2700.000 ;
        RECT 1280.340 2699.940 1280.630 2700.000 ;
        RECT 1290.460 2699.940 1290.750 2700.000 ;
        RECT 1301.040 2699.940 1301.330 2700.000 ;
        RECT 1311.160 2699.940 1311.450 2700.000 ;
        RECT 1321.740 2699.940 1322.030 2700.000 ;
        RECT 1332.320 2699.940 1332.610 2700.000 ;
        RECT 1342.440 2699.940 1342.730 2700.000 ;
        RECT 1353.020 2699.940 1353.310 2700.000 ;
        RECT 1363.140 2699.940 1363.430 2700.000 ;
        RECT 1373.720 2699.940 1374.010 2700.000 ;
        RECT 1383.840 2699.940 1384.130 2700.000 ;
        RECT 1394.420 2699.940 1394.710 2700.000 ;
        RECT 1124.410 2696.000 1124.690 2699.870 ;
        RECT 1134.990 2696.000 1135.270 2699.940 ;
        RECT 1145.570 2696.000 1145.850 2699.940 ;
        RECT 1155.690 2696.000 1155.970 2699.940 ;
        RECT 1166.270 2696.000 1166.550 2699.940 ;
        RECT 1176.390 2696.000 1176.670 2699.940 ;
        RECT 1186.970 2696.000 1187.250 2699.940 ;
        RECT 1197.090 2696.000 1197.370 2699.940 ;
        RECT 1207.670 2696.000 1207.950 2699.940 ;
        RECT 1217.790 2696.000 1218.070 2699.940 ;
        RECT 1228.370 2696.000 1228.650 2699.940 ;
        RECT 1238.950 2696.000 1239.230 2699.940 ;
        RECT 1249.070 2696.000 1249.350 2699.940 ;
        RECT 1259.650 2696.000 1259.930 2699.940 ;
        RECT 1269.770 2696.000 1270.050 2699.940 ;
        RECT 1280.350 2696.000 1280.630 2699.940 ;
        RECT 1290.470 2696.000 1290.750 2699.940 ;
        RECT 1301.050 2696.000 1301.330 2699.940 ;
        RECT 1311.170 2696.000 1311.450 2699.940 ;
        RECT 1321.750 2696.000 1322.030 2699.940 ;
        RECT 1332.330 2696.000 1332.610 2699.940 ;
        RECT 1342.450 2696.000 1342.730 2699.940 ;
        RECT 1353.030 2696.000 1353.310 2699.940 ;
        RECT 1363.150 2696.000 1363.430 2699.940 ;
        RECT 1373.730 2696.000 1374.010 2699.940 ;
        RECT 1383.850 2696.000 1384.130 2699.940 ;
        RECT 1394.430 2696.000 1394.710 2699.940 ;
      LAYER met2 ;
        RECT 300.090 2695.720 304.870 2696.000 ;
        RECT 305.710 2695.720 314.990 2696.000 ;
        RECT 315.830 2695.720 325.570 2696.000 ;
        RECT 326.410 2695.720 335.690 2696.000 ;
        RECT 336.530 2695.720 346.270 2696.000 ;
        RECT 347.110 2695.720 356.390 2696.000 ;
        RECT 357.230 2695.720 366.970 2696.000 ;
        RECT 367.810 2695.720 377.090 2696.000 ;
        RECT 377.930 2695.720 387.670 2696.000 ;
        RECT 388.510 2695.720 398.250 2696.000 ;
        RECT 399.090 2695.720 408.370 2696.000 ;
        RECT 409.210 2695.720 418.950 2696.000 ;
        RECT 419.790 2695.720 429.070 2696.000 ;
        RECT 429.910 2695.720 439.650 2696.000 ;
        RECT 440.490 2695.720 449.770 2696.000 ;
        RECT 450.610 2695.720 460.350 2696.000 ;
        RECT 461.190 2695.720 470.470 2696.000 ;
        RECT 471.310 2695.720 481.050 2696.000 ;
        RECT 481.890 2695.720 491.630 2696.000 ;
        RECT 492.470 2695.720 501.750 2696.000 ;
        RECT 502.590 2695.720 512.330 2696.000 ;
        RECT 513.170 2695.720 522.450 2696.000 ;
        RECT 523.290 2695.720 533.030 2696.000 ;
        RECT 533.870 2695.720 543.150 2696.000 ;
        RECT 543.990 2695.720 553.730 2696.000 ;
        RECT 554.570 2695.720 563.850 2696.000 ;
        RECT 564.690 2695.720 574.430 2696.000 ;
        RECT 575.270 2695.720 585.010 2696.000 ;
        RECT 585.850 2695.720 595.130 2696.000 ;
        RECT 595.970 2695.720 605.710 2696.000 ;
        RECT 606.550 2695.720 615.830 2696.000 ;
        RECT 616.670 2695.720 626.410 2696.000 ;
        RECT 627.250 2695.720 636.530 2696.000 ;
        RECT 637.370 2695.720 647.110 2696.000 ;
        RECT 647.950 2695.720 657.230 2696.000 ;
        RECT 658.070 2695.720 667.810 2696.000 ;
        RECT 668.650 2695.720 678.390 2696.000 ;
        RECT 679.230 2695.720 688.510 2696.000 ;
        RECT 689.350 2695.720 699.090 2696.000 ;
        RECT 699.930 2695.720 709.210 2696.000 ;
        RECT 710.050 2695.720 719.790 2696.000 ;
        RECT 720.630 2695.720 729.910 2696.000 ;
        RECT 730.750 2695.720 740.490 2696.000 ;
        RECT 741.330 2695.720 750.610 2696.000 ;
        RECT 751.450 2695.720 761.190 2696.000 ;
        RECT 762.030 2695.720 771.770 2696.000 ;
        RECT 772.610 2695.720 781.890 2696.000 ;
        RECT 782.730 2695.720 792.470 2696.000 ;
        RECT 793.310 2695.720 802.590 2696.000 ;
        RECT 803.430 2695.720 813.170 2696.000 ;
        RECT 814.010 2695.720 823.290 2696.000 ;
        RECT 824.130 2695.720 833.870 2696.000 ;
        RECT 834.710 2695.720 843.990 2696.000 ;
        RECT 844.830 2695.720 854.570 2696.000 ;
        RECT 855.410 2695.720 865.150 2696.000 ;
        RECT 865.990 2695.720 875.270 2696.000 ;
        RECT 876.110 2695.720 885.850 2696.000 ;
        RECT 886.690 2695.720 895.970 2696.000 ;
        RECT 896.810 2695.720 906.550 2696.000 ;
        RECT 907.390 2695.720 916.670 2696.000 ;
        RECT 917.510 2695.720 927.250 2696.000 ;
        RECT 928.090 2695.720 937.370 2696.000 ;
        RECT 938.210 2695.720 947.950 2696.000 ;
        RECT 948.790 2695.720 958.530 2696.000 ;
        RECT 959.370 2695.720 968.650 2696.000 ;
        RECT 969.490 2695.720 979.230 2696.000 ;
        RECT 980.070 2695.720 989.350 2696.000 ;
        RECT 990.190 2695.720 999.930 2696.000 ;
        RECT 1000.770 2695.720 1010.050 2696.000 ;
        RECT 1010.890 2695.720 1020.630 2696.000 ;
        RECT 1021.470 2695.720 1030.750 2696.000 ;
        RECT 1031.590 2695.720 1041.330 2696.000 ;
        RECT 1042.170 2695.720 1051.910 2696.000 ;
        RECT 1052.750 2695.720 1062.030 2696.000 ;
        RECT 1062.870 2695.720 1072.610 2696.000 ;
        RECT 1073.450 2695.720 1082.730 2696.000 ;
        RECT 1083.570 2695.720 1093.310 2696.000 ;
        RECT 1094.150 2695.720 1103.430 2696.000 ;
        RECT 1104.270 2695.720 1114.010 2696.000 ;
        RECT 1114.850 2695.720 1124.130 2696.000 ;
        RECT 1124.970 2695.720 1134.710 2696.000 ;
        RECT 1135.550 2695.720 1145.290 2696.000 ;
        RECT 1146.130 2695.720 1155.410 2696.000 ;
        RECT 1156.250 2695.720 1165.990 2696.000 ;
        RECT 1166.830 2695.720 1176.110 2696.000 ;
        RECT 1176.950 2695.720 1186.690 2696.000 ;
        RECT 1187.530 2695.720 1196.810 2696.000 ;
        RECT 1197.650 2695.720 1207.390 2696.000 ;
        RECT 1208.230 2695.720 1217.510 2696.000 ;
        RECT 1218.350 2695.720 1228.090 2696.000 ;
        RECT 1228.930 2695.720 1238.670 2696.000 ;
        RECT 1239.510 2695.720 1248.790 2696.000 ;
        RECT 1249.630 2695.720 1259.370 2696.000 ;
        RECT 1260.210 2695.720 1269.490 2696.000 ;
        RECT 1270.330 2695.720 1280.070 2696.000 ;
        RECT 1280.910 2695.720 1290.190 2696.000 ;
        RECT 1291.030 2695.720 1300.770 2696.000 ;
        RECT 1301.610 2695.720 1310.890 2696.000 ;
        RECT 1311.730 2695.720 1321.470 2696.000 ;
        RECT 1322.310 2695.720 1332.050 2696.000 ;
        RECT 1332.890 2695.720 1342.170 2696.000 ;
        RECT 1343.010 2695.720 1352.750 2696.000 ;
        RECT 1353.590 2695.720 1362.870 2696.000 ;
        RECT 1363.710 2695.720 1373.450 2696.000 ;
        RECT 1374.290 2695.720 1383.570 2696.000 ;
        RECT 1384.410 2695.720 1394.150 2696.000 ;
        RECT 1394.990 2695.720 1395.630 2696.000 ;
        RECT 300.090 1604.280 1395.630 2695.720 ;
      LAYER met2 ;
        RECT 1407.690 2146.915 1407.970 2147.285 ;
        RECT 1407.760 2146.070 1407.900 2146.915 ;
        RECT 1407.700 2145.750 1407.960 2146.070 ;
        RECT 1407.690 2142.155 1407.970 2142.525 ;
        RECT 1407.760 2139.270 1407.900 2142.155 ;
        RECT 1407.700 2138.950 1407.960 2139.270 ;
        RECT 1408.150 2136.715 1408.430 2137.085 ;
        RECT 1408.220 2132.810 1408.360 2136.715 ;
        RECT 1408.160 2132.490 1408.420 2132.810 ;
        RECT 1407.700 2132.325 1407.960 2132.470 ;
        RECT 1407.690 2131.955 1407.970 2132.325 ;
        RECT 1407.690 2126.515 1407.970 2126.885 ;
        RECT 1407.760 2125.670 1407.900 2126.515 ;
        RECT 1407.700 2125.350 1407.960 2125.670 ;
        RECT 1407.690 2121.755 1407.970 2122.125 ;
        RECT 1407.760 2118.530 1407.900 2121.755 ;
        RECT 1407.700 2118.210 1407.960 2118.530 ;
        RECT 1408.150 2116.995 1408.430 2117.365 ;
        RECT 1408.220 2112.070 1408.360 2116.995 ;
        RECT 1407.690 2111.555 1407.970 2111.925 ;
        RECT 1408.160 2111.750 1408.420 2112.070 ;
        RECT 1407.700 2111.410 1407.960 2111.555 ;
        RECT 1407.690 2106.795 1407.970 2107.165 ;
        RECT 1407.760 2104.930 1407.900 2106.795 ;
        RECT 1407.700 2104.610 1407.960 2104.930 ;
        RECT 1407.690 2101.355 1407.970 2101.725 ;
        RECT 1407.760 2097.790 1407.900 2101.355 ;
        RECT 1407.700 2097.470 1407.960 2097.790 ;
        RECT 1408.150 2096.595 1408.430 2096.965 ;
        RECT 1407.690 2091.155 1407.970 2091.525 ;
        RECT 1408.220 2091.330 1408.360 2096.595 ;
        RECT 1407.760 2090.990 1407.900 2091.155 ;
        RECT 1408.160 2091.010 1408.420 2091.330 ;
        RECT 1407.700 2090.670 1407.960 2090.990 ;
        RECT 1414.130 2086.395 1414.410 2086.765 ;
        RECT 1414.200 2084.190 1414.340 2086.395 ;
        RECT 1414.140 2083.870 1414.400 2084.190 ;
        RECT 1411.370 2081.635 1411.650 2082.005 ;
        RECT 1411.440 2077.390 1411.580 2081.635 ;
        RECT 1411.380 2077.070 1411.640 2077.390 ;
        RECT 1408.610 2076.195 1408.890 2076.565 ;
        RECT 1408.680 2070.590 1408.820 2076.195 ;
        RECT 1410.450 2071.435 1410.730 2071.805 ;
        RECT 1408.620 2070.270 1408.880 2070.590 ;
        RECT 1410.520 2070.250 1410.660 2071.435 ;
        RECT 1410.460 2069.930 1410.720 2070.250 ;
        RECT 1413.220 2068.230 1413.480 2068.550 ;
        RECT 1407.700 2067.890 1407.960 2068.210 ;
        RECT 1407.760 2064.210 1407.900 2067.890 ;
        RECT 1409.080 2067.210 1409.340 2067.530 ;
        RECT 1407.300 2064.070 1407.900 2064.210 ;
        RECT 1407.300 2062.170 1407.440 2064.070 ;
        RECT 1407.700 2063.470 1407.960 2063.790 ;
        RECT 1408.160 2063.470 1408.420 2063.790 ;
        RECT 1407.760 2063.110 1407.900 2063.470 ;
        RECT 1407.700 2062.790 1407.960 2063.110 ;
        RECT 1408.220 2062.850 1408.360 2063.470 ;
        RECT 1408.220 2062.710 1408.820 2062.850 ;
        RECT 1409.140 2062.770 1409.280 2067.210 ;
        RECT 1410.920 2066.530 1411.180 2066.850 ;
        RECT 1410.000 2065.170 1410.260 2065.490 ;
        RECT 1407.300 2062.030 1408.360 2062.170 ;
        RECT 1407.700 2061.430 1407.960 2061.750 ;
        RECT 1407.760 1650.090 1407.900 2061.430 ;
        RECT 1408.220 2039.310 1408.360 2062.030 ;
        RECT 1408.160 2038.990 1408.420 2039.310 ;
        RECT 1408.160 2038.310 1408.420 2038.630 ;
        RECT 1408.220 2015.250 1408.360 2038.310 ;
        RECT 1408.680 2026.245 1408.820 2062.710 ;
        RECT 1409.080 2062.450 1409.340 2062.770 ;
        RECT 1409.080 2061.770 1409.340 2062.090 ;
        RECT 1409.140 2031.005 1409.280 2061.770 ;
        RECT 1409.540 2059.730 1409.800 2060.050 ;
        RECT 1409.600 2056.650 1409.740 2059.730 ;
        RECT 1409.540 2056.330 1409.800 2056.650 ;
        RECT 1409.540 2055.650 1409.800 2055.970 ;
        RECT 1409.600 2051.405 1409.740 2055.650 ;
        RECT 1409.530 2051.035 1409.810 2051.405 ;
        RECT 1409.540 2050.550 1409.800 2050.870 ;
        RECT 1409.600 2038.630 1409.740 2050.550 ;
        RECT 1410.060 2039.050 1410.200 2065.170 ;
        RECT 1410.460 2063.810 1410.720 2064.130 ;
        RECT 1410.520 2062.090 1410.660 2063.810 ;
        RECT 1410.460 2061.770 1410.720 2062.090 ;
        RECT 1410.450 2061.235 1410.730 2061.605 ;
        RECT 1410.520 2059.030 1410.660 2061.235 ;
        RECT 1410.460 2058.710 1410.720 2059.030 ;
        RECT 1410.460 2057.690 1410.720 2058.010 ;
        RECT 1410.520 2039.650 1410.660 2057.690 ;
        RECT 1410.980 2039.650 1411.120 2066.530 ;
        RECT 1411.840 2065.510 1412.100 2065.830 ;
        RECT 1411.380 2064.490 1411.640 2064.810 ;
        RECT 1410.460 2039.330 1410.720 2039.650 ;
        RECT 1410.920 2039.330 1411.180 2039.650 ;
        RECT 1410.060 2038.910 1411.120 2039.050 ;
        RECT 1409.540 2038.310 1409.800 2038.630 ;
        RECT 1410.000 2038.370 1410.260 2038.630 ;
        RECT 1410.000 2038.310 1410.660 2038.370 ;
        RECT 1410.060 2038.230 1410.660 2038.310 ;
        RECT 1409.540 2037.630 1409.800 2037.950 ;
        RECT 1410.000 2037.630 1410.260 2037.950 ;
        RECT 1409.070 2030.635 1409.350 2031.005 ;
        RECT 1408.610 2025.875 1408.890 2026.245 ;
        RECT 1409.600 2016.045 1409.740 2037.630 ;
        RECT 1409.530 2015.675 1409.810 2016.045 ;
        RECT 1408.220 2015.110 1409.740 2015.250 ;
        RECT 1408.160 2005.845 1408.420 2005.990 ;
        RECT 1408.150 2005.475 1408.430 2005.845 ;
        RECT 1408.150 2000.715 1408.430 2001.085 ;
        RECT 1408.160 2000.570 1408.420 2000.715 ;
        RECT 1408.160 1997.510 1408.420 1997.830 ;
        RECT 1408.220 1995.645 1408.360 1997.510 ;
        RECT 1408.150 1995.275 1408.430 1995.645 ;
        RECT 1408.160 1972.690 1408.420 1973.010 ;
        RECT 1408.220 1970.485 1408.360 1972.690 ;
        RECT 1408.150 1970.115 1408.430 1970.485 ;
        RECT 1408.610 1966.035 1408.890 1966.405 ;
        RECT 1408.160 1965.725 1408.420 1965.870 ;
        RECT 1408.150 1965.355 1408.430 1965.725 ;
        RECT 1408.160 1961.810 1408.420 1962.130 ;
        RECT 1408.220 1960.285 1408.360 1961.810 ;
        RECT 1408.150 1959.915 1408.430 1960.285 ;
        RECT 1408.160 1940.730 1408.420 1941.050 ;
        RECT 1408.220 1940.565 1408.360 1940.730 ;
        RECT 1408.150 1940.195 1408.430 1940.565 ;
        RECT 1408.160 1935.125 1408.420 1935.270 ;
        RECT 1408.150 1934.755 1408.430 1935.125 ;
        RECT 1408.680 1930.930 1408.820 1966.035 ;
        RECT 1409.080 1965.890 1409.340 1966.210 ;
        RECT 1408.220 1930.790 1408.820 1930.930 ;
        RECT 1408.220 1928.890 1408.360 1930.790 ;
        RECT 1408.620 1930.365 1408.880 1930.510 ;
        RECT 1408.610 1929.995 1408.890 1930.365 ;
        RECT 1408.220 1928.750 1408.820 1928.890 ;
        RECT 1408.160 1927.810 1408.420 1928.130 ;
        RECT 1408.220 1925.605 1408.360 1927.810 ;
        RECT 1408.150 1925.235 1408.430 1925.605 ;
        RECT 1408.160 1924.410 1408.420 1924.730 ;
        RECT 1408.220 1920.165 1408.360 1924.410 ;
        RECT 1408.150 1919.795 1408.430 1920.165 ;
        RECT 1408.680 1919.290 1408.820 1928.750 ;
        RECT 1408.620 1918.970 1408.880 1919.290 ;
        RECT 1409.140 1918.950 1409.280 1965.890 ;
        RECT 1409.600 1950.765 1409.740 2015.110 ;
        RECT 1409.530 1950.395 1409.810 1950.765 ;
        RECT 1409.080 1918.630 1409.340 1918.950 ;
        RECT 1408.620 1910.810 1408.880 1911.130 ;
        RECT 1408.160 1909.965 1408.420 1910.110 ;
        RECT 1408.150 1909.595 1408.430 1909.965 ;
        RECT 1408.680 1905.205 1408.820 1910.810 ;
        RECT 1408.610 1904.835 1408.890 1905.205 ;
        RECT 1409.540 1869.670 1409.800 1869.990 ;
        RECT 1409.080 1868.990 1409.340 1869.310 ;
        RECT 1408.620 1868.650 1408.880 1868.970 ;
        RECT 1408.680 1822.730 1408.820 1868.650 ;
        RECT 1408.620 1822.410 1408.880 1822.730 ;
        RECT 1409.140 1822.390 1409.280 1868.990 ;
        RECT 1409.080 1822.070 1409.340 1822.390 ;
        RECT 1409.600 1822.050 1409.740 1869.670 ;
        RECT 1409.540 1821.730 1409.800 1822.050 ;
        RECT 1408.620 1807.450 1408.880 1807.770 ;
        RECT 1408.680 1803.885 1408.820 1807.450 ;
        RECT 1408.610 1803.515 1408.890 1803.885 ;
        RECT 1409.540 1793.510 1409.800 1793.830 ;
        RECT 1409.600 1788.925 1409.740 1793.510 ;
        RECT 1409.530 1788.555 1409.810 1788.925 ;
        RECT 1410.060 1784.165 1410.200 2037.630 ;
        RECT 1409.990 1783.795 1410.270 1784.165 ;
        RECT 1410.520 1778.725 1410.660 2038.230 ;
        RECT 1410.980 2013.890 1411.120 2038.910 ;
        RECT 1411.440 2014.490 1411.580 2064.490 ;
        RECT 1411.900 2039.050 1412.040 2065.510 ;
        RECT 1412.300 2064.830 1412.560 2065.150 ;
        RECT 1412.360 2057.410 1412.500 2064.830 ;
        RECT 1412.360 2057.270 1412.960 2057.410 ;
        RECT 1412.300 2056.670 1412.560 2056.990 ;
        RECT 1412.360 2039.845 1412.500 2056.670 ;
        RECT 1412.290 2039.475 1412.570 2039.845 ;
        RECT 1411.900 2038.910 1412.500 2039.050 ;
        RECT 1411.380 2014.170 1411.640 2014.490 ;
        RECT 1410.980 2013.750 1412.040 2013.890 ;
        RECT 1411.380 2013.150 1411.640 2013.470 ;
        RECT 1410.920 2012.810 1411.180 2013.130 ;
        RECT 1410.980 2011.285 1411.120 2012.810 ;
        RECT 1410.910 2010.915 1411.190 2011.285 ;
        RECT 1410.920 1990.885 1411.180 1991.030 ;
        RECT 1410.910 1990.515 1411.190 1990.885 ;
        RECT 1410.920 1966.230 1411.180 1966.550 ;
        RECT 1410.980 1918.610 1411.120 1966.230 ;
        RECT 1410.920 1918.290 1411.180 1918.610 ;
        RECT 1410.920 1890.070 1411.180 1890.390 ;
        RECT 1410.980 1884.805 1411.120 1890.070 ;
        RECT 1410.910 1884.435 1411.190 1884.805 ;
        RECT 1410.920 1869.330 1411.180 1869.650 ;
        RECT 1410.980 1864.405 1411.120 1869.330 ;
        RECT 1410.910 1864.035 1411.190 1864.405 ;
        RECT 1410.920 1855.390 1411.180 1855.710 ;
        RECT 1410.980 1849.445 1411.120 1855.390 ;
        RECT 1410.910 1849.075 1411.190 1849.445 ;
        RECT 1410.920 1834.650 1411.180 1834.970 ;
        RECT 1410.980 1829.045 1411.120 1834.650 ;
        RECT 1410.910 1828.675 1411.190 1829.045 ;
        RECT 1410.920 1814.590 1411.180 1814.910 ;
        RECT 1410.450 1778.355 1410.730 1778.725 ;
        RECT 1410.980 1773.965 1411.120 1814.590 ;
        RECT 1410.910 1773.595 1411.190 1773.965 ;
        RECT 1409.990 1772.915 1410.270 1773.285 ;
        RECT 1410.060 1759.005 1410.200 1772.915 ;
        RECT 1410.460 1772.770 1410.720 1773.090 ;
        RECT 1410.520 1763.765 1410.660 1772.770 ;
        RECT 1410.450 1763.395 1410.730 1763.765 ;
        RECT 1409.990 1758.635 1410.270 1759.005 ;
        RECT 1411.440 1748.805 1411.580 2013.150 ;
        RECT 1411.900 1966.210 1412.040 2013.750 ;
        RECT 1412.360 1966.405 1412.500 2038.910 ;
        RECT 1412.820 1966.550 1412.960 2057.270 ;
        RECT 1413.280 2040.410 1413.420 2068.230 ;
        RECT 1414.140 2066.365 1414.400 2066.510 ;
        RECT 1414.130 2065.995 1414.410 2066.365 ;
        RECT 1413.680 2064.150 1413.940 2064.470 ;
        RECT 1413.740 2062.850 1413.880 2064.150 ;
        RECT 1413.740 2062.710 1414.340 2062.850 ;
        RECT 1413.680 2062.110 1413.940 2062.430 ;
        RECT 1413.740 2041.090 1413.880 2062.110 ;
        RECT 1414.200 2056.990 1414.340 2062.710 ;
        RECT 1417.360 2060.750 1417.620 2061.070 ;
        RECT 1416.900 2060.410 1417.160 2060.730 ;
        RECT 1414.600 2060.070 1414.860 2060.390 ;
        RECT 1414.140 2056.670 1414.400 2056.990 ;
        RECT 1414.140 2056.165 1414.400 2056.310 ;
        RECT 1414.130 2055.795 1414.410 2056.165 ;
        RECT 1414.660 2055.370 1414.800 2060.070 ;
        RECT 1415.060 2058.370 1415.320 2058.690 ;
        RECT 1414.200 2055.230 1414.800 2055.370 ;
        RECT 1414.200 2041.770 1414.340 2055.230 ;
        RECT 1414.600 2052.930 1414.860 2053.250 ;
        RECT 1414.660 2042.565 1414.800 2052.930 ;
        RECT 1415.120 2046.645 1415.260 2058.370 ;
        RECT 1415.520 2057.350 1415.780 2057.670 ;
        RECT 1415.050 2046.275 1415.330 2046.645 ;
        RECT 1414.590 2042.195 1414.870 2042.565 ;
        RECT 1414.200 2041.630 1415.260 2041.770 ;
        RECT 1413.740 2040.950 1414.340 2041.090 ;
        RECT 1413.280 2040.270 1413.880 2040.410 ;
        RECT 1413.220 2039.330 1413.480 2039.650 ;
        RECT 1411.840 1965.890 1412.100 1966.210 ;
        RECT 1412.290 1966.035 1412.570 1966.405 ;
        RECT 1412.760 1966.230 1413.020 1966.550 ;
        RECT 1411.840 1918.630 1412.100 1918.950 ;
        RECT 1412.300 1918.630 1412.560 1918.950 ;
        RECT 1411.900 1869.310 1412.040 1918.630 ;
        RECT 1412.360 1869.310 1412.500 1918.630 ;
        RECT 1412.760 1918.290 1413.020 1918.610 ;
        RECT 1412.820 1869.990 1412.960 1918.290 ;
        RECT 1412.760 1869.670 1413.020 1869.990 ;
        RECT 1411.840 1868.990 1412.100 1869.310 ;
        RECT 1412.300 1868.990 1412.560 1869.310 ;
        RECT 1411.840 1822.070 1412.100 1822.390 ;
        RECT 1412.300 1822.070 1412.560 1822.390 ;
        RECT 1411.900 1773.285 1412.040 1822.070 ;
        RECT 1411.830 1772.915 1412.110 1773.285 ;
        RECT 1412.360 1773.090 1412.500 1822.070 ;
        RECT 1412.760 1821.730 1413.020 1822.050 ;
        RECT 1412.300 1772.770 1412.560 1773.090 ;
        RECT 1412.820 1753.565 1412.960 1821.730 ;
        RECT 1413.280 1768.525 1413.420 2039.330 ;
        RECT 1413.740 2037.950 1413.880 2040.270 ;
        RECT 1413.680 2037.630 1413.940 2037.950 ;
        RECT 1414.200 2037.010 1414.340 2040.950 ;
        RECT 1413.740 2036.870 1414.340 2037.010 ;
        RECT 1413.740 1814.910 1413.880 2036.870 ;
        RECT 1415.120 2036.330 1415.260 2041.630 ;
        RECT 1414.200 2036.190 1415.260 2036.330 ;
        RECT 1414.200 2022.050 1414.340 2036.190 ;
        RECT 1414.200 2021.910 1414.800 2022.050 ;
        RECT 1414.140 2021.485 1414.400 2021.630 ;
        RECT 1414.130 2021.115 1414.410 2021.485 ;
        RECT 1414.660 2020.690 1414.800 2021.910 ;
        RECT 1414.200 2020.550 1414.800 2020.690 ;
        RECT 1414.200 1945.325 1414.340 2020.550 ;
        RECT 1415.580 2005.990 1415.720 2057.350 ;
        RECT 1416.440 2057.010 1416.700 2057.330 ;
        RECT 1415.980 2056.330 1416.240 2056.650 ;
        RECT 1415.520 2005.670 1415.780 2005.990 ;
        RECT 1416.040 1997.830 1416.180 2056.330 ;
        RECT 1416.500 2000.890 1416.640 2057.010 ;
        RECT 1416.440 2000.570 1416.700 2000.890 ;
        RECT 1415.980 1997.510 1416.240 1997.830 ;
        RECT 1414.130 1944.955 1414.410 1945.325 ;
        RECT 1416.960 1941.050 1417.100 2060.410 ;
        RECT 1416.900 1940.730 1417.160 1941.050 ;
        RECT 1417.420 1935.270 1417.560 2060.750 ;
        RECT 1417.880 1965.870 1418.020 2788.010 ;
        RECT 1417.820 1965.550 1418.080 1965.870 ;
        RECT 1418.340 1962.130 1418.480 2788.350 ;
        RECT 1418.800 1973.010 1418.940 2790.390 ;
        RECT 1420.580 2061.770 1420.840 2062.090 ;
        RECT 1420.120 2061.430 1420.380 2061.750 ;
        RECT 1419.660 2053.270 1419.920 2053.590 ;
        RECT 1419.200 2052.590 1419.460 2052.910 ;
        RECT 1418.740 1972.690 1419.000 1973.010 ;
        RECT 1418.280 1961.810 1418.540 1962.130 ;
        RECT 1417.360 1934.950 1417.620 1935.270 ;
        RECT 1414.140 1917.950 1414.400 1918.270 ;
        RECT 1414.200 1915.405 1414.340 1917.950 ;
        RECT 1414.130 1915.035 1414.410 1915.405 ;
        RECT 1414.140 1904.010 1414.400 1904.330 ;
        RECT 1414.200 1899.765 1414.340 1904.010 ;
        RECT 1414.130 1899.395 1414.410 1899.765 ;
        RECT 1414.140 1897.210 1414.400 1897.530 ;
        RECT 1414.200 1895.005 1414.340 1897.210 ;
        RECT 1414.130 1894.635 1414.410 1895.005 ;
        RECT 1414.140 1890.410 1414.400 1890.730 ;
        RECT 1414.200 1890.245 1414.340 1890.410 ;
        RECT 1414.130 1889.875 1414.410 1890.245 ;
        RECT 1414.140 1883.270 1414.400 1883.590 ;
        RECT 1414.200 1880.045 1414.340 1883.270 ;
        RECT 1414.130 1879.675 1414.410 1880.045 ;
        RECT 1414.140 1876.470 1414.400 1876.790 ;
        RECT 1414.200 1874.605 1414.340 1876.470 ;
        RECT 1414.130 1874.235 1414.410 1874.605 ;
        RECT 1414.140 1869.845 1414.400 1869.990 ;
        RECT 1414.130 1869.475 1414.410 1869.845 ;
        RECT 1414.140 1862.530 1414.400 1862.850 ;
        RECT 1414.200 1859.645 1414.340 1862.530 ;
        RECT 1414.130 1859.275 1414.410 1859.645 ;
        RECT 1414.140 1855.730 1414.400 1856.050 ;
        RECT 1414.200 1854.885 1414.340 1855.730 ;
        RECT 1414.130 1854.515 1414.410 1854.885 ;
        RECT 1414.140 1848.930 1414.400 1849.250 ;
        RECT 1414.200 1844.685 1414.340 1848.930 ;
        RECT 1414.130 1844.315 1414.410 1844.685 ;
        RECT 1414.140 1842.130 1414.400 1842.450 ;
        RECT 1414.200 1839.245 1414.340 1842.130 ;
        RECT 1414.130 1838.875 1414.410 1839.245 ;
        RECT 1414.140 1834.990 1414.400 1835.310 ;
        RECT 1414.200 1834.485 1414.340 1834.990 ;
        RECT 1414.130 1834.115 1414.410 1834.485 ;
        RECT 1414.140 1828.190 1414.400 1828.510 ;
        RECT 1414.200 1824.285 1414.340 1828.190 ;
        RECT 1414.130 1823.915 1414.410 1824.285 ;
        RECT 1414.140 1821.390 1414.400 1821.710 ;
        RECT 1414.200 1819.525 1414.340 1821.390 ;
        RECT 1414.130 1819.155 1414.410 1819.525 ;
        RECT 1413.680 1814.590 1413.940 1814.910 ;
        RECT 1414.140 1814.250 1414.400 1814.570 ;
        RECT 1413.680 1813.910 1413.940 1814.230 ;
        RECT 1414.200 1814.085 1414.340 1814.250 ;
        RECT 1413.740 1809.325 1413.880 1813.910 ;
        RECT 1414.130 1813.715 1414.410 1814.085 ;
        RECT 1413.670 1808.955 1413.950 1809.325 ;
        RECT 1414.140 1800.650 1414.400 1800.970 ;
        RECT 1413.680 1800.310 1413.940 1800.630 ;
        RECT 1413.740 1794.365 1413.880 1800.310 ;
        RECT 1414.200 1799.125 1414.340 1800.650 ;
        RECT 1414.130 1798.755 1414.410 1799.125 ;
        RECT 1413.670 1793.995 1413.950 1794.365 ;
        RECT 1413.210 1768.155 1413.490 1768.525 ;
        RECT 1412.750 1753.195 1413.030 1753.565 ;
        RECT 1411.370 1748.435 1411.650 1748.805 ;
        RECT 1414.140 1745.230 1414.400 1745.550 ;
        RECT 1414.200 1743.365 1414.340 1745.230 ;
        RECT 1414.130 1742.995 1414.410 1743.365 ;
        RECT 1414.140 1738.605 1414.400 1738.750 ;
        RECT 1411.380 1738.090 1411.640 1738.410 ;
        RECT 1414.130 1738.235 1414.410 1738.605 ;
        RECT 1411.440 1733.165 1411.580 1738.090 ;
        RECT 1411.370 1732.795 1411.650 1733.165 ;
        RECT 1410.460 1731.630 1410.720 1731.950 ;
        RECT 1410.520 1728.405 1410.660 1731.630 ;
        RECT 1410.450 1728.035 1410.730 1728.405 ;
        RECT 1414.130 1723.275 1414.410 1723.645 ;
        RECT 1414.200 1722.770 1414.340 1723.275 ;
        RECT 1414.140 1722.450 1414.400 1722.770 ;
        RECT 1412.760 1717.690 1413.020 1718.010 ;
        RECT 1413.670 1717.835 1413.950 1718.205 ;
        RECT 1412.820 1713.445 1412.960 1717.690 ;
        RECT 1413.740 1717.670 1413.880 1717.835 ;
        RECT 1413.680 1717.350 1413.940 1717.670 ;
        RECT 1412.750 1713.075 1413.030 1713.445 ;
        RECT 1414.140 1710.890 1414.400 1711.210 ;
        RECT 1414.200 1708.005 1414.340 1710.890 ;
        RECT 1414.130 1707.635 1414.410 1708.005 ;
        RECT 1412.290 1702.875 1412.570 1703.245 ;
        RECT 1410.450 1698.115 1410.730 1698.485 ;
        RECT 1409.990 1682.475 1410.270 1682.845 ;
        RECT 1409.070 1672.275 1409.350 1672.645 ;
        RECT 1408.160 1667.885 1408.420 1668.030 ;
        RECT 1408.150 1667.515 1408.430 1667.885 ;
        RECT 1408.160 1655.810 1408.420 1656.130 ;
        RECT 1408.220 1652.925 1408.360 1655.810 ;
        RECT 1408.150 1652.555 1408.430 1652.925 ;
        RECT 1407.760 1649.950 1408.820 1650.090 ;
        RECT 1408.160 1648.670 1408.420 1648.990 ;
        RECT 1407.700 1648.330 1407.960 1648.650 ;
        RECT 1407.760 1647.485 1407.900 1648.330 ;
        RECT 1407.690 1647.115 1407.970 1647.485 ;
        RECT 1408.220 1642.725 1408.360 1648.670 ;
        RECT 1408.150 1642.355 1408.430 1642.725 ;
        RECT 1407.700 1641.870 1407.960 1642.190 ;
        RECT 1407.760 1637.285 1407.900 1641.870 ;
        RECT 1407.690 1636.915 1407.970 1637.285 ;
        RECT 1407.700 1635.070 1407.960 1635.390 ;
        RECT 1407.760 1632.525 1407.900 1635.070 ;
        RECT 1407.690 1632.155 1407.970 1632.525 ;
        RECT 1407.700 1627.930 1407.960 1628.250 ;
        RECT 1407.760 1622.325 1407.900 1627.930 ;
        RECT 1408.680 1627.765 1408.820 1649.950 ;
        RECT 1409.140 1631.650 1409.280 1672.275 ;
        RECT 1410.060 1659.190 1410.200 1682.475 ;
        RECT 1410.000 1658.870 1410.260 1659.190 ;
        RECT 1409.530 1657.315 1409.810 1657.685 ;
        RECT 1409.600 1631.990 1409.740 1657.315 ;
        RECT 1410.520 1633.090 1410.660 1698.115 ;
        RECT 1411.830 1692.675 1412.110 1693.045 ;
        RECT 1410.920 1669.410 1411.180 1669.730 ;
        RECT 1410.980 1663.125 1411.120 1669.410 ;
        RECT 1410.910 1662.755 1411.190 1663.125 ;
        RECT 1410.060 1632.950 1410.660 1633.090 ;
        RECT 1409.540 1631.670 1409.800 1631.990 ;
        RECT 1409.080 1631.330 1409.340 1631.650 ;
        RECT 1408.610 1627.395 1408.890 1627.765 ;
        RECT 1407.690 1621.955 1407.970 1622.325 ;
        RECT 1407.700 1621.130 1407.960 1621.450 ;
        RECT 1407.760 1617.565 1407.900 1621.130 ;
        RECT 1407.690 1617.195 1407.970 1617.565 ;
        RECT 1407.700 1614.330 1407.960 1614.650 ;
        RECT 1407.760 1612.125 1407.900 1614.330 ;
        RECT 1407.690 1611.755 1407.970 1612.125 ;
      LAYER met2 ;
        RECT 300.090 1602.195 304.410 1604.280 ;
        RECT 305.250 1602.195 314.070 1604.280 ;
        RECT 314.910 1602.195 323.730 1604.280 ;
        RECT 324.570 1602.195 333.390 1604.280 ;
        RECT 334.230 1602.195 343.050 1604.280 ;
        RECT 343.890 1602.195 352.710 1604.280 ;
        RECT 353.550 1602.195 362.370 1604.280 ;
        RECT 363.210 1602.195 372.490 1604.280 ;
        RECT 373.330 1602.195 382.150 1604.280 ;
        RECT 382.990 1602.195 391.810 1604.280 ;
        RECT 392.650 1602.195 401.470 1604.280 ;
        RECT 402.310 1602.195 411.130 1604.280 ;
        RECT 411.970 1602.195 420.790 1604.280 ;
        RECT 421.630 1602.195 430.910 1604.280 ;
        RECT 431.750 1602.195 440.570 1604.280 ;
        RECT 441.410 1602.195 450.230 1604.280 ;
        RECT 451.070 1602.195 459.890 1604.280 ;
        RECT 460.730 1602.195 469.550 1604.280 ;
        RECT 470.390 1602.195 479.210 1604.280 ;
        RECT 480.050 1602.195 489.330 1604.280 ;
        RECT 490.170 1602.195 498.990 1604.280 ;
        RECT 499.830 1602.195 508.650 1604.280 ;
        RECT 509.490 1602.195 518.310 1604.280 ;
        RECT 519.150 1602.195 527.970 1604.280 ;
        RECT 528.810 1602.195 537.630 1604.280 ;
        RECT 538.470 1602.195 547.290 1604.280 ;
        RECT 548.130 1602.195 557.410 1604.280 ;
        RECT 558.250 1602.195 567.070 1604.280 ;
        RECT 567.910 1602.195 576.730 1604.280 ;
        RECT 577.570 1602.195 586.390 1604.280 ;
        RECT 587.230 1602.195 596.050 1604.280 ;
        RECT 596.890 1602.195 605.710 1604.280 ;
        RECT 606.550 1602.195 615.830 1604.280 ;
        RECT 616.670 1602.195 625.490 1604.280 ;
        RECT 626.330 1602.195 635.150 1604.280 ;
        RECT 635.990 1602.195 644.810 1604.280 ;
        RECT 645.650 1602.195 654.470 1604.280 ;
        RECT 655.310 1602.195 664.130 1604.280 ;
        RECT 664.970 1602.195 674.250 1604.280 ;
        RECT 675.090 1602.195 683.910 1604.280 ;
        RECT 684.750 1602.195 693.570 1604.280 ;
        RECT 694.410 1602.195 703.230 1604.280 ;
        RECT 704.070 1602.195 712.890 1604.280 ;
        RECT 713.730 1602.195 722.550 1604.280 ;
        RECT 723.390 1602.195 732.670 1604.280 ;
        RECT 733.510 1602.195 742.330 1604.280 ;
        RECT 743.170 1602.195 751.990 1604.280 ;
        RECT 752.830 1602.195 761.650 1604.280 ;
        RECT 762.490 1602.195 771.310 1604.280 ;
        RECT 772.150 1602.195 780.970 1604.280 ;
        RECT 781.810 1602.195 790.630 1604.280 ;
        RECT 791.470 1602.195 800.750 1604.280 ;
        RECT 801.590 1602.195 810.410 1604.280 ;
        RECT 811.250 1602.195 820.070 1604.280 ;
        RECT 820.910 1602.195 829.730 1604.280 ;
        RECT 830.570 1602.195 839.390 1604.280 ;
        RECT 840.230 1602.195 849.050 1604.280 ;
        RECT 849.890 1602.195 859.170 1604.280 ;
        RECT 860.010 1602.195 868.830 1604.280 ;
        RECT 869.670 1602.195 878.490 1604.280 ;
        RECT 879.330 1602.195 888.150 1604.280 ;
        RECT 888.990 1602.195 897.810 1604.280 ;
        RECT 898.650 1602.195 907.470 1604.280 ;
        RECT 908.310 1602.195 917.590 1604.280 ;
        RECT 918.430 1602.195 927.250 1604.280 ;
        RECT 928.090 1602.195 936.910 1604.280 ;
        RECT 937.750 1602.195 946.570 1604.280 ;
        RECT 947.410 1602.195 956.230 1604.280 ;
        RECT 957.070 1602.195 965.890 1604.280 ;
        RECT 966.730 1602.195 975.550 1604.280 ;
        RECT 976.390 1602.195 985.670 1604.280 ;
        RECT 986.510 1602.195 995.330 1604.280 ;
        RECT 996.170 1602.195 1004.990 1604.280 ;
        RECT 1005.830 1602.195 1014.650 1604.280 ;
        RECT 1015.490 1602.195 1024.310 1604.280 ;
        RECT 1025.150 1602.195 1033.970 1604.280 ;
        RECT 1034.810 1602.195 1044.090 1604.280 ;
        RECT 1044.930 1602.195 1053.750 1604.280 ;
        RECT 1054.590 1602.195 1063.410 1604.280 ;
        RECT 1064.250 1602.195 1073.070 1604.280 ;
        RECT 1073.910 1602.195 1082.730 1604.280 ;
        RECT 1083.570 1602.195 1092.390 1604.280 ;
        RECT 1093.230 1602.195 1102.510 1604.280 ;
        RECT 1103.350 1602.195 1112.170 1604.280 ;
        RECT 1113.010 1602.195 1121.830 1604.280 ;
        RECT 1122.670 1602.195 1131.490 1604.280 ;
        RECT 1132.330 1602.195 1141.150 1604.280 ;
        RECT 1141.990 1602.195 1150.810 1604.280 ;
        RECT 1151.650 1602.195 1160.930 1604.280 ;
        RECT 1161.770 1602.195 1170.590 1604.280 ;
        RECT 1171.430 1602.195 1180.250 1604.280 ;
        RECT 1181.090 1602.195 1189.910 1604.280 ;
        RECT 1190.750 1602.195 1199.570 1604.280 ;
        RECT 1200.410 1602.195 1209.230 1604.280 ;
        RECT 1210.070 1602.195 1218.890 1604.280 ;
        RECT 1219.730 1602.195 1229.010 1604.280 ;
        RECT 1229.850 1602.195 1238.670 1604.280 ;
        RECT 1239.510 1602.195 1248.330 1604.280 ;
        RECT 1249.170 1602.195 1257.990 1604.280 ;
        RECT 1258.830 1602.195 1267.650 1604.280 ;
        RECT 1268.490 1602.195 1277.310 1604.280 ;
        RECT 1278.150 1602.195 1287.430 1604.280 ;
        RECT 1288.270 1602.195 1297.090 1604.280 ;
        RECT 1297.930 1602.195 1306.750 1604.280 ;
        RECT 1307.590 1602.195 1316.410 1604.280 ;
        RECT 1317.250 1602.195 1326.070 1604.280 ;
        RECT 1326.910 1602.195 1335.730 1604.280 ;
        RECT 1336.570 1602.195 1345.850 1604.280 ;
        RECT 1346.690 1602.195 1355.510 1604.280 ;
        RECT 1356.350 1602.195 1365.170 1604.280 ;
        RECT 1366.010 1602.195 1374.830 1604.280 ;
        RECT 1375.670 1602.195 1384.490 1604.280 ;
        RECT 1385.330 1602.195 1394.150 1604.280 ;
        RECT 1394.990 1602.195 1395.630 1604.280 ;
      LAYER met2 ;
        RECT 1410.060 1602.750 1410.200 1632.950 ;
        RECT 1410.460 1632.010 1410.720 1632.330 ;
        RECT 1410.000 1602.430 1410.260 1602.750 ;
        RECT 1410.520 1601.390 1410.660 1632.010 ;
        RECT 1410.920 1631.670 1411.180 1631.990 ;
        RECT 1411.380 1631.670 1411.640 1631.990 ;
        RECT 1410.980 1604.790 1411.120 1631.670 ;
        RECT 1410.920 1604.470 1411.180 1604.790 ;
        RECT 1411.440 1602.070 1411.580 1631.670 ;
        RECT 1411.900 1603.090 1412.040 1692.675 ;
        RECT 1411.840 1602.770 1412.100 1603.090 ;
        RECT 1412.360 1602.410 1412.500 1702.875 ;
        RECT 1412.750 1687.915 1413.030 1688.285 ;
        RECT 1412.820 1604.450 1412.960 1687.915 ;
        RECT 1413.210 1677.715 1413.490 1678.085 ;
        RECT 1413.280 1631.990 1413.420 1677.715 ;
        RECT 1419.260 1668.030 1419.400 2052.590 ;
        RECT 1419.720 1910.110 1419.860 2053.270 ;
        RECT 1420.180 1924.730 1420.320 2061.430 ;
        RECT 1420.640 1928.130 1420.780 2061.770 ;
        RECT 1421.040 2061.090 1421.300 2061.410 ;
        RECT 1421.100 1930.510 1421.240 2061.090 ;
        RECT 1425.180 2058.030 1425.440 2058.350 ;
        RECT 1424.720 2056.670 1424.980 2056.990 ;
        RECT 1424.780 1991.030 1424.920 2056.670 ;
        RECT 1425.240 2013.130 1425.380 2058.030 ;
        RECT 1425.180 2012.810 1425.440 2013.130 ;
        RECT 1424.720 1990.710 1424.980 1991.030 ;
        RECT 1421.040 1930.190 1421.300 1930.510 ;
        RECT 1420.580 1927.810 1420.840 1928.130 ;
        RECT 1420.120 1924.410 1420.380 1924.730 ;
        RECT 1419.660 1909.790 1419.920 1910.110 ;
        RECT 1419.200 1667.710 1419.460 1668.030 ;
        RECT 1413.680 1658.870 1413.940 1659.190 ;
        RECT 1413.740 1632.330 1413.880 1658.870 ;
        RECT 1413.680 1632.010 1413.940 1632.330 ;
        RECT 1413.220 1631.670 1413.480 1631.990 ;
        RECT 1413.680 1631.330 1413.940 1631.650 ;
        RECT 1412.760 1604.130 1413.020 1604.450 ;
        RECT 1412.300 1602.090 1412.560 1602.410 ;
        RECT 1411.380 1601.750 1411.640 1602.070 ;
        RECT 1413.740 1601.730 1413.880 1631.330 ;
        RECT 1428.000 1611.250 1428.140 3250.750 ;
        RECT 1535.570 3231.515 1535.850 3231.885 ;
        RECT 1535.640 3229.650 1535.780 3231.515 ;
        RECT 1486.820 3229.330 1487.080 3229.650 ;
        RECT 1535.580 3229.330 1535.840 3229.650 ;
        RECT 1473.020 3222.190 1473.280 3222.510 ;
        RECT 1459.220 3215.390 1459.480 3215.710 ;
        RECT 1452.320 3208.590 1452.580 3208.910 ;
        RECT 1438.520 3201.450 1438.780 3201.770 ;
        RECT 1431.620 3194.650 1431.880 3194.970 ;
        RECT 1431.680 1717.670 1431.820 3194.650 ;
        RECT 1435.760 2066.870 1436.020 2067.190 ;
        RECT 1435.300 2065.850 1435.560 2066.170 ;
        RECT 1435.360 2065.150 1435.500 2065.850 ;
        RECT 1435.820 2065.490 1435.960 2066.870 ;
        RECT 1435.760 2065.170 1436.020 2065.490 ;
        RECT 1435.300 2064.830 1435.560 2065.150 ;
        RECT 1438.580 1722.770 1438.720 3201.450 ;
        RECT 1452.380 1731.950 1452.520 3208.590 ;
        RECT 1459.280 1738.410 1459.420 3215.390 ;
        RECT 1473.080 1738.750 1473.220 3222.190 ;
        RECT 1482.680 2066.870 1482.940 2067.190 ;
        RECT 1482.740 2065.490 1482.880 2066.870 ;
        RECT 1483.140 2065.850 1483.400 2066.170 ;
        RECT 1482.680 2065.170 1482.940 2065.490 ;
        RECT 1483.200 2065.150 1483.340 2065.850 ;
        RECT 1483.140 2064.830 1483.400 2065.150 ;
        RECT 1486.880 1745.550 1487.020 3229.330 ;
        RECT 1535.570 3224.715 1535.850 3225.085 ;
        RECT 1535.640 3222.510 1535.780 3224.715 ;
        RECT 1535.580 3222.190 1535.840 3222.510 ;
        RECT 1535.570 3217.235 1535.850 3217.605 ;
        RECT 1535.640 3215.710 1535.780 3217.235 ;
        RECT 1535.580 3215.390 1535.840 3215.710 ;
        RECT 1538.330 3210.435 1538.610 3210.805 ;
        RECT 1538.400 3208.910 1538.540 3210.435 ;
        RECT 1538.340 3208.590 1538.600 3208.910 ;
        RECT 1538.330 3202.275 1538.610 3202.645 ;
        RECT 1538.400 3201.770 1538.540 3202.275 ;
        RECT 1538.340 3201.450 1538.600 3201.770 ;
        RECT 1533.270 3196.835 1533.550 3197.205 ;
        RECT 1533.340 3194.970 1533.480 3196.835 ;
        RECT 1533.280 3194.650 1533.540 3194.970 ;
        RECT 1534.190 3189.355 1534.470 3189.725 ;
        RECT 1534.260 3188.170 1534.400 3189.355 ;
        RECT 1507.520 3187.850 1507.780 3188.170 ;
        RECT 1534.200 3187.850 1534.460 3188.170 ;
        RECT 1487.280 2789.030 1487.540 2789.350 ;
        RECT 1486.820 1745.230 1487.080 1745.550 ;
        RECT 1473.020 1738.430 1473.280 1738.750 ;
        RECT 1459.220 1738.090 1459.480 1738.410 ;
        RECT 1452.320 1731.630 1452.580 1731.950 ;
        RECT 1438.520 1722.450 1438.780 1722.770 ;
        RECT 1431.620 1717.350 1431.880 1717.670 ;
        RECT 1487.340 1648.650 1487.480 2789.030 ;
        RECT 1493.720 2053.610 1493.980 2053.930 ;
        RECT 1493.780 1918.270 1493.920 2053.610 ;
        RECT 1493.720 1917.950 1493.980 1918.270 ;
        RECT 1507.580 1718.010 1507.720 3187.850 ;
        RECT 1548.920 2946.450 1549.180 2946.770 ;
        RECT 1535.110 2898.315 1535.390 2898.685 ;
        RECT 1528.210 2891.515 1528.490 2891.885 ;
        RECT 1528.280 2804.650 1528.420 2891.515 ;
        RECT 1528.220 2804.330 1528.480 2804.650 ;
        RECT 1514.420 2789.370 1514.680 2789.690 ;
        RECT 1507.520 1717.690 1507.780 1718.010 ;
        RECT 1487.280 1648.330 1487.540 1648.650 ;
        RECT 1514.480 1642.190 1514.620 2789.370 ;
        RECT 1528.280 2059.710 1528.420 2804.330 ;
        RECT 1532.360 2066.870 1532.620 2067.190 ;
        RECT 1531.900 2065.850 1532.160 2066.170 ;
        RECT 1531.960 2065.150 1532.100 2065.850 ;
        RECT 1532.420 2065.490 1532.560 2066.870 ;
        RECT 1532.360 2065.170 1532.620 2065.490 ;
        RECT 1531.900 2064.830 1532.160 2065.150 ;
        RECT 1528.220 2059.390 1528.480 2059.710 ;
        RECT 1514.420 1641.870 1514.680 1642.190 ;
        RECT 1528.280 1614.650 1528.420 2059.390 ;
        RECT 1535.180 1669.730 1535.320 2898.315 ;
        RECT 1548.980 2801.250 1549.120 2946.450 ;
      LAYER met2 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met2 ;
        RECT 1932.160 3249.565 1932.300 3251.430 ;
        RECT 1932.090 3249.195 1932.370 3249.565 ;
        RECT 1939.060 2948.325 1939.200 3264.010 ;
        RECT 1938.990 2947.955 1939.270 2948.325 ;
        RECT 1945.890 2904.435 1946.170 2904.805 ;
        RECT 1945.960 2801.250 1946.100 2904.435 ;
        RECT 1548.920 2800.930 1549.180 2801.250 ;
        RECT 1552.140 2800.930 1552.400 2801.250 ;
        RECT 1945.900 2800.930 1946.160 2801.250 ;
        RECT 1552.200 1949.210 1552.340 2800.930 ;
        RECT 1645.510 2799.035 1645.790 2799.405 ;
        RECT 1688.750 2799.035 1689.030 2799.405 ;
        RECT 1788.570 2799.035 1788.850 2799.405 ;
        RECT 1607.790 2794.275 1608.070 2794.645 ;
        RECT 1614.690 2794.275 1614.970 2794.645 ;
        RECT 1621.590 2794.275 1621.870 2794.645 ;
        RECT 1628.490 2794.275 1628.770 2794.645 ;
        RECT 1635.390 2794.275 1635.670 2794.645 ;
        RECT 1587.090 2789.515 1587.370 2789.885 ;
        RECT 1600.890 2789.515 1601.170 2789.885 ;
        RECT 1587.100 2789.370 1587.360 2789.515 ;
        RECT 1600.960 2789.350 1601.100 2789.515 ;
        RECT 1600.900 2789.030 1601.160 2789.350 ;
        RECT 1580.190 2787.475 1580.470 2787.845 ;
        RECT 1593.990 2787.475 1594.270 2787.845 ;
        RECT 1601.350 2787.475 1601.630 2787.845 ;
        RECT 1579.280 2066.870 1579.540 2067.190 ;
        RECT 1579.340 2065.490 1579.480 2066.870 ;
        RECT 1579.740 2065.850 1580.000 2066.170 ;
        RECT 1579.280 2065.170 1579.540 2065.490 ;
        RECT 1579.800 2065.150 1579.940 2065.850 ;
        RECT 1579.740 2064.830 1580.000 2065.150 ;
        RECT 1555.820 2059.050 1556.080 2059.370 ;
        RECT 1555.880 2021.630 1556.020 2059.050 ;
        RECT 1555.820 2021.310 1556.080 2021.630 ;
        RECT 1552.140 1948.890 1552.400 1949.210 ;
        RECT 1580.260 1711.210 1580.400 2787.475 ;
        RECT 1591.240 2067.550 1591.500 2067.870 ;
        RECT 1590.780 2066.870 1591.040 2067.190 ;
        RECT 1590.320 2065.850 1590.580 2066.170 ;
        RECT 1580.200 1710.890 1580.460 1711.210 ;
        RECT 1535.120 1669.410 1535.380 1669.730 ;
        RECT 1590.380 1621.450 1590.520 2065.850 ;
        RECT 1590.840 1628.250 1590.980 2066.870 ;
        RECT 1591.300 1635.390 1591.440 2067.550 ;
        RECT 1594.060 1648.990 1594.200 2787.475 ;
        RECT 1601.420 1656.130 1601.560 2787.475 ;
        RECT 1607.860 1834.970 1608.000 2794.275 ;
        RECT 1611.010 2793.595 1611.290 2793.965 ;
        RECT 1611.080 2789.350 1611.220 2793.595 ;
        RECT 1611.020 2789.030 1611.280 2789.350 ;
        RECT 1607.800 1834.650 1608.060 1834.970 ;
        RECT 1611.080 1793.830 1611.220 2789.030 ;
        RECT 1614.760 1835.310 1614.900 2794.275 ;
        RECT 1617.910 2793.595 1618.190 2793.965 ;
        RECT 1617.980 2789.690 1618.120 2793.595 ;
        RECT 1617.920 2789.370 1618.180 2789.690 ;
        RECT 1614.700 1834.990 1614.960 1835.310 ;
        RECT 1617.980 1800.630 1618.120 2789.370 ;
        RECT 1621.660 1842.450 1621.800 2794.275 ;
        RECT 1624.810 2793.595 1625.090 2793.965 ;
        RECT 1624.880 2789.010 1625.020 2793.595 ;
        RECT 1624.820 2788.690 1625.080 2789.010 ;
        RECT 1621.600 1842.130 1621.860 1842.450 ;
        RECT 1624.880 1800.970 1625.020 2788.690 ;
        RECT 1628.560 1849.250 1628.700 2794.275 ;
        RECT 1631.710 2793.595 1631.990 2793.965 ;
        RECT 1631.780 2790.030 1631.920 2793.595 ;
        RECT 1631.720 2789.710 1631.980 2790.030 ;
        RECT 1629.420 2068.910 1629.680 2069.230 ;
        RECT 1628.960 2068.570 1629.220 2068.890 ;
        RECT 1629.020 2065.150 1629.160 2068.570 ;
        RECT 1629.480 2065.490 1629.620 2068.910 ;
        RECT 1629.420 2065.170 1629.680 2065.490 ;
        RECT 1628.960 2064.830 1629.220 2065.150 ;
        RECT 1628.500 1848.930 1628.760 1849.250 ;
        RECT 1631.780 1807.770 1631.920 2789.710 ;
        RECT 1635.460 1855.710 1635.600 2794.275 ;
        RECT 1642.300 2793.965 1642.560 2794.110 ;
        RECT 1638.610 2793.595 1638.890 2793.965 ;
        RECT 1642.290 2793.595 1642.570 2793.965 ;
        RECT 1638.680 2787.990 1638.820 2793.595 ;
        RECT 1642.760 2793.450 1643.020 2793.770 ;
        RECT 1642.820 2792.660 1642.960 2793.450 ;
        RECT 1642.360 2792.605 1642.960 2792.660 ;
        RECT 1642.290 2792.520 1642.960 2792.605 ;
        RECT 1642.290 2792.235 1642.570 2792.520 ;
        RECT 1638.620 2787.670 1638.880 2787.990 ;
        RECT 1635.400 1855.390 1635.660 1855.710 ;
        RECT 1638.680 1814.230 1638.820 2787.670 ;
        RECT 1642.290 2785.435 1642.570 2785.805 ;
        RECT 1642.360 1856.050 1642.500 2785.435 ;
        RECT 1642.300 1855.730 1642.560 1856.050 ;
        RECT 1645.580 1814.570 1645.720 2799.035 ;
        RECT 1646.430 2794.275 1646.710 2794.645 ;
        RECT 1649.190 2794.275 1649.470 2794.645 ;
        RECT 1652.410 2794.275 1652.690 2794.645 ;
        RECT 1656.090 2794.275 1656.370 2794.645 ;
        RECT 1662.990 2794.275 1663.270 2794.645 ;
        RECT 1669.890 2794.275 1670.170 2794.645 ;
        RECT 1676.790 2794.275 1677.070 2794.645 ;
        RECT 1646.500 2792.070 1646.640 2794.275 ;
        RECT 1646.440 2791.750 1646.700 2792.070 ;
        RECT 1646.500 1821.710 1646.640 2791.750 ;
        RECT 1649.260 1862.850 1649.400 2794.275 ;
        RECT 1649.650 2793.595 1649.930 2793.965 ;
        RECT 1649.720 1869.650 1649.860 2793.595 ;
        RECT 1652.480 2792.750 1652.620 2794.275 ;
        RECT 1652.420 2792.430 1652.680 2792.750 ;
        RECT 1649.660 1869.330 1649.920 1869.650 ;
        RECT 1649.200 1862.530 1649.460 1862.850 ;
        RECT 1652.480 1828.510 1652.620 2792.430 ;
        RECT 1656.160 1869.990 1656.300 2794.275 ;
        RECT 1658.850 2793.595 1659.130 2793.965 ;
        RECT 1658.920 2791.390 1659.060 2793.595 ;
        RECT 1656.560 2791.070 1656.820 2791.390 ;
        RECT 1658.860 2791.070 1659.120 2791.390 ;
        RECT 1656.620 2789.350 1656.760 2791.070 ;
        RECT 1656.560 2789.030 1656.820 2789.350 ;
        RECT 1663.060 1876.790 1663.200 2794.275 ;
        RECT 1663.450 2793.595 1663.730 2793.965 ;
        RECT 1663.520 2791.730 1663.660 2793.595 ;
        RECT 1663.460 2791.410 1663.720 2791.730 ;
        RECT 1663.520 2789.690 1663.660 2791.410 ;
        RECT 1663.460 2789.370 1663.720 2789.690 ;
        RECT 1669.960 1883.590 1670.100 2794.275 ;
        RECT 1670.350 2793.595 1670.630 2793.965 ;
        RECT 1670.420 2791.050 1670.560 2793.595 ;
        RECT 1670.360 2790.730 1670.620 2791.050 ;
        RECT 1670.420 2789.010 1670.560 2790.730 ;
        RECT 1670.360 2788.690 1670.620 2789.010 ;
        RECT 1675.880 2068.910 1676.140 2069.230 ;
        RECT 1675.940 2065.490 1676.080 2068.910 ;
        RECT 1676.340 2068.570 1676.600 2068.890 ;
        RECT 1675.880 2065.170 1676.140 2065.490 ;
        RECT 1676.400 2065.150 1676.540 2068.570 ;
        RECT 1676.340 2064.830 1676.600 2065.150 ;
        RECT 1676.860 1890.390 1677.000 2794.275 ;
        RECT 1677.260 2794.130 1677.520 2794.450 ;
        RECT 1683.690 2794.275 1683.970 2794.645 ;
        RECT 1677.320 2793.965 1677.460 2794.130 ;
        RECT 1677.250 2793.595 1677.530 2793.965 ;
        RECT 1682.310 2793.595 1682.590 2793.965 ;
        RECT 1677.320 2790.030 1677.460 2793.595 ;
        RECT 1682.380 2793.090 1682.520 2793.595 ;
        RECT 1682.320 2792.770 1682.580 2793.090 ;
        RECT 1677.260 2789.710 1677.520 2790.030 ;
        RECT 1682.380 2787.990 1682.520 2792.770 ;
        RECT 1682.320 2787.670 1682.580 2787.990 ;
        RECT 1683.760 1890.730 1683.900 2794.275 ;
        RECT 1688.820 2792.410 1688.960 2799.035 ;
        RECT 1740.730 2796.315 1741.010 2796.685 ;
        RECT 1740.270 2795.635 1740.550 2796.005 ;
        RECT 1690.590 2794.275 1690.870 2794.645 ;
        RECT 1697.490 2794.275 1697.770 2794.645 ;
        RECT 1706.230 2794.275 1706.510 2794.645 ;
        RECT 1712.670 2794.275 1712.950 2794.645 ;
        RECT 1718.190 2794.275 1718.470 2794.645 ;
        RECT 1724.170 2794.275 1724.450 2794.645 ;
        RECT 1728.770 2794.275 1729.050 2794.645 ;
        RECT 1734.290 2794.275 1734.570 2794.645 ;
        RECT 1690.140 2793.965 1690.400 2794.110 ;
        RECT 1689.680 2793.450 1689.940 2793.770 ;
        RECT 1690.130 2793.595 1690.410 2793.965 ;
        RECT 1689.740 2792.660 1689.880 2793.450 ;
        RECT 1689.740 2792.605 1690.340 2792.660 ;
        RECT 1689.740 2792.520 1690.410 2792.605 ;
        RECT 1688.760 2792.090 1689.020 2792.410 ;
        RECT 1690.130 2792.235 1690.410 2792.520 ;
        RECT 1684.150 2789.515 1684.430 2789.885 ;
        RECT 1684.220 1897.530 1684.360 2789.515 ;
        RECT 1690.130 1949.035 1690.410 1949.405 ;
        RECT 1690.140 1948.890 1690.400 1949.035 ;
        RECT 1686.910 1906.195 1687.190 1906.565 ;
        RECT 1684.160 1897.210 1684.420 1897.530 ;
        RECT 1683.700 1890.410 1683.960 1890.730 ;
        RECT 1676.800 1890.070 1677.060 1890.390 ;
        RECT 1669.900 1883.270 1670.160 1883.590 ;
        RECT 1663.000 1876.470 1663.260 1876.790 ;
        RECT 1656.100 1869.670 1656.360 1869.990 ;
        RECT 1652.420 1828.190 1652.680 1828.510 ;
        RECT 1646.440 1821.390 1646.700 1821.710 ;
        RECT 1645.520 1814.250 1645.780 1814.570 ;
        RECT 1638.620 1813.910 1638.880 1814.230 ;
        RECT 1631.720 1807.450 1631.980 1807.770 ;
        RECT 1624.820 1800.650 1625.080 1800.970 ;
        RECT 1617.920 1800.310 1618.180 1800.630 ;
        RECT 1611.020 1793.510 1611.280 1793.830 ;
        RECT 1601.360 1655.810 1601.620 1656.130 ;
        RECT 1594.000 1648.670 1594.260 1648.990 ;
        RECT 1591.240 1635.070 1591.500 1635.390 ;
        RECT 1590.780 1627.930 1591.040 1628.250 ;
        RECT 1590.320 1621.130 1590.580 1621.450 ;
        RECT 1528.220 1614.330 1528.480 1614.650 ;
        RECT 1421.500 1610.930 1421.760 1611.250 ;
        RECT 1427.940 1610.930 1428.200 1611.250 ;
        RECT 1421.560 1607.850 1421.700 1610.930 ;
        RECT 1414.140 1607.530 1414.400 1607.850 ;
        RECT 1421.500 1607.530 1421.760 1607.850 ;
        RECT 1414.200 1607.365 1414.340 1607.530 ;
        RECT 1414.130 1606.995 1414.410 1607.365 ;
        RECT 1686.980 1605.130 1687.120 1906.195 ;
        RECT 1690.660 1904.330 1690.800 2794.275 ;
        RECT 1695.190 2793.595 1695.470 2793.965 ;
        RECT 1695.260 2792.070 1695.400 2793.595 ;
        RECT 1695.200 2791.750 1695.460 2792.070 ;
        RECT 1697.560 1911.130 1697.700 2794.275 ;
        RECT 1699.330 2793.595 1699.610 2793.965 ;
        RECT 1699.400 2792.750 1699.540 2793.595 ;
        RECT 1699.340 2792.430 1699.600 2792.750 ;
        RECT 1706.300 2791.390 1706.440 2794.275 ;
        RECT 1712.740 2791.730 1712.880 2794.275 ;
        RECT 1712.680 2791.410 1712.940 2791.730 ;
        RECT 1706.240 2791.070 1706.500 2791.390 ;
        RECT 1718.260 2791.050 1718.400 2794.275 ;
        RECT 1724.180 2794.130 1724.440 2794.275 ;
        RECT 1724.240 2793.430 1724.380 2794.130 ;
        RECT 1724.180 2793.110 1724.440 2793.430 ;
        RECT 1728.840 2793.090 1728.980 2794.275 ;
        RECT 1728.780 2792.770 1729.040 2793.090 ;
        RECT 1728.310 2792.235 1728.590 2792.605 ;
        RECT 1734.360 2792.410 1734.500 2794.275 ;
        RECT 1740.340 2793.285 1740.480 2795.635 ;
        RECT 1740.270 2792.915 1740.550 2793.285 ;
        RECT 1718.200 2790.730 1718.460 2791.050 ;
        RECT 1728.380 2790.565 1728.520 2792.235 ;
        RECT 1734.300 2792.090 1734.560 2792.410 ;
        RECT 1740.800 2791.730 1740.940 2796.315 ;
        RECT 1741.190 2794.275 1741.470 2794.645 ;
        RECT 1747.630 2794.275 1747.910 2794.645 ;
        RECT 1758.670 2794.275 1758.950 2794.645 ;
        RECT 1741.260 2792.070 1741.400 2794.275 ;
        RECT 1747.700 2792.750 1747.840 2794.275 ;
        RECT 1747.640 2792.430 1747.900 2792.750 ;
        RECT 1752.690 2792.235 1752.970 2792.605 ;
        RECT 1741.200 2791.750 1741.460 2792.070 ;
        RECT 1740.740 2791.410 1741.000 2791.730 ;
        RECT 1752.760 2791.390 1752.900 2792.235 ;
        RECT 1752.700 2791.070 1752.960 2791.390 ;
        RECT 1758.740 2791.245 1758.880 2794.275 ;
        RECT 1766.490 2793.595 1766.770 2793.965 ;
        RECT 1773.390 2793.595 1773.670 2793.965 ;
        RECT 1780.290 2793.595 1780.570 2793.965 ;
        RECT 1766.560 2793.430 1766.700 2793.595 ;
        RECT 1766.500 2793.110 1766.760 2793.430 ;
        RECT 1773.460 2793.090 1773.600 2793.595 ;
        RECT 1773.400 2792.770 1773.660 2793.090 ;
        RECT 1780.360 2792.410 1780.500 2793.595 ;
        RECT 1788.640 2792.750 1788.780 2799.035 ;
        RECT 1780.300 2792.090 1780.560 2792.410 ;
        RECT 1787.190 2792.235 1787.470 2792.605 ;
        RECT 1788.580 2792.430 1788.840 2792.750 ;
        RECT 1787.260 2792.070 1787.400 2792.235 ;
        RECT 1787.200 2791.750 1787.460 2792.070 ;
        RECT 1758.670 2790.875 1758.950 2791.245 ;
        RECT 1759.590 2790.875 1759.870 2791.245 ;
        RECT 1773.390 2790.875 1773.670 2791.245 ;
        RECT 1759.600 2790.730 1759.860 2790.875 ;
        RECT 1773.460 2790.710 1773.600 2790.875 ;
        RECT 1728.310 2790.195 1728.590 2790.565 ;
        RECT 1759.590 2790.195 1759.870 2790.565 ;
        RECT 1773.400 2790.390 1773.660 2790.710 ;
        RECT 1759.660 2788.670 1759.800 2790.195 ;
        RECT 1766.490 2789.515 1766.770 2789.885 ;
        RECT 1718.650 2788.155 1718.930 2788.525 ;
        RECT 1759.600 2788.350 1759.860 2788.670 ;
        RECT 1766.560 2788.330 1766.700 2789.515 ;
        RECT 1704.390 2787.475 1704.670 2787.845 ;
        RECT 1711.290 2787.475 1711.570 2787.845 ;
        RECT 1718.190 2787.475 1718.470 2787.845 ;
        RECT 1704.460 2053.590 1704.600 2787.475 ;
        RECT 1711.360 2053.930 1711.500 2787.475 ;
        RECT 1718.260 2061.750 1718.400 2787.475 ;
        RECT 1718.720 2062.090 1718.860 2788.155 ;
        RECT 1766.500 2788.010 1766.760 2788.330 ;
        RECT 1725.090 2787.475 1725.370 2787.845 ;
        RECT 1731.990 2787.475 1732.270 2787.845 ;
        RECT 1738.890 2787.475 1739.170 2787.845 ;
        RECT 1745.790 2787.475 1746.070 2787.845 ;
        RECT 1753.150 2787.475 1753.430 2787.845 ;
        RECT 1718.660 2061.770 1718.920 2062.090 ;
        RECT 1718.200 2061.430 1718.460 2061.750 ;
        RECT 1725.160 2061.410 1725.300 2787.475 ;
        RECT 1726.020 2068.910 1726.280 2069.230 ;
        RECT 1725.560 2068.570 1725.820 2068.890 ;
        RECT 1725.620 2065.150 1725.760 2068.570 ;
        RECT 1726.080 2065.490 1726.220 2068.910 ;
        RECT 1726.020 2065.170 1726.280 2065.490 ;
        RECT 1725.560 2064.830 1725.820 2065.150 ;
        RECT 1725.100 2061.090 1725.360 2061.410 ;
        RECT 1732.060 2061.070 1732.200 2787.475 ;
        RECT 1732.000 2060.750 1732.260 2061.070 ;
        RECT 1738.960 2060.730 1739.100 2787.475 ;
        RECT 1738.900 2060.410 1739.160 2060.730 ;
        RECT 1745.860 2060.390 1746.000 2787.475 ;
        RECT 1745.800 2060.070 1746.060 2060.390 ;
        RECT 1753.220 2060.050 1753.360 2787.475 ;
        RECT 1835.500 2145.750 1835.760 2146.070 ;
        RECT 1835.560 2069.765 1835.700 2145.750 ;
        RECT 1842.400 2138.950 1842.660 2139.270 ;
        RECT 1842.460 2069.765 1842.600 2138.950 ;
        RECT 1849.300 2132.490 1849.560 2132.810 ;
        RECT 1849.360 2069.765 1849.500 2132.490 ;
        RECT 1856.200 2132.150 1856.460 2132.470 ;
        RECT 1856.260 2069.765 1856.400 2132.150 ;
        RECT 1863.100 2125.350 1863.360 2125.670 ;
        RECT 1863.160 2069.765 1863.300 2125.350 ;
        RECT 1870.000 2118.210 1870.260 2118.530 ;
        RECT 1870.060 2069.765 1870.200 2118.210 ;
        RECT 1870.460 2111.750 1870.720 2112.070 ;
        RECT 1835.490 2069.395 1835.770 2069.765 ;
        RECT 1842.390 2069.395 1842.670 2069.765 ;
        RECT 1849.290 2069.395 1849.570 2069.765 ;
        RECT 1856.190 2069.395 1856.470 2069.765 ;
        RECT 1863.090 2069.395 1863.370 2069.765 ;
        RECT 1869.990 2069.395 1870.270 2069.765 ;
        RECT 1772.480 2068.910 1772.740 2069.230 ;
        RECT 1870.520 2069.085 1870.660 2111.750 ;
        RECT 1876.900 2111.410 1877.160 2111.730 ;
        RECT 1876.960 2069.765 1877.100 2111.410 ;
        RECT 1883.800 2104.610 1884.060 2104.930 ;
        RECT 1883.860 2069.765 1884.000 2104.610 ;
        RECT 1890.700 2097.470 1890.960 2097.790 ;
        RECT 1890.760 2069.765 1890.900 2097.470 ;
        RECT 1897.600 2091.010 1897.860 2091.330 ;
        RECT 1897.660 2069.765 1897.800 2091.010 ;
        RECT 1904.500 2090.670 1904.760 2090.990 ;
        RECT 1904.560 2069.765 1904.700 2090.670 ;
        RECT 1911.400 2083.870 1911.660 2084.190 ;
        RECT 1911.460 2069.765 1911.600 2083.870 ;
        RECT 1911.860 2077.070 1912.120 2077.390 ;
        RECT 1876.890 2069.395 1877.170 2069.765 ;
        RECT 1883.790 2069.395 1884.070 2069.765 ;
        RECT 1890.690 2069.395 1890.970 2069.765 ;
        RECT 1897.590 2069.395 1897.870 2069.765 ;
        RECT 1904.490 2069.395 1904.770 2069.765 ;
        RECT 1911.390 2069.395 1911.670 2069.765 ;
        RECT 1772.540 2065.490 1772.680 2068.910 ;
        RECT 1772.940 2068.570 1773.200 2068.890 ;
        RECT 1848.840 2068.570 1849.100 2068.890 ;
        RECT 1870.450 2068.715 1870.730 2069.085 ;
        RECT 1890.240 2068.910 1890.500 2069.230 ;
        RECT 1911.920 2069.085 1912.060 2077.070 ;
        RECT 1919.220 2070.270 1919.480 2070.590 ;
        RECT 1917.840 2069.250 1918.100 2069.570 ;
        RECT 1772.480 2065.170 1772.740 2065.490 ;
        RECT 1773.000 2065.150 1773.140 2068.570 ;
        RECT 1841.480 2068.230 1841.740 2068.550 ;
        RECT 1841.540 2067.045 1841.680 2068.230 ;
        RECT 1843.780 2067.890 1844.040 2068.210 ;
        RECT 1844.240 2067.890 1844.500 2068.210 ;
        RECT 1843.840 2067.045 1843.980 2067.890 ;
        RECT 1844.300 2067.530 1844.440 2067.890 ;
        RECT 1844.240 2067.210 1844.500 2067.530 ;
        RECT 1844.700 2067.210 1844.960 2067.530 ;
        RECT 1841.470 2066.675 1841.750 2067.045 ;
        RECT 1843.770 2066.675 1844.050 2067.045 ;
        RECT 1844.760 2065.830 1844.900 2067.210 ;
        RECT 1848.900 2067.045 1849.040 2068.570 ;
        RECT 1890.300 2068.550 1890.440 2068.910 ;
        RECT 1893.920 2068.570 1894.180 2068.890 ;
        RECT 1911.850 2068.715 1912.130 2069.085 ;
        RECT 1890.240 2068.230 1890.500 2068.550 ;
        RECT 1849.300 2067.890 1849.560 2068.210 ;
        RECT 1848.830 2066.675 1849.110 2067.045 ;
        RECT 1849.360 2066.365 1849.500 2067.890 ;
        RECT 1864.940 2067.210 1865.200 2067.530 ;
        RECT 1859.880 2066.530 1860.140 2066.850 ;
        RECT 1849.290 2065.995 1849.570 2066.365 ;
        RECT 1844.700 2065.510 1844.960 2065.830 ;
        RECT 1859.940 2065.685 1860.080 2066.530 ;
        RECT 1865.000 2065.685 1865.140 2067.210 ;
        RECT 1890.300 2067.045 1890.440 2068.230 ;
        RECT 1890.230 2066.675 1890.510 2067.045 ;
        RECT 1893.980 2065.685 1894.120 2068.570 ;
        RECT 1898.060 2067.890 1898.320 2068.210 ;
        RECT 1898.120 2066.365 1898.260 2067.890 ;
        RECT 1911.400 2067.210 1911.660 2067.530 ;
        RECT 1907.720 2066.530 1907.980 2066.850 ;
        RECT 1898.050 2065.995 1898.330 2066.365 ;
        RECT 1907.780 2065.685 1907.920 2066.530 ;
        RECT 1911.460 2065.830 1911.600 2067.210 ;
        RECT 1911.400 2065.685 1911.660 2065.830 ;
        RECT 1844.240 2065.170 1844.500 2065.490 ;
        RECT 1859.870 2065.315 1860.150 2065.685 ;
        RECT 1864.930 2065.315 1865.210 2065.685 ;
        RECT 1877.360 2065.170 1877.620 2065.490 ;
        RECT 1893.910 2065.315 1894.190 2065.685 ;
        RECT 1907.710 2065.315 1907.990 2065.685 ;
        RECT 1911.390 2065.315 1911.670 2065.685 ;
        RECT 1772.940 2064.830 1773.200 2065.150 ;
        RECT 1844.300 2064.890 1844.440 2065.170 ;
        RECT 1846.540 2064.890 1846.800 2065.150 ;
        RECT 1871.840 2065.005 1872.100 2065.150 ;
        RECT 1844.300 2064.830 1846.800 2064.890 ;
        RECT 1844.300 2064.750 1846.740 2064.830 ;
        RECT 1871.830 2064.635 1872.110 2065.005 ;
        RECT 1877.420 2064.325 1877.560 2065.170 ;
        RECT 1917.380 2064.890 1917.640 2065.150 ;
        RECT 1917.900 2065.005 1918.040 2069.250 ;
        RECT 1919.280 2069.085 1919.420 2070.270 ;
        RECT 1925.200 2069.930 1925.460 2070.250 ;
        RECT 1925.260 2069.765 1925.400 2069.930 ;
        RECT 1925.190 2069.395 1925.470 2069.765 ;
        RECT 1965.680 2069.250 1965.940 2069.570 ;
        RECT 1919.210 2068.715 1919.490 2069.085 ;
        RECT 1936.700 2068.910 1936.960 2069.230 ;
        RECT 1930.260 2068.230 1930.520 2068.550 ;
        RECT 1924.740 2067.210 1925.000 2067.530 ;
        RECT 1924.800 2065.150 1924.940 2067.210 ;
        RECT 1924.740 2065.005 1925.000 2065.150 ;
        RECT 1930.320 2065.005 1930.460 2068.230 ;
        RECT 1932.100 2066.365 1932.360 2066.510 ;
        RECT 1932.090 2065.995 1932.370 2066.365 ;
        RECT 1936.760 2065.685 1936.900 2068.910 ;
        RECT 1941.760 2068.570 1942.020 2068.890 ;
        RECT 1941.820 2067.045 1941.960 2068.570 ;
        RECT 1948.200 2067.890 1948.460 2068.210 ;
        RECT 1941.750 2066.675 1942.030 2067.045 ;
        RECT 1936.690 2065.315 1936.970 2065.685 ;
        RECT 1917.830 2064.890 1918.110 2065.005 ;
        RECT 1917.380 2064.830 1918.110 2064.890 ;
        RECT 1882.880 2064.490 1883.140 2064.810 ;
        RECT 1917.440 2064.750 1918.110 2064.830 ;
        RECT 1917.830 2064.635 1918.110 2064.750 ;
        RECT 1924.730 2064.635 1925.010 2065.005 ;
        RECT 1930.250 2064.635 1930.530 2065.005 ;
        RECT 1948.260 2064.810 1948.400 2067.890 ;
        RECT 1965.740 2066.850 1965.880 2069.250 ;
        RECT 1980.400 2068.910 1980.660 2069.230 ;
        RECT 1973.500 2068.230 1973.760 2068.550 ;
        RECT 1980.460 2068.405 1980.600 2068.910 ;
        RECT 1987.300 2068.570 1987.560 2068.890 ;
        RECT 1987.360 2068.405 1987.500 2068.570 ;
        RECT 1973.560 2067.530 1973.700 2068.230 ;
        RECT 1980.390 2068.035 1980.670 2068.405 ;
        RECT 1987.290 2068.035 1987.570 2068.405 ;
        RECT 2028.700 2067.725 2028.960 2067.870 ;
        RECT 1969.820 2067.210 1970.080 2067.530 ;
        RECT 1973.500 2067.210 1973.760 2067.530 ;
        RECT 1976.720 2067.210 1976.980 2067.530 ;
        RECT 2021.800 2067.210 2022.060 2067.530 ;
        RECT 2028.690 2067.355 2028.970 2067.725 ;
        RECT 1954.640 2066.530 1954.900 2066.850 ;
        RECT 1959.240 2066.530 1959.500 2066.850 ;
        RECT 1965.680 2066.530 1965.940 2066.850 ;
        RECT 1930.260 2064.490 1930.520 2064.635 ;
        RECT 1948.200 2064.490 1948.460 2064.810 ;
        RECT 1882.940 2064.325 1883.080 2064.490 ;
        RECT 1930.320 2064.335 1930.460 2064.490 ;
        RECT 1877.350 2063.955 1877.630 2064.325 ;
        RECT 1882.870 2063.955 1883.150 2064.325 ;
        RECT 1948.260 2063.645 1948.400 2064.490 ;
        RECT 1954.700 2063.645 1954.840 2066.530 ;
        RECT 1959.300 2065.830 1959.440 2066.530 ;
        RECT 1958.780 2065.510 1959.040 2065.830 ;
        RECT 1959.240 2065.510 1959.500 2065.830 ;
        RECT 1958.840 2063.645 1958.980 2065.510 ;
        RECT 1965.740 2063.645 1965.880 2066.530 ;
        RECT 1969.880 2066.510 1970.020 2067.210 ;
        RECT 1969.820 2066.190 1970.080 2066.510 ;
        RECT 1966.600 2064.325 1966.860 2064.470 ;
        RECT 1966.590 2063.955 1966.870 2064.325 ;
        RECT 1969.880 2063.645 1970.020 2066.190 ;
        RECT 1973.500 2063.810 1973.760 2064.130 ;
        RECT 1973.560 2063.645 1973.700 2063.810 ;
        RECT 1976.780 2063.645 1976.920 2067.210 ;
        RECT 2021.860 2067.045 2022.000 2067.210 ;
        RECT 2008.000 2066.530 2008.260 2066.850 ;
        RECT 2021.790 2066.675 2022.070 2067.045 ;
        RECT 2035.600 2066.870 2035.860 2067.190 ;
        RECT 2008.060 2066.365 2008.200 2066.530 ;
        RECT 2015.820 2066.365 2016.080 2066.510 ;
        RECT 2035.660 2066.365 2035.800 2066.870 ;
        RECT 2007.990 2065.995 2008.270 2066.365 ;
        RECT 2015.810 2065.995 2016.090 2066.365 ;
        RECT 2035.590 2065.995 2035.870 2066.365 ;
        RECT 2042.500 2065.850 2042.760 2066.170 ;
        RECT 1994.200 2065.685 1994.460 2065.830 ;
        RECT 2042.560 2065.685 2042.700 2065.850 ;
        RECT 1994.190 2065.315 1994.470 2065.685 ;
        RECT 2001.100 2065.170 2001.360 2065.490 ;
        RECT 2042.490 2065.315 2042.770 2065.685 ;
        RECT 2001.160 2065.005 2001.300 2065.170 ;
        RECT 1987.300 2064.490 1987.560 2064.810 ;
        RECT 2001.090 2064.635 2001.370 2065.005 ;
        RECT 1987.360 2064.325 1987.500 2064.490 ;
        RECT 1987.290 2063.955 1987.570 2064.325 ;
        RECT 1980.400 2063.645 1980.660 2063.790 ;
        RECT 1948.190 2063.275 1948.470 2063.645 ;
        RECT 1954.630 2063.275 1954.910 2063.645 ;
        RECT 1958.770 2063.275 1959.050 2063.645 ;
        RECT 1965.670 2063.275 1965.950 2063.645 ;
        RECT 1969.810 2063.275 1970.090 2063.645 ;
        RECT 1973.490 2063.275 1973.770 2063.645 ;
        RECT 1976.710 2063.275 1976.990 2063.645 ;
        RECT 1980.390 2063.275 1980.670 2063.645 ;
        RECT 2028.690 2063.275 2028.970 2063.645 ;
        RECT 2028.700 2063.130 2028.960 2063.275 ;
        RECT 1753.160 2059.730 1753.420 2060.050 ;
        RECT 2097.700 2059.390 2097.960 2059.710 ;
        RECT 1987.300 2059.050 1987.560 2059.370 ;
        RECT 1940.380 2058.885 1940.640 2059.030 ;
        RECT 1940.370 2058.515 1940.650 2058.885 ;
        RECT 1955.100 2058.370 1955.360 2058.690 ;
        RECT 1955.160 2058.205 1955.300 2058.370 ;
        RECT 1987.360 2058.205 1987.500 2059.050 ;
        RECT 1995.580 2058.205 1995.840 2058.350 ;
        RECT 1955.090 2057.835 1955.370 2058.205 ;
        RECT 1987.290 2057.835 1987.570 2058.205 ;
        RECT 1990.060 2057.690 1990.320 2058.010 ;
        RECT 1995.570 2057.835 1995.850 2058.205 ;
        RECT 1990.120 2057.525 1990.260 2057.690 ;
        RECT 2004.780 2057.525 2005.040 2057.670 ;
        RECT 1946.350 2057.155 1946.630 2057.525 ;
        RECT 1990.050 2057.155 1990.330 2057.525 ;
        RECT 2004.770 2057.155 2005.050 2057.525 ;
        RECT 1946.420 2056.310 1946.560 2057.155 ;
        RECT 2008.460 2057.010 2008.720 2057.330 ;
        RECT 2016.270 2057.155 2016.550 2057.525 ;
        RECT 2008.520 2056.845 2008.660 2057.010 ;
        RECT 2008.450 2056.475 2008.730 2056.845 ;
        RECT 2016.340 2056.650 2016.480 2057.155 ;
        RECT 2021.800 2056.845 2022.060 2056.990 ;
        RECT 2016.280 2056.330 2016.540 2056.650 ;
        RECT 2021.790 2056.475 2022.070 2056.845 ;
        RECT 1946.360 2055.990 1946.620 2056.310 ;
        RECT 1948.660 2055.650 1948.920 2055.970 ;
        RECT 1948.720 2055.485 1948.860 2055.650 ;
        RECT 1948.650 2055.115 1948.930 2055.485 ;
        RECT 1711.300 2053.610 1711.560 2053.930 ;
        RECT 1704.400 2053.270 1704.660 2053.590 ;
        RECT 1961.540 2052.930 1961.800 2053.250 ;
        RECT 1961.600 2052.085 1961.740 2052.930 ;
        RECT 2049.860 2052.590 2050.120 2052.910 ;
        RECT 2049.920 2052.085 2050.060 2052.590 ;
        RECT 1961.530 2051.715 1961.810 2052.085 ;
        RECT 2049.850 2051.715 2050.130 2052.085 ;
        RECT 1697.500 1910.810 1697.760 1911.130 ;
        RECT 1690.600 1904.010 1690.860 1904.330 ;
        RECT 1688.760 1610.930 1689.020 1611.250 ;
        RECT 1688.820 1610.085 1688.960 1610.930 ;
        RECT 1688.750 1609.715 1689.030 1610.085 ;
        RECT 1414.140 1604.810 1414.400 1605.130 ;
        RECT 1686.920 1604.810 1687.180 1605.130 ;
        RECT 1690.140 1604.810 1690.400 1605.130 ;
      LAYER met2 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met2 ;
        RECT 2097.760 1965.045 2097.900 2059.390 ;
        RECT 2097.690 1964.675 2097.970 1965.045 ;
        RECT 2097.690 1953.115 2097.970 1953.485 ;
        RECT 2082.050 1619.915 2082.330 1620.285 ;
        RECT 1414.200 1603.965 1414.340 1604.810 ;
        RECT 1414.130 1603.595 1414.410 1603.965 ;
        RECT 1413.680 1601.410 1413.940 1601.730 ;
        RECT 1410.460 1601.070 1410.720 1601.390 ;
        RECT 1690.200 1593.910 1690.340 1604.810 ;
        RECT 2082.120 1602.410 2082.260 1619.915 ;
        RECT 2097.760 1604.790 2097.900 1953.115 ;
        RECT 2099.530 1662.755 2099.810 1663.125 ;
        RECT 2099.070 1643.035 2099.350 1643.405 ;
        RECT 2098.610 1635.555 2098.890 1635.925 ;
        RECT 2098.150 1628.755 2098.430 1629.125 ;
        RECT 2097.700 1604.470 2097.960 1604.790 ;
        RECT 2098.220 1602.750 2098.360 1628.755 ;
        RECT 2098.680 1603.090 2098.820 1635.555 ;
        RECT 2099.140 1604.450 2099.280 1643.035 ;
        RECT 2099.080 1604.130 2099.340 1604.450 ;
        RECT 2098.620 1602.770 2098.880 1603.090 ;
        RECT 2098.160 1602.430 2098.420 1602.750 ;
        RECT 2082.060 1602.090 2082.320 1602.410 ;
        RECT 2099.600 1601.730 2099.740 1662.755 ;
        RECT 2100.910 1655.955 2101.190 1656.325 ;
        RECT 2099.990 1649.155 2100.270 1649.525 ;
        RECT 2099.540 1601.410 2099.800 1601.730 ;
        RECT 2100.060 1601.390 2100.200 1649.155 ;
        RECT 2100.980 1602.070 2101.120 1655.955 ;
        RECT 2100.920 1601.750 2101.180 1602.070 ;
        RECT 2100.000 1601.070 2100.260 1601.390 ;
        RECT 1720.100 1593.910 1720.240 1594.065 ;
        RECT 1690.140 1593.590 1690.400 1593.910 ;
        RECT 1720.040 1593.765 1720.300 1593.910 ;
        RECT 1720.030 1593.395 1720.310 1593.765 ;
        RECT 1720.100 1590.510 1720.240 1593.395 ;
        RECT 1738.890 1592.035 1739.170 1592.405 ;
        RECT 1738.960 1590.510 1739.100 1592.035 ;
        RECT 1720.040 1590.190 1720.300 1590.510 ;
        RECT 1738.900 1590.190 1739.160 1590.510 ;
      LAYER via2 ;
        RECT 646.390 3264.200 646.670 3264.480 ;
        RECT 668.470 3264.200 668.750 3264.480 ;
        RECT 1293.150 3264.200 1293.430 3264.480 ;
        RECT 288.050 3230.200 288.330 3230.480 ;
        RECT 287.590 3224.760 287.870 3225.040 ;
        RECT 287.130 3215.920 287.410 3216.200 ;
        RECT 286.670 3209.800 286.950 3210.080 ;
        RECT 286.210 3201.640 286.490 3201.920 ;
        RECT 285.290 3196.200 285.570 3196.480 ;
        RECT 284.830 2898.360 285.110 2898.640 ;
        RECT 284.370 2891.560 284.650 2891.840 ;
        RECT 285.750 3188.040 286.030 3188.320 ;
        RECT 688.250 3248.275 688.530 3248.555 ;
        RECT 1890.690 3264.200 1890.970 3264.480 ;
        RECT 1917.370 3264.200 1917.650 3264.480 ;
        RECT 1317.530 3258.080 1317.810 3258.360 ;
        RECT 1186.890 3252.640 1187.170 3252.920 ;
        RECT 1187.810 3252.640 1188.090 3252.920 ;
        RECT 941.710 3230.200 941.990 3230.480 ;
        RECT 941.250 3188.040 941.530 3188.320 ;
        RECT 696.990 2948.000 697.270 2948.280 ;
        RECT 337.730 2794.320 338.010 2794.600 ;
        RECT 344.630 2794.320 344.910 2794.600 ;
        RECT 351.530 2794.320 351.810 2794.600 ;
        RECT 358.430 2794.320 358.710 2794.600 ;
        RECT 363.030 2794.320 363.310 2794.600 ;
        RECT 365.330 2794.320 365.610 2794.600 ;
        RECT 369.010 2794.320 369.290 2794.600 ;
        RECT 371.310 2794.320 371.590 2794.600 ;
        RECT 374.990 2794.320 375.270 2794.600 ;
        RECT 380.050 2794.320 380.330 2794.600 ;
        RECT 384.190 2794.320 384.470 2794.600 ;
        RECT 386.950 2794.320 387.230 2794.600 ;
        RECT 392.470 2794.320 392.750 2794.600 ;
        RECT 397.070 2794.320 397.350 2794.600 ;
        RECT 399.830 2794.320 400.110 2794.600 ;
        RECT 403.970 2794.320 404.250 2794.600 ;
        RECT 406.270 2794.320 406.550 2794.600 ;
        RECT 409.490 2794.320 409.770 2794.600 ;
        RECT 413.630 2794.320 413.910 2794.600 ;
        RECT 419.150 2794.320 419.430 2794.600 ;
        RECT 420.990 2794.320 421.270 2794.600 ;
        RECT 427.430 2794.320 427.710 2794.600 ;
        RECT 432.030 2794.320 432.310 2794.600 ;
        RECT 434.330 2794.320 434.610 2794.600 ;
        RECT 439.390 2794.320 439.670 2794.600 ;
        RECT 441.230 2794.320 441.510 2794.600 ;
        RECT 444.450 2794.320 444.730 2794.600 ;
        RECT 448.130 2794.320 448.410 2794.600 ;
        RECT 449.050 2794.320 449.330 2794.600 ;
        RECT 455.030 2794.320 455.310 2794.600 ;
        RECT 462.390 2794.320 462.670 2794.600 ;
        RECT 468.370 2794.320 468.650 2794.600 ;
        RECT 474.350 2794.320 474.630 2794.600 ;
        RECT 475.730 2794.320 476.010 2794.600 ;
        RECT 478.950 2794.320 479.230 2794.600 ;
        RECT 482.630 2794.320 482.910 2794.600 ;
        RECT 484.930 2794.320 485.210 2794.600 ;
        RECT 489.070 2794.320 489.350 2794.600 ;
        RECT 490.450 2794.320 490.730 2794.600 ;
        RECT 496.430 2794.320 496.710 2794.600 ;
        RECT 497.810 2794.320 498.090 2794.600 ;
        RECT 501.950 2794.320 502.230 2794.600 ;
        RECT 510.230 2794.320 510.510 2794.600 ;
        RECT 517.130 2794.320 517.410 2794.600 ;
        RECT 524.030 2794.320 524.310 2794.600 ;
        RECT 527.710 2794.320 527.990 2794.600 ;
        RECT 530.930 2794.320 531.210 2794.600 ;
        RECT 537.370 2794.320 537.650 2794.600 ;
        RECT 542.430 2794.320 542.710 2794.600 ;
        RECT 551.630 2794.320 551.910 2794.600 ;
        RECT 351.070 2792.960 351.350 2793.240 ;
        RECT 379.130 2790.920 379.410 2791.200 ;
        RECT 392.930 2791.600 393.210 2791.880 ;
        RECT 397.990 2792.960 398.270 2793.240 ;
        RECT 414.090 2792.960 414.370 2793.240 ;
        RECT 426.050 2792.960 426.330 2793.240 ;
        RECT 419.150 2721.560 419.430 2721.840 ;
        RECT 433.870 2792.960 434.150 2793.240 ;
        RECT 429.270 2722.240 429.550 2722.520 ;
        RECT 439.850 2722.920 440.130 2723.200 ;
        RECT 455.490 2792.960 455.770 2793.240 ;
        RECT 461.930 2791.600 462.210 2791.880 ;
        RECT 466.530 2792.960 466.810 2793.240 ;
        RECT 460.550 2723.600 460.830 2723.880 ;
        RECT 468.830 2792.960 469.110 2793.240 ;
        RECT 489.990 2791.600 490.270 2791.880 ;
        RECT 500.110 2792.960 500.390 2793.240 ;
        RECT 509.770 2792.960 510.050 2793.240 ;
        RECT 507.010 2791.600 507.290 2791.880 ;
        RECT 513.910 2792.960 514.190 2793.240 ;
        RECT 519.430 2792.960 519.710 2793.240 ;
        RECT 534.610 2792.960 534.890 2793.240 ;
        RECT 530.930 2714.760 531.210 2715.040 ;
        RECT 538.750 2792.960 539.030 2793.240 ;
        RECT 541.510 2792.960 541.790 2793.240 ;
        RECT 707.570 2716.120 707.850 2716.400 ;
        RECT 720.910 2715.440 721.190 2715.720 ;
        RECT 942.170 3224.760 942.450 3225.040 ;
        RECT 942.630 3215.920 942.910 3216.200 ;
        RECT 943.090 3209.800 943.370 3210.080 ;
        RECT 942.630 2723.600 942.910 2723.880 ;
        RECT 943.550 3201.640 943.830 3201.920 ;
        RECT 944.470 3196.200 944.750 3196.480 ;
        RECT 944.010 2898.360 944.290 2898.640 ;
        RECT 943.550 2722.920 943.830 2723.200 ;
        RECT 944.930 2891.560 945.210 2891.840 ;
        RECT 1352.490 3249.920 1352.770 3250.200 ;
        RECT 1400.330 3249.920 1400.610 3250.200 ;
        RECT 1332.250 3249.240 1332.530 3249.520 ;
        RECT 1345.590 2946.640 1345.870 2946.920 ;
        RECT 1352.030 2946.640 1352.310 2946.920 ;
        RECT 1345.590 2938.480 1345.870 2938.760 ;
        RECT 1054.870 2799.760 1055.150 2800.040 ;
        RECT 979.890 2794.320 980.170 2794.600 ;
        RECT 986.790 2794.320 987.070 2794.600 ;
        RECT 1007.490 2794.320 1007.770 2794.600 ;
        RECT 1013.930 2794.320 1014.210 2794.600 ;
        RECT 1020.830 2794.320 1021.110 2794.600 ;
        RECT 1027.730 2794.320 1028.010 2794.600 ;
        RECT 1030.490 2794.320 1030.770 2794.600 ;
        RECT 1041.990 2794.320 1042.270 2794.600 ;
        RECT 1053.030 2794.320 1053.310 2794.600 ;
        RECT 944.470 2722.240 944.750 2722.520 ;
        RECT 941.250 2721.560 941.530 2721.840 ;
        RECT 1010.710 2792.960 1010.990 2793.240 ;
        RECT 1001.050 2788.880 1001.330 2789.160 ;
        RECT 993.690 2788.200 993.970 2788.480 ;
        RECT 1017.610 2793.640 1017.890 2793.920 ;
        RECT 1024.510 2792.960 1024.790 2793.240 ;
        RECT 1045.210 2792.960 1045.490 2793.240 ;
        RECT 1038.310 2788.200 1038.590 2788.480 ;
        RECT 1034.630 2787.520 1034.910 2787.800 ;
        RECT 1041.530 2787.520 1041.810 2787.800 ;
        RECT 1048.430 2787.520 1048.710 2787.800 ;
        RECT 1041.530 2716.120 1041.810 2716.400 ;
        RECT 1100.410 2795.000 1100.690 2795.280 ;
        RECT 1059.010 2794.320 1059.290 2794.600 ;
        RECT 1065.450 2794.320 1065.730 2794.600 ;
        RECT 1069.590 2794.320 1069.870 2794.600 ;
        RECT 1076.490 2794.320 1076.770 2794.600 ;
        RECT 1089.830 2794.320 1090.110 2794.600 ;
        RECT 1094.890 2794.320 1095.170 2794.600 ;
        RECT 1075.570 2791.600 1075.850 2791.880 ;
        RECT 1088.910 2793.640 1089.190 2793.920 ;
        RECT 1055.330 2788.200 1055.610 2788.480 ;
        RECT 1111.910 2794.320 1112.190 2794.600 ;
        RECT 1117.890 2794.320 1118.170 2794.600 ;
        RECT 1122.490 2794.320 1122.770 2794.600 ;
        RECT 1129.390 2794.320 1129.670 2794.600 ;
        RECT 1135.830 2794.320 1136.110 2794.600 ;
        RECT 1140.890 2794.320 1141.170 2794.600 ;
        RECT 1147.790 2794.320 1148.070 2794.600 ;
        RECT 1107.770 2791.600 1108.050 2791.880 ;
        RECT 1159.290 2793.640 1159.570 2793.920 ;
        RECT 1166.190 2793.640 1166.470 2793.920 ;
        RECT 1174.470 2792.960 1174.750 2793.240 ;
        RECT 1186.890 2792.960 1187.170 2793.240 ;
        RECT 1159.750 2792.280 1160.030 2792.560 ;
        RECT 1152.390 2791.600 1152.670 2791.880 ;
        RECT 1159.290 2791.600 1159.570 2791.880 ;
        RECT 1193.790 2792.280 1194.070 2792.560 ;
        RECT 1089.370 2788.200 1089.650 2788.480 ;
        RECT 1130.770 2788.200 1131.050 2788.480 ;
        RECT 1165.730 2788.200 1166.010 2788.480 ;
        RECT 1062.230 2787.520 1062.510 2787.800 ;
        RECT 1069.130 2787.520 1069.410 2787.800 ;
        RECT 1076.030 2787.520 1076.310 2787.800 ;
        RECT 1082.930 2787.520 1083.210 2787.800 ;
        RECT 1030.950 2714.760 1031.230 2715.040 ;
        RECT 1052.110 2715.440 1052.390 2715.720 ;
        RECT 1089.830 2787.520 1090.110 2787.800 ;
        RECT 1096.730 2787.520 1097.010 2787.800 ;
        RECT 1103.630 2787.520 1103.910 2787.800 ;
        RECT 1110.530 2787.520 1110.810 2787.800 ;
        RECT 1117.430 2787.520 1117.710 2787.800 ;
        RECT 1124.330 2787.520 1124.610 2787.800 ;
        RECT 1131.230 2787.520 1131.510 2787.800 ;
        RECT 1138.130 2787.520 1138.410 2787.800 ;
        RECT 1145.030 2787.520 1145.310 2787.800 ;
        RECT 1151.930 2787.520 1152.210 2787.800 ;
        RECT 1158.830 2787.520 1159.110 2787.800 ;
        RECT 1165.270 2787.520 1165.550 2787.800 ;
        RECT 1172.630 2787.520 1172.910 2787.800 ;
        RECT 1179.530 2787.520 1179.810 2787.800 ;
        RECT 1186.430 2787.520 1186.710 2787.800 ;
        RECT 1193.330 2787.520 1193.610 2787.800 ;
        RECT 1200.230 2787.520 1200.510 2787.800 ;
        RECT 1407.690 2146.960 1407.970 2147.240 ;
        RECT 1407.690 2142.200 1407.970 2142.480 ;
        RECT 1408.150 2136.760 1408.430 2137.040 ;
        RECT 1407.690 2132.000 1407.970 2132.280 ;
        RECT 1407.690 2126.560 1407.970 2126.840 ;
        RECT 1407.690 2121.800 1407.970 2122.080 ;
        RECT 1408.150 2117.040 1408.430 2117.320 ;
        RECT 1407.690 2111.600 1407.970 2111.880 ;
        RECT 1407.690 2106.840 1407.970 2107.120 ;
        RECT 1407.690 2101.400 1407.970 2101.680 ;
        RECT 1408.150 2096.640 1408.430 2096.920 ;
        RECT 1407.690 2091.200 1407.970 2091.480 ;
        RECT 1414.130 2086.440 1414.410 2086.720 ;
        RECT 1411.370 2081.680 1411.650 2081.960 ;
        RECT 1408.610 2076.240 1408.890 2076.520 ;
        RECT 1410.450 2071.480 1410.730 2071.760 ;
        RECT 1409.530 2051.080 1409.810 2051.360 ;
        RECT 1410.450 2061.280 1410.730 2061.560 ;
        RECT 1409.070 2030.680 1409.350 2030.960 ;
        RECT 1408.610 2025.920 1408.890 2026.200 ;
        RECT 1409.530 2015.720 1409.810 2016.000 ;
        RECT 1408.150 2005.520 1408.430 2005.800 ;
        RECT 1408.150 2000.760 1408.430 2001.040 ;
        RECT 1408.150 1995.320 1408.430 1995.600 ;
        RECT 1408.150 1970.160 1408.430 1970.440 ;
        RECT 1408.610 1966.080 1408.890 1966.360 ;
        RECT 1408.150 1965.400 1408.430 1965.680 ;
        RECT 1408.150 1959.960 1408.430 1960.240 ;
        RECT 1408.150 1940.240 1408.430 1940.520 ;
        RECT 1408.150 1934.800 1408.430 1935.080 ;
        RECT 1408.610 1930.040 1408.890 1930.320 ;
        RECT 1408.150 1925.280 1408.430 1925.560 ;
        RECT 1408.150 1919.840 1408.430 1920.120 ;
        RECT 1409.530 1950.440 1409.810 1950.720 ;
        RECT 1408.150 1909.640 1408.430 1909.920 ;
        RECT 1408.610 1904.880 1408.890 1905.160 ;
        RECT 1408.610 1803.560 1408.890 1803.840 ;
        RECT 1409.530 1788.600 1409.810 1788.880 ;
        RECT 1409.990 1783.840 1410.270 1784.120 ;
        RECT 1412.290 2039.520 1412.570 2039.800 ;
        RECT 1410.910 2010.960 1411.190 2011.240 ;
        RECT 1410.910 1990.560 1411.190 1990.840 ;
        RECT 1410.910 1884.480 1411.190 1884.760 ;
        RECT 1410.910 1864.080 1411.190 1864.360 ;
        RECT 1410.910 1849.120 1411.190 1849.400 ;
        RECT 1410.910 1828.720 1411.190 1829.000 ;
        RECT 1410.450 1778.400 1410.730 1778.680 ;
        RECT 1410.910 1773.640 1411.190 1773.920 ;
        RECT 1409.990 1772.960 1410.270 1773.240 ;
        RECT 1410.450 1763.440 1410.730 1763.720 ;
        RECT 1409.990 1758.680 1410.270 1758.960 ;
        RECT 1414.130 2066.040 1414.410 2066.320 ;
        RECT 1414.130 2055.840 1414.410 2056.120 ;
        RECT 1415.050 2046.320 1415.330 2046.600 ;
        RECT 1414.590 2042.240 1414.870 2042.520 ;
        RECT 1412.290 1966.080 1412.570 1966.360 ;
        RECT 1411.830 1772.960 1412.110 1773.240 ;
        RECT 1414.130 2021.160 1414.410 2021.440 ;
        RECT 1414.130 1945.000 1414.410 1945.280 ;
        RECT 1414.130 1915.080 1414.410 1915.360 ;
        RECT 1414.130 1899.440 1414.410 1899.720 ;
        RECT 1414.130 1894.680 1414.410 1894.960 ;
        RECT 1414.130 1889.920 1414.410 1890.200 ;
        RECT 1414.130 1879.720 1414.410 1880.000 ;
        RECT 1414.130 1874.280 1414.410 1874.560 ;
        RECT 1414.130 1869.520 1414.410 1869.800 ;
        RECT 1414.130 1859.320 1414.410 1859.600 ;
        RECT 1414.130 1854.560 1414.410 1854.840 ;
        RECT 1414.130 1844.360 1414.410 1844.640 ;
        RECT 1414.130 1838.920 1414.410 1839.200 ;
        RECT 1414.130 1834.160 1414.410 1834.440 ;
        RECT 1414.130 1823.960 1414.410 1824.240 ;
        RECT 1414.130 1819.200 1414.410 1819.480 ;
        RECT 1414.130 1813.760 1414.410 1814.040 ;
        RECT 1413.670 1809.000 1413.950 1809.280 ;
        RECT 1414.130 1798.800 1414.410 1799.080 ;
        RECT 1413.670 1794.040 1413.950 1794.320 ;
        RECT 1413.210 1768.200 1413.490 1768.480 ;
        RECT 1412.750 1753.240 1413.030 1753.520 ;
        RECT 1411.370 1748.480 1411.650 1748.760 ;
        RECT 1414.130 1743.040 1414.410 1743.320 ;
        RECT 1414.130 1738.280 1414.410 1738.560 ;
        RECT 1411.370 1732.840 1411.650 1733.120 ;
        RECT 1410.450 1728.080 1410.730 1728.360 ;
        RECT 1414.130 1723.320 1414.410 1723.600 ;
        RECT 1413.670 1717.880 1413.950 1718.160 ;
        RECT 1412.750 1713.120 1413.030 1713.400 ;
        RECT 1414.130 1707.680 1414.410 1707.960 ;
        RECT 1412.290 1702.920 1412.570 1703.200 ;
        RECT 1410.450 1698.160 1410.730 1698.440 ;
        RECT 1409.990 1682.520 1410.270 1682.800 ;
        RECT 1409.070 1672.320 1409.350 1672.600 ;
        RECT 1408.150 1667.560 1408.430 1667.840 ;
        RECT 1408.150 1652.600 1408.430 1652.880 ;
        RECT 1407.690 1647.160 1407.970 1647.440 ;
        RECT 1408.150 1642.400 1408.430 1642.680 ;
        RECT 1407.690 1636.960 1407.970 1637.240 ;
        RECT 1407.690 1632.200 1407.970 1632.480 ;
        RECT 1409.530 1657.360 1409.810 1657.640 ;
        RECT 1411.830 1692.720 1412.110 1693.000 ;
        RECT 1410.910 1662.800 1411.190 1663.080 ;
        RECT 1408.610 1627.440 1408.890 1627.720 ;
        RECT 1407.690 1622.000 1407.970 1622.280 ;
        RECT 1407.690 1617.240 1407.970 1617.520 ;
        RECT 1407.690 1611.800 1407.970 1612.080 ;
        RECT 1412.750 1687.960 1413.030 1688.240 ;
        RECT 1413.210 1677.760 1413.490 1678.040 ;
        RECT 1535.570 3231.560 1535.850 3231.840 ;
        RECT 1535.570 3224.760 1535.850 3225.040 ;
        RECT 1535.570 3217.280 1535.850 3217.560 ;
        RECT 1538.330 3210.480 1538.610 3210.760 ;
        RECT 1538.330 3202.320 1538.610 3202.600 ;
        RECT 1533.270 3196.880 1533.550 3197.160 ;
        RECT 1534.190 3189.400 1534.470 3189.680 ;
        RECT 1535.110 2898.360 1535.390 2898.640 ;
        RECT 1528.210 2891.560 1528.490 2891.840 ;
        RECT 1932.090 3249.240 1932.370 3249.520 ;
        RECT 1938.990 2948.000 1939.270 2948.280 ;
        RECT 1945.890 2904.480 1946.170 2904.760 ;
        RECT 1645.510 2799.080 1645.790 2799.360 ;
        RECT 1688.750 2799.080 1689.030 2799.360 ;
        RECT 1788.570 2799.080 1788.850 2799.360 ;
        RECT 1607.790 2794.320 1608.070 2794.600 ;
        RECT 1614.690 2794.320 1614.970 2794.600 ;
        RECT 1621.590 2794.320 1621.870 2794.600 ;
        RECT 1628.490 2794.320 1628.770 2794.600 ;
        RECT 1635.390 2794.320 1635.670 2794.600 ;
        RECT 1587.090 2789.560 1587.370 2789.840 ;
        RECT 1600.890 2789.560 1601.170 2789.840 ;
        RECT 1580.190 2787.520 1580.470 2787.800 ;
        RECT 1593.990 2787.520 1594.270 2787.800 ;
        RECT 1601.350 2787.520 1601.630 2787.800 ;
        RECT 1611.010 2793.640 1611.290 2793.920 ;
        RECT 1617.910 2793.640 1618.190 2793.920 ;
        RECT 1624.810 2793.640 1625.090 2793.920 ;
        RECT 1631.710 2793.640 1631.990 2793.920 ;
        RECT 1638.610 2793.640 1638.890 2793.920 ;
        RECT 1642.290 2793.640 1642.570 2793.920 ;
        RECT 1642.290 2792.280 1642.570 2792.560 ;
        RECT 1642.290 2785.480 1642.570 2785.760 ;
        RECT 1646.430 2794.320 1646.710 2794.600 ;
        RECT 1649.190 2794.320 1649.470 2794.600 ;
        RECT 1652.410 2794.320 1652.690 2794.600 ;
        RECT 1656.090 2794.320 1656.370 2794.600 ;
        RECT 1662.990 2794.320 1663.270 2794.600 ;
        RECT 1669.890 2794.320 1670.170 2794.600 ;
        RECT 1676.790 2794.320 1677.070 2794.600 ;
        RECT 1649.650 2793.640 1649.930 2793.920 ;
        RECT 1658.850 2793.640 1659.130 2793.920 ;
        RECT 1663.450 2793.640 1663.730 2793.920 ;
        RECT 1670.350 2793.640 1670.630 2793.920 ;
        RECT 1683.690 2794.320 1683.970 2794.600 ;
        RECT 1677.250 2793.640 1677.530 2793.920 ;
        RECT 1682.310 2793.640 1682.590 2793.920 ;
        RECT 1740.730 2796.360 1741.010 2796.640 ;
        RECT 1740.270 2795.680 1740.550 2795.960 ;
        RECT 1690.590 2794.320 1690.870 2794.600 ;
        RECT 1697.490 2794.320 1697.770 2794.600 ;
        RECT 1706.230 2794.320 1706.510 2794.600 ;
        RECT 1712.670 2794.320 1712.950 2794.600 ;
        RECT 1718.190 2794.320 1718.470 2794.600 ;
        RECT 1724.170 2794.320 1724.450 2794.600 ;
        RECT 1728.770 2794.320 1729.050 2794.600 ;
        RECT 1734.290 2794.320 1734.570 2794.600 ;
        RECT 1690.130 2793.640 1690.410 2793.920 ;
        RECT 1690.130 2792.280 1690.410 2792.560 ;
        RECT 1684.150 2789.560 1684.430 2789.840 ;
        RECT 1690.130 1949.080 1690.410 1949.360 ;
        RECT 1686.910 1906.240 1687.190 1906.520 ;
        RECT 1414.130 1607.040 1414.410 1607.320 ;
        RECT 1695.190 2793.640 1695.470 2793.920 ;
        RECT 1699.330 2793.640 1699.610 2793.920 ;
        RECT 1728.310 2792.280 1728.590 2792.560 ;
        RECT 1740.270 2792.960 1740.550 2793.240 ;
        RECT 1741.190 2794.320 1741.470 2794.600 ;
        RECT 1747.630 2794.320 1747.910 2794.600 ;
        RECT 1758.670 2794.320 1758.950 2794.600 ;
        RECT 1752.690 2792.280 1752.970 2792.560 ;
        RECT 1766.490 2793.640 1766.770 2793.920 ;
        RECT 1773.390 2793.640 1773.670 2793.920 ;
        RECT 1780.290 2793.640 1780.570 2793.920 ;
        RECT 1787.190 2792.280 1787.470 2792.560 ;
        RECT 1758.670 2790.920 1758.950 2791.200 ;
        RECT 1759.590 2790.920 1759.870 2791.200 ;
        RECT 1773.390 2790.920 1773.670 2791.200 ;
        RECT 1728.310 2790.240 1728.590 2790.520 ;
        RECT 1759.590 2790.240 1759.870 2790.520 ;
        RECT 1766.490 2789.560 1766.770 2789.840 ;
        RECT 1718.650 2788.200 1718.930 2788.480 ;
        RECT 1704.390 2787.520 1704.670 2787.800 ;
        RECT 1711.290 2787.520 1711.570 2787.800 ;
        RECT 1718.190 2787.520 1718.470 2787.800 ;
        RECT 1725.090 2787.520 1725.370 2787.800 ;
        RECT 1731.990 2787.520 1732.270 2787.800 ;
        RECT 1738.890 2787.520 1739.170 2787.800 ;
        RECT 1745.790 2787.520 1746.070 2787.800 ;
        RECT 1753.150 2787.520 1753.430 2787.800 ;
        RECT 1835.490 2069.440 1835.770 2069.720 ;
        RECT 1842.390 2069.440 1842.670 2069.720 ;
        RECT 1849.290 2069.440 1849.570 2069.720 ;
        RECT 1856.190 2069.440 1856.470 2069.720 ;
        RECT 1863.090 2069.440 1863.370 2069.720 ;
        RECT 1869.990 2069.440 1870.270 2069.720 ;
        RECT 1876.890 2069.440 1877.170 2069.720 ;
        RECT 1883.790 2069.440 1884.070 2069.720 ;
        RECT 1890.690 2069.440 1890.970 2069.720 ;
        RECT 1897.590 2069.440 1897.870 2069.720 ;
        RECT 1904.490 2069.440 1904.770 2069.720 ;
        RECT 1911.390 2069.440 1911.670 2069.720 ;
        RECT 1870.450 2068.760 1870.730 2069.040 ;
        RECT 1841.470 2066.720 1841.750 2067.000 ;
        RECT 1843.770 2066.720 1844.050 2067.000 ;
        RECT 1911.850 2068.760 1912.130 2069.040 ;
        RECT 1848.830 2066.720 1849.110 2067.000 ;
        RECT 1849.290 2066.040 1849.570 2066.320 ;
        RECT 1890.230 2066.720 1890.510 2067.000 ;
        RECT 1898.050 2066.040 1898.330 2066.320 ;
        RECT 1859.870 2065.360 1860.150 2065.640 ;
        RECT 1864.930 2065.360 1865.210 2065.640 ;
        RECT 1893.910 2065.360 1894.190 2065.640 ;
        RECT 1907.710 2065.360 1907.990 2065.640 ;
        RECT 1911.390 2065.360 1911.670 2065.640 ;
        RECT 1871.830 2064.680 1872.110 2064.960 ;
        RECT 1925.190 2069.440 1925.470 2069.720 ;
        RECT 1919.210 2068.760 1919.490 2069.040 ;
        RECT 1932.090 2066.040 1932.370 2066.320 ;
        RECT 1941.750 2066.720 1942.030 2067.000 ;
        RECT 1936.690 2065.360 1936.970 2065.640 ;
        RECT 1917.830 2064.680 1918.110 2064.960 ;
        RECT 1924.730 2064.680 1925.010 2064.960 ;
        RECT 1930.250 2064.680 1930.530 2064.960 ;
        RECT 1980.390 2068.080 1980.670 2068.360 ;
        RECT 1987.290 2068.080 1987.570 2068.360 ;
        RECT 2028.690 2067.400 2028.970 2067.680 ;
        RECT 1877.350 2064.000 1877.630 2064.280 ;
        RECT 1882.870 2064.000 1883.150 2064.280 ;
        RECT 1966.590 2064.000 1966.870 2064.280 ;
        RECT 2021.790 2066.720 2022.070 2067.000 ;
        RECT 2007.990 2066.040 2008.270 2066.320 ;
        RECT 2015.810 2066.040 2016.090 2066.320 ;
        RECT 2035.590 2066.040 2035.870 2066.320 ;
        RECT 1994.190 2065.360 1994.470 2065.640 ;
        RECT 2042.490 2065.360 2042.770 2065.640 ;
        RECT 2001.090 2064.680 2001.370 2064.960 ;
        RECT 1987.290 2064.000 1987.570 2064.280 ;
        RECT 1948.190 2063.320 1948.470 2063.600 ;
        RECT 1954.630 2063.320 1954.910 2063.600 ;
        RECT 1958.770 2063.320 1959.050 2063.600 ;
        RECT 1965.670 2063.320 1965.950 2063.600 ;
        RECT 1969.810 2063.320 1970.090 2063.600 ;
        RECT 1973.490 2063.320 1973.770 2063.600 ;
        RECT 1976.710 2063.320 1976.990 2063.600 ;
        RECT 1980.390 2063.320 1980.670 2063.600 ;
        RECT 2028.690 2063.320 2028.970 2063.600 ;
        RECT 1940.370 2058.560 1940.650 2058.840 ;
        RECT 1955.090 2057.880 1955.370 2058.160 ;
        RECT 1987.290 2057.880 1987.570 2058.160 ;
        RECT 1995.570 2057.880 1995.850 2058.160 ;
        RECT 1946.350 2057.200 1946.630 2057.480 ;
        RECT 1990.050 2057.200 1990.330 2057.480 ;
        RECT 2004.770 2057.200 2005.050 2057.480 ;
        RECT 2016.270 2057.200 2016.550 2057.480 ;
        RECT 2008.450 2056.520 2008.730 2056.800 ;
        RECT 2021.790 2056.520 2022.070 2056.800 ;
        RECT 1948.650 2055.160 1948.930 2055.440 ;
        RECT 1961.530 2051.760 1961.810 2052.040 ;
        RECT 2049.850 2051.760 2050.130 2052.040 ;
        RECT 1688.750 1609.760 1689.030 1610.040 ;
        RECT 2097.690 1964.720 2097.970 1965.000 ;
        RECT 2097.690 1953.160 2097.970 1953.440 ;
        RECT 2082.050 1619.960 2082.330 1620.240 ;
        RECT 1414.130 1603.640 1414.410 1603.920 ;
        RECT 2099.530 1662.800 2099.810 1663.080 ;
        RECT 2099.070 1643.080 2099.350 1643.360 ;
        RECT 2098.610 1635.600 2098.890 1635.880 ;
        RECT 2098.150 1628.800 2098.430 1629.080 ;
        RECT 2100.910 1656.000 2101.190 1656.280 ;
        RECT 2099.990 1649.200 2100.270 1649.480 ;
        RECT 1720.030 1593.440 1720.310 1593.720 ;
        RECT 1738.890 1592.080 1739.170 1592.360 ;
      LAYER met3 ;
        RECT 646.365 3264.500 646.695 3264.505 ;
        RECT 668.445 3264.500 668.775 3264.505 ;
        RECT 1293.125 3264.500 1293.455 3264.505 ;
        RECT 646.110 3264.490 646.695 3264.500 ;
        RECT 668.190 3264.490 668.775 3264.500 ;
        RECT 1292.870 3264.490 1293.455 3264.500 ;
        RECT 645.910 3264.190 646.695 3264.490 ;
        RECT 667.990 3264.190 668.775 3264.490 ;
        RECT 1292.670 3264.190 1293.455 3264.490 ;
        RECT 646.110 3264.180 646.695 3264.190 ;
        RECT 668.190 3264.180 668.775 3264.190 ;
        RECT 1292.870 3264.180 1293.455 3264.190 ;
        RECT 646.365 3264.175 646.695 3264.180 ;
        RECT 668.445 3264.175 668.775 3264.180 ;
        RECT 1293.125 3264.175 1293.455 3264.180 ;
        RECT 1890.665 3264.500 1890.995 3264.505 ;
        RECT 1917.345 3264.500 1917.675 3264.505 ;
        RECT 1890.665 3264.490 1891.250 3264.500 ;
        RECT 1917.345 3264.490 1917.930 3264.500 ;
        RECT 1890.665 3264.190 1891.450 3264.490 ;
        RECT 1917.345 3264.190 1918.130 3264.490 ;
        RECT 1890.665 3264.180 1891.250 3264.190 ;
        RECT 1917.345 3264.180 1917.930 3264.190 ;
        RECT 1890.665 3264.175 1890.995 3264.180 ;
        RECT 1917.345 3264.175 1917.675 3264.180 ;
        RECT 1317.505 3258.380 1317.835 3258.385 ;
        RECT 1317.505 3258.370 1318.205 3258.380 ;
        RECT 1317.505 3258.070 1318.290 3258.370 ;
        RECT 1317.505 3258.060 1318.205 3258.070 ;
        RECT 1317.505 3258.055 1317.835 3258.060 ;
        RECT 1186.865 3252.930 1187.195 3252.945 ;
        RECT 1187.785 3252.930 1188.115 3252.945 ;
        RECT 1186.865 3252.630 1188.115 3252.930 ;
        RECT 1186.865 3252.615 1187.195 3252.630 ;
        RECT 1187.785 3252.615 1188.115 3252.630 ;
        RECT 659.280 3251.235 661.020 3252.140 ;
        RECT 1309.280 3251.235 1311.020 3252.140 ;
        RECT 1909.280 3251.235 1911.020 3252.140 ;
        RECT 300.000 3232.785 304.600 3233.085 ;
        RECT 288.025 3230.490 288.355 3230.505 ;
        RECT 300.230 3230.490 300.530 3232.785 ;
        RECT 288.025 3230.190 300.530 3230.490 ;
        RECT 288.025 3230.175 288.355 3230.190 ;
        RECT 300.000 3227.145 304.600 3227.445 ;
        RECT 287.565 3225.050 287.895 3225.065 ;
        RECT 300.230 3225.050 300.530 3227.145 ;
        RECT 287.565 3224.750 300.530 3225.050 ;
        RECT 287.565 3224.735 287.895 3224.750 ;
        RECT 300.000 3218.645 304.600 3218.945 ;
        RECT 287.105 3216.210 287.435 3216.225 ;
        RECT 300.230 3216.210 300.530 3218.645 ;
        RECT 287.105 3215.910 300.530 3216.210 ;
        RECT 287.105 3215.895 287.435 3215.910 ;
        RECT 300.000 3213.005 304.600 3213.305 ;
        RECT 286.645 3210.090 286.975 3210.105 ;
        RECT 300.230 3210.090 300.530 3213.005 ;
        RECT 286.645 3209.790 300.530 3210.090 ;
        RECT 286.645 3209.775 286.975 3209.790 ;
        RECT 300.000 3204.505 304.600 3204.805 ;
        RECT 286.185 3201.930 286.515 3201.945 ;
        RECT 300.230 3201.930 300.530 3204.505 ;
        RECT 286.185 3201.630 300.530 3201.930 ;
        RECT 286.185 3201.615 286.515 3201.630 ;
        RECT 300.000 3198.865 304.600 3199.165 ;
        RECT 285.265 3196.490 285.595 3196.505 ;
        RECT 300.230 3196.490 300.530 3198.865 ;
        RECT 285.265 3196.190 300.530 3196.490 ;
        RECT 285.265 3196.175 285.595 3196.190 ;
        RECT 300.000 3190.365 304.600 3190.665 ;
        RECT 285.725 3188.330 286.055 3188.345 ;
        RECT 300.230 3188.330 300.530 3190.365 ;
        RECT 285.725 3188.030 300.530 3188.330 ;
        RECT 285.725 3188.015 286.055 3188.030 ;
        RECT 300.000 2901.125 304.600 2901.425 ;
        RECT 284.805 2898.650 285.135 2898.665 ;
        RECT 300.230 2898.650 300.530 2901.125 ;
        RECT 284.805 2898.350 300.530 2898.650 ;
        RECT 284.805 2898.335 285.135 2898.350 ;
        RECT 300.000 2892.625 304.600 2892.925 ;
        RECT 284.345 2891.850 284.675 2891.865 ;
        RECT 300.230 2891.850 300.530 2892.625 ;
        RECT 284.345 2891.550 300.530 2891.850 ;
        RECT 284.345 2891.535 284.675 2891.550 ;
      LAYER met3 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
      LAYER met3 ;
        RECT 688.225 3248.565 688.555 3248.580 ;
        RECT 681.880 3248.265 688.555 3248.565 ;
        RECT 688.225 3248.250 688.555 3248.265 ;
        RECT 950.000 3232.785 954.600 3233.085 ;
        RECT 941.685 3230.490 942.015 3230.505 ;
        RECT 950.670 3230.490 950.970 3232.785 ;
        RECT 941.685 3230.190 950.970 3230.490 ;
        RECT 941.685 3230.175 942.015 3230.190 ;
        RECT 950.000 3227.145 954.600 3227.445 ;
        RECT 942.145 3225.050 942.475 3225.065 ;
        RECT 950.670 3225.050 950.970 3227.145 ;
        RECT 942.145 3224.750 950.970 3225.050 ;
        RECT 942.145 3224.735 942.475 3224.750 ;
        RECT 950.000 3218.645 954.600 3218.945 ;
        RECT 942.605 3216.210 942.935 3216.225 ;
        RECT 950.670 3216.210 950.970 3218.645 ;
        RECT 942.605 3215.910 950.970 3216.210 ;
        RECT 942.605 3215.895 942.935 3215.910 ;
        RECT 950.000 3213.005 954.600 3213.305 ;
        RECT 943.065 3210.090 943.395 3210.105 ;
        RECT 950.670 3210.090 950.970 3213.005 ;
        RECT 943.065 3209.790 950.970 3210.090 ;
        RECT 943.065 3209.775 943.395 3209.790 ;
        RECT 950.000 3204.505 954.600 3204.805 ;
        RECT 943.525 3201.930 943.855 3201.945 ;
        RECT 950.670 3201.930 950.970 3204.505 ;
        RECT 943.525 3201.630 950.970 3201.930 ;
        RECT 943.525 3201.615 943.855 3201.630 ;
        RECT 950.000 3198.865 954.600 3199.165 ;
        RECT 944.445 3196.490 944.775 3196.505 ;
        RECT 950.670 3196.490 950.970 3198.865 ;
        RECT 944.445 3196.190 950.970 3196.490 ;
        RECT 944.445 3196.175 944.775 3196.190 ;
        RECT 950.000 3190.365 954.600 3190.665 ;
        RECT 941.225 3188.330 941.555 3188.345 ;
        RECT 950.670 3188.330 950.970 3190.365 ;
        RECT 941.225 3188.030 950.970 3188.330 ;
        RECT 941.225 3188.015 941.555 3188.030 ;
        RECT 696.965 2948.290 697.295 2948.305 ;
        RECT 684.790 2947.990 697.295 2948.290 ;
        RECT 684.790 2947.210 685.090 2947.990 ;
        RECT 696.965 2947.975 697.295 2947.990 ;
        RECT 681.880 2946.910 686.480 2947.210 ;
        RECT 684.790 2938.710 685.090 2946.910 ;
        RECT 681.880 2938.410 686.480 2938.710 ;
        RECT 684.790 2933.070 685.090 2938.410 ;
        RECT 681.880 2932.770 686.480 2933.070 ;
        RECT 685.710 2924.570 686.010 2932.770 ;
        RECT 681.880 2924.270 686.480 2924.570 ;
        RECT 685.710 2918.930 686.010 2924.270 ;
        RECT 681.880 2918.630 686.480 2918.930 ;
        RECT 685.710 2910.430 686.010 2918.630 ;
        RECT 681.880 2910.130 686.480 2910.430 ;
        RECT 685.710 2904.790 686.010 2910.130 ;
        RECT 681.880 2904.490 686.480 2904.790 ;
        RECT 950.000 2901.125 954.600 2901.425 ;
        RECT 943.985 2898.650 944.315 2898.665 ;
        RECT 950.670 2898.650 950.970 2901.125 ;
        RECT 943.985 2898.350 950.970 2898.650 ;
        RECT 943.985 2898.335 944.315 2898.350 ;
        RECT 950.000 2892.625 954.600 2892.925 ;
        RECT 944.905 2891.850 945.235 2891.865 ;
        RECT 950.670 2891.850 950.970 2892.625 ;
        RECT 944.905 2891.550 950.970 2891.850 ;
        RECT 944.905 2891.535 945.235 2891.550 ;
      LAYER met3 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
      LAYER met3 ;
        RECT 1352.465 3250.210 1352.795 3250.225 ;
        RECT 1400.305 3250.210 1400.635 3250.225 ;
        RECT 1352.465 3249.910 1400.635 3250.210 ;
        RECT 1352.465 3249.895 1352.795 3249.910 ;
        RECT 1400.305 3249.895 1400.635 3249.910 ;
        RECT 1332.225 3249.530 1332.555 3249.545 ;
        RECT 1332.225 3249.215 1332.770 3249.530 ;
        RECT 1332.470 3248.565 1332.770 3249.215 ;
        RECT 1331.880 3248.265 1336.480 3248.565 ;
        RECT 1550.000 3232.785 1554.600 3233.085 ;
        RECT 1535.545 3231.850 1535.875 3231.865 ;
        RECT 1550.510 3231.850 1550.810 3232.785 ;
        RECT 1535.545 3231.550 1550.810 3231.850 ;
        RECT 1535.545 3231.535 1535.875 3231.550 ;
        RECT 1550.000 3227.145 1554.600 3227.445 ;
        RECT 1535.545 3225.050 1535.875 3225.065 ;
        RECT 1550.510 3225.050 1550.810 3227.145 ;
        RECT 1535.545 3224.750 1550.810 3225.050 ;
        RECT 1535.545 3224.735 1535.875 3224.750 ;
        RECT 1550.000 3218.645 1554.600 3218.945 ;
        RECT 1535.545 3217.570 1535.875 3217.585 ;
        RECT 1550.510 3217.570 1550.810 3218.645 ;
        RECT 1535.545 3217.270 1550.810 3217.570 ;
        RECT 1535.545 3217.255 1535.875 3217.270 ;
        RECT 1550.000 3213.005 1554.600 3213.305 ;
        RECT 1538.305 3210.770 1538.635 3210.785 ;
        RECT 1550.510 3210.770 1550.810 3213.005 ;
        RECT 1538.305 3210.470 1550.810 3210.770 ;
        RECT 1538.305 3210.455 1538.635 3210.470 ;
        RECT 1550.000 3204.505 1554.600 3204.805 ;
        RECT 1538.305 3202.610 1538.635 3202.625 ;
        RECT 1550.510 3202.610 1550.810 3204.505 ;
        RECT 1538.305 3202.310 1550.810 3202.610 ;
        RECT 1538.305 3202.295 1538.635 3202.310 ;
        RECT 1550.000 3198.865 1554.600 3199.165 ;
        RECT 1533.245 3197.170 1533.575 3197.185 ;
        RECT 1550.510 3197.170 1550.810 3198.865 ;
        RECT 1533.245 3196.870 1550.810 3197.170 ;
        RECT 1533.245 3196.855 1533.575 3196.870 ;
        RECT 1550.000 3190.365 1554.600 3190.665 ;
        RECT 1534.165 3189.690 1534.495 3189.705 ;
        RECT 1550.510 3189.690 1550.810 3190.365 ;
        RECT 1534.165 3189.390 1550.810 3189.690 ;
        RECT 1534.165 3189.375 1534.495 3189.390 ;
        RECT 1331.880 2946.930 1336.480 2947.210 ;
        RECT 1345.565 2946.930 1345.895 2946.945 ;
        RECT 1352.005 2946.930 1352.335 2946.945 ;
        RECT 1331.880 2946.910 1352.335 2946.930 ;
        RECT 1336.150 2946.630 1352.335 2946.910 ;
        RECT 1345.565 2946.615 1345.895 2946.630 ;
        RECT 1352.005 2946.615 1352.335 2946.630 ;
        RECT 1345.565 2938.770 1345.895 2938.785 ;
        RECT 1336.150 2938.710 1345.895 2938.770 ;
        RECT 1331.880 2938.470 1345.895 2938.710 ;
        RECT 1331.880 2938.410 1336.480 2938.470 ;
        RECT 1345.565 2938.455 1345.895 2938.470 ;
        RECT 1336.150 2933.070 1336.450 2938.410 ;
        RECT 1331.880 2932.770 1336.480 2933.070 ;
        RECT 1336.150 2924.570 1336.450 2932.770 ;
        RECT 1331.880 2924.270 1336.480 2924.570 ;
        RECT 1336.150 2918.930 1336.450 2924.270 ;
        RECT 1331.880 2918.630 1336.480 2918.930 ;
        RECT 1336.150 2910.430 1336.450 2918.630 ;
        RECT 1331.880 2910.130 1336.480 2910.430 ;
        RECT 1336.150 2904.790 1336.450 2910.130 ;
        RECT 1331.880 2904.490 1336.480 2904.790 ;
        RECT 1550.000 2901.125 1554.600 2901.425 ;
        RECT 1535.085 2898.650 1535.415 2898.665 ;
        RECT 1550.510 2898.650 1550.810 2901.125 ;
        RECT 1535.085 2898.350 1550.810 2898.650 ;
        RECT 1535.085 2898.335 1535.415 2898.350 ;
        RECT 1550.000 2892.625 1554.600 2892.925 ;
        RECT 1528.185 2891.850 1528.515 2891.865 ;
        RECT 1550.510 2891.850 1550.810 2892.625 ;
        RECT 1528.185 2891.550 1550.810 2891.850 ;
        RECT 1528.185 2891.535 1528.515 2891.550 ;
      LAYER met3 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met3 ;
        RECT 1932.065 3249.530 1932.395 3249.545 ;
        RECT 1932.065 3249.215 1932.610 3249.530 ;
        RECT 1932.310 3248.565 1932.610 3249.215 ;
        RECT 1931.880 3248.265 1936.480 3248.565 ;
        RECT 1938.965 2948.290 1939.295 2948.305 ;
        RECT 1935.070 2947.990 1939.295 2948.290 ;
        RECT 1935.070 2947.210 1935.370 2947.990 ;
        RECT 1938.965 2947.975 1939.295 2947.990 ;
        RECT 1931.880 2946.910 1936.480 2947.210 ;
        RECT 1935.070 2938.710 1935.370 2946.910 ;
        RECT 1931.880 2938.410 1936.480 2938.710 ;
        RECT 1935.070 2933.070 1935.370 2938.410 ;
        RECT 1931.880 2932.770 1936.480 2933.070 ;
        RECT 1935.990 2924.570 1936.290 2932.770 ;
        RECT 1931.880 2924.270 1936.480 2924.570 ;
        RECT 1935.990 2918.930 1936.290 2924.270 ;
        RECT 1931.880 2918.630 1936.480 2918.930 ;
        RECT 1935.990 2910.430 1936.290 2918.630 ;
        RECT 1931.880 2910.130 1936.480 2910.430 ;
        RECT 1935.990 2904.790 1936.290 2910.130 ;
        RECT 1931.880 2904.770 1936.480 2904.790 ;
        RECT 1945.865 2904.770 1946.195 2904.785 ;
        RECT 1931.880 2904.490 1946.195 2904.770 ;
        RECT 1935.990 2904.470 1946.195 2904.490 ;
        RECT 1945.865 2904.455 1946.195 2904.470 ;
        RECT 1054.845 2800.050 1055.175 2800.065 ;
        RECT 1055.510 2800.050 1055.890 2800.060 ;
        RECT 1054.845 2799.750 1055.890 2800.050 ;
        RECT 1054.845 2799.735 1055.175 2799.750 ;
        RECT 1055.510 2799.740 1055.890 2799.750 ;
        RECT 1642.370 2799.370 1642.750 2799.380 ;
        RECT 1645.485 2799.370 1645.815 2799.385 ;
        RECT 1688.725 2799.380 1689.055 2799.385 ;
        RECT 1688.470 2799.370 1689.055 2799.380 ;
        RECT 1788.545 2799.370 1788.875 2799.385 ;
        RECT 1794.210 2799.370 1794.590 2799.380 ;
        RECT 1642.370 2799.070 1689.460 2799.370 ;
        RECT 1788.545 2799.070 1794.590 2799.370 ;
        RECT 1642.370 2799.060 1642.750 2799.070 ;
        RECT 1645.485 2799.055 1645.815 2799.070 ;
        RECT 1688.470 2799.060 1689.055 2799.070 ;
        RECT 1688.725 2799.055 1689.055 2799.060 ;
        RECT 1788.545 2799.055 1788.875 2799.070 ;
        RECT 1794.210 2799.060 1794.590 2799.070 ;
        RECT 1794.270 2798.690 1794.650 2798.700 ;
        RECT 1797.030 2798.690 1797.410 2798.700 ;
        RECT 1794.270 2798.390 1797.410 2798.690 ;
        RECT 1794.270 2798.380 1794.650 2798.390 ;
        RECT 1797.030 2798.380 1797.410 2798.390 ;
        RECT 1740.705 2796.650 1741.035 2796.665 ;
        RECT 1759.310 2796.650 1759.690 2796.660 ;
        RECT 1740.705 2796.350 1759.690 2796.650 ;
        RECT 1740.705 2796.335 1741.035 2796.350 ;
        RECT 1759.310 2796.340 1759.690 2796.350 ;
        RECT 1740.245 2795.970 1740.575 2795.985 ;
        RECT 1761.150 2795.970 1761.530 2795.980 ;
        RECT 1740.245 2795.670 1761.530 2795.970 ;
        RECT 1740.245 2795.655 1740.575 2795.670 ;
        RECT 1761.150 2795.660 1761.530 2795.670 ;
        RECT 1100.385 2795.300 1100.715 2795.305 ;
        RECT 1100.385 2795.290 1100.970 2795.300 ;
        RECT 1100.385 2794.990 1101.170 2795.290 ;
        RECT 1100.385 2794.980 1100.970 2794.990 ;
        RECT 1100.385 2794.975 1100.715 2794.980 ;
        RECT 336.990 2794.610 337.370 2794.620 ;
        RECT 337.705 2794.610 338.035 2794.625 ;
        RECT 336.990 2794.310 338.035 2794.610 ;
        RECT 336.990 2794.300 337.370 2794.310 ;
        RECT 337.705 2794.295 338.035 2794.310 ;
        RECT 342.510 2794.610 342.890 2794.620 ;
        RECT 344.605 2794.610 344.935 2794.625 ;
        RECT 342.510 2794.310 344.935 2794.610 ;
        RECT 342.510 2794.300 342.890 2794.310 ;
        RECT 344.605 2794.295 344.935 2794.310 ;
        RECT 350.790 2794.610 351.170 2794.620 ;
        RECT 351.505 2794.610 351.835 2794.625 ;
        RECT 358.405 2794.620 358.735 2794.625 ;
        RECT 350.790 2794.310 351.835 2794.610 ;
        RECT 350.790 2794.300 351.170 2794.310 ;
        RECT 351.505 2794.295 351.835 2794.310 ;
        RECT 358.150 2794.610 358.735 2794.620 ;
        RECT 361.830 2794.610 362.210 2794.620 ;
        RECT 363.005 2794.610 363.335 2794.625 ;
        RECT 358.150 2794.310 358.960 2794.610 ;
        RECT 361.830 2794.310 363.335 2794.610 ;
        RECT 358.150 2794.300 358.735 2794.310 ;
        RECT 361.830 2794.300 362.210 2794.310 ;
        RECT 358.405 2794.295 358.735 2794.300 ;
        RECT 363.005 2794.295 363.335 2794.310 ;
        RECT 364.590 2794.610 364.970 2794.620 ;
        RECT 365.305 2794.610 365.635 2794.625 ;
        RECT 364.590 2794.310 365.635 2794.610 ;
        RECT 364.590 2794.300 364.970 2794.310 ;
        RECT 365.305 2794.295 365.635 2794.310 ;
        RECT 368.270 2794.610 368.650 2794.620 ;
        RECT 368.985 2794.610 369.315 2794.625 ;
        RECT 371.285 2794.620 371.615 2794.625 ;
        RECT 374.965 2794.620 375.295 2794.625 ;
        RECT 371.030 2794.610 371.615 2794.620 ;
        RECT 374.710 2794.610 375.295 2794.620 ;
        RECT 368.270 2794.310 369.315 2794.610 ;
        RECT 370.830 2794.310 371.615 2794.610 ;
        RECT 374.510 2794.310 375.295 2794.610 ;
        RECT 368.270 2794.300 368.650 2794.310 ;
        RECT 368.985 2794.295 369.315 2794.310 ;
        RECT 371.030 2794.300 371.615 2794.310 ;
        RECT 374.710 2794.300 375.295 2794.310 ;
        RECT 379.310 2794.610 379.690 2794.620 ;
        RECT 380.025 2794.610 380.355 2794.625 ;
        RECT 384.165 2794.620 384.495 2794.625 ;
        RECT 386.925 2794.620 387.255 2794.625 ;
        RECT 392.445 2794.620 392.775 2794.625 ;
        RECT 383.910 2794.610 384.495 2794.620 ;
        RECT 386.670 2794.610 387.255 2794.620 ;
        RECT 392.190 2794.610 392.775 2794.620 ;
        RECT 379.310 2794.310 380.355 2794.610 ;
        RECT 383.710 2794.310 384.495 2794.610 ;
        RECT 386.470 2794.310 387.255 2794.610 ;
        RECT 391.990 2794.310 392.775 2794.610 ;
        RECT 379.310 2794.300 379.690 2794.310 ;
        RECT 371.285 2794.295 371.615 2794.300 ;
        RECT 374.965 2794.295 375.295 2794.300 ;
        RECT 380.025 2794.295 380.355 2794.310 ;
        RECT 383.910 2794.300 384.495 2794.310 ;
        RECT 386.670 2794.300 387.255 2794.310 ;
        RECT 392.190 2794.300 392.775 2794.310 ;
        RECT 395.870 2794.610 396.250 2794.620 ;
        RECT 397.045 2794.610 397.375 2794.625 ;
        RECT 399.805 2794.620 400.135 2794.625 ;
        RECT 399.550 2794.610 400.135 2794.620 ;
        RECT 395.870 2794.310 397.375 2794.610 ;
        RECT 399.350 2794.310 400.135 2794.610 ;
        RECT 395.870 2794.300 396.250 2794.310 ;
        RECT 384.165 2794.295 384.495 2794.300 ;
        RECT 386.925 2794.295 387.255 2794.300 ;
        RECT 392.445 2794.295 392.775 2794.300 ;
        RECT 397.045 2794.295 397.375 2794.310 ;
        RECT 399.550 2794.300 400.135 2794.310 ;
        RECT 403.230 2794.610 403.610 2794.620 ;
        RECT 403.945 2794.610 404.275 2794.625 ;
        RECT 406.245 2794.620 406.575 2794.625 ;
        RECT 405.990 2794.610 406.575 2794.620 ;
        RECT 403.230 2794.310 404.275 2794.610 ;
        RECT 405.790 2794.310 406.575 2794.610 ;
        RECT 403.230 2794.300 403.610 2794.310 ;
        RECT 399.805 2794.295 400.135 2794.300 ;
        RECT 403.945 2794.295 404.275 2794.310 ;
        RECT 405.990 2794.300 406.575 2794.310 ;
        RECT 406.245 2794.295 406.575 2794.300 ;
        RECT 409.465 2794.620 409.795 2794.625 ;
        RECT 413.605 2794.620 413.935 2794.625 ;
        RECT 419.125 2794.620 419.455 2794.625 ;
        RECT 420.965 2794.620 421.295 2794.625 ;
        RECT 409.465 2794.610 410.050 2794.620 ;
        RECT 413.350 2794.610 413.935 2794.620 ;
        RECT 418.870 2794.610 419.455 2794.620 ;
        RECT 409.465 2794.310 410.250 2794.610 ;
        RECT 413.350 2794.310 414.160 2794.610 ;
        RECT 418.670 2794.310 419.455 2794.610 ;
        RECT 409.465 2794.300 410.050 2794.310 ;
        RECT 413.350 2794.300 413.935 2794.310 ;
        RECT 418.870 2794.300 419.455 2794.310 ;
        RECT 420.710 2794.610 421.295 2794.620 ;
        RECT 425.310 2794.610 425.690 2794.620 ;
        RECT 427.405 2794.610 427.735 2794.625 ;
        RECT 432.005 2794.620 432.335 2794.625 ;
        RECT 431.750 2794.610 432.335 2794.620 ;
        RECT 420.710 2794.310 421.520 2794.610 ;
        RECT 425.310 2794.310 427.735 2794.610 ;
        RECT 431.550 2794.310 432.335 2794.610 ;
        RECT 420.710 2794.300 421.295 2794.310 ;
        RECT 425.310 2794.300 425.690 2794.310 ;
        RECT 409.465 2794.295 409.795 2794.300 ;
        RECT 413.605 2794.295 413.935 2794.300 ;
        RECT 419.125 2794.295 419.455 2794.300 ;
        RECT 420.965 2794.295 421.295 2794.300 ;
        RECT 427.405 2794.295 427.735 2794.310 ;
        RECT 431.750 2794.300 432.335 2794.310 ;
        RECT 433.590 2794.610 433.970 2794.620 ;
        RECT 434.305 2794.610 434.635 2794.625 ;
        RECT 439.365 2794.620 439.695 2794.625 ;
        RECT 441.205 2794.620 441.535 2794.625 ;
        RECT 439.110 2794.610 439.695 2794.620 ;
        RECT 433.590 2794.310 434.635 2794.610 ;
        RECT 438.910 2794.310 439.695 2794.610 ;
        RECT 433.590 2794.300 433.970 2794.310 ;
        RECT 432.005 2794.295 432.335 2794.300 ;
        RECT 434.305 2794.295 434.635 2794.310 ;
        RECT 439.110 2794.300 439.695 2794.310 ;
        RECT 440.950 2794.610 441.535 2794.620 ;
        RECT 444.425 2794.620 444.755 2794.625 ;
        RECT 444.425 2794.610 445.010 2794.620 ;
        RECT 440.950 2794.310 441.760 2794.610 ;
        RECT 444.200 2794.310 445.010 2794.610 ;
        RECT 440.950 2794.300 441.535 2794.310 ;
        RECT 439.365 2794.295 439.695 2794.300 ;
        RECT 441.205 2794.295 441.535 2794.300 ;
        RECT 444.425 2794.300 445.010 2794.310 ;
        RECT 445.550 2794.610 445.930 2794.620 ;
        RECT 448.105 2794.610 448.435 2794.625 ;
        RECT 445.550 2794.310 448.435 2794.610 ;
        RECT 445.550 2794.300 445.930 2794.310 ;
        RECT 444.425 2794.295 444.755 2794.300 ;
        RECT 448.105 2794.295 448.435 2794.310 ;
        RECT 449.025 2794.620 449.355 2794.625 ;
        RECT 455.005 2794.620 455.335 2794.625 ;
        RECT 462.365 2794.620 462.695 2794.625 ;
        RECT 449.025 2794.610 449.610 2794.620 ;
        RECT 454.750 2794.610 455.335 2794.620 ;
        RECT 462.110 2794.610 462.695 2794.620 ;
        RECT 449.025 2794.310 449.810 2794.610 ;
        RECT 454.750 2794.310 455.560 2794.610 ;
        RECT 461.910 2794.310 462.695 2794.610 ;
        RECT 449.025 2794.300 449.610 2794.310 ;
        RECT 454.750 2794.300 455.335 2794.310 ;
        RECT 462.110 2794.300 462.695 2794.310 ;
        RECT 465.790 2794.610 466.170 2794.620 ;
        RECT 468.345 2794.610 468.675 2794.625 ;
        RECT 474.325 2794.620 474.655 2794.625 ;
        RECT 474.070 2794.610 474.655 2794.620 ;
        RECT 465.790 2794.310 468.675 2794.610 ;
        RECT 473.870 2794.310 474.655 2794.610 ;
        RECT 465.790 2794.300 466.170 2794.310 ;
        RECT 449.025 2794.295 449.355 2794.300 ;
        RECT 455.005 2794.295 455.335 2794.300 ;
        RECT 462.365 2794.295 462.695 2794.300 ;
        RECT 468.345 2794.295 468.675 2794.310 ;
        RECT 474.070 2794.300 474.655 2794.310 ;
        RECT 474.990 2794.610 475.370 2794.620 ;
        RECT 475.705 2794.610 476.035 2794.625 ;
        RECT 478.925 2794.620 479.255 2794.625 ;
        RECT 482.605 2794.620 482.935 2794.625 ;
        RECT 478.670 2794.610 479.255 2794.620 ;
        RECT 474.990 2794.310 476.035 2794.610 ;
        RECT 478.470 2794.310 479.255 2794.610 ;
        RECT 474.990 2794.300 475.370 2794.310 ;
        RECT 474.325 2794.295 474.655 2794.300 ;
        RECT 475.705 2794.295 476.035 2794.310 ;
        RECT 478.670 2794.300 479.255 2794.310 ;
        RECT 482.350 2794.610 482.935 2794.620 ;
        RECT 484.905 2794.620 485.235 2794.625 ;
        RECT 489.045 2794.620 489.375 2794.625 ;
        RECT 484.905 2794.610 485.490 2794.620 ;
        RECT 488.790 2794.610 489.375 2794.620 ;
        RECT 482.350 2794.310 483.160 2794.610 ;
        RECT 484.905 2794.310 485.690 2794.610 ;
        RECT 488.590 2794.310 489.375 2794.610 ;
        RECT 482.350 2794.300 482.935 2794.310 ;
        RECT 478.925 2794.295 479.255 2794.300 ;
        RECT 482.605 2794.295 482.935 2794.300 ;
        RECT 484.905 2794.300 485.490 2794.310 ;
        RECT 488.790 2794.300 489.375 2794.310 ;
        RECT 484.905 2794.295 485.235 2794.300 ;
        RECT 489.045 2794.295 489.375 2794.300 ;
        RECT 490.425 2794.620 490.755 2794.625 ;
        RECT 490.425 2794.610 491.010 2794.620 ;
        RECT 495.230 2794.610 495.610 2794.620 ;
        RECT 496.405 2794.610 496.735 2794.625 ;
        RECT 490.425 2794.310 491.210 2794.610 ;
        RECT 495.230 2794.310 496.735 2794.610 ;
        RECT 490.425 2794.300 491.010 2794.310 ;
        RECT 495.230 2794.300 495.610 2794.310 ;
        RECT 490.425 2794.295 490.755 2794.300 ;
        RECT 496.405 2794.295 496.735 2794.310 ;
        RECT 497.785 2794.620 498.115 2794.625 ;
        RECT 497.785 2794.610 498.370 2794.620 ;
        RECT 500.750 2794.610 501.130 2794.620 ;
        RECT 501.925 2794.610 502.255 2794.625 ;
        RECT 497.785 2794.310 498.570 2794.610 ;
        RECT 500.750 2794.310 502.255 2794.610 ;
        RECT 497.785 2794.300 498.370 2794.310 ;
        RECT 500.750 2794.300 501.130 2794.310 ;
        RECT 497.785 2794.295 498.115 2794.300 ;
        RECT 501.925 2794.295 502.255 2794.310 ;
        RECT 507.190 2794.610 507.570 2794.620 ;
        RECT 510.205 2794.610 510.535 2794.625 ;
        RECT 507.190 2794.310 510.535 2794.610 ;
        RECT 507.190 2794.300 507.570 2794.310 ;
        RECT 510.205 2794.295 510.535 2794.310 ;
        RECT 516.390 2794.610 516.770 2794.620 ;
        RECT 517.105 2794.610 517.435 2794.625 ;
        RECT 524.005 2794.620 524.335 2794.625 ;
        RECT 523.750 2794.610 524.335 2794.620 ;
        RECT 516.390 2794.310 517.435 2794.610 ;
        RECT 523.550 2794.310 524.335 2794.610 ;
        RECT 516.390 2794.300 516.770 2794.310 ;
        RECT 517.105 2794.295 517.435 2794.310 ;
        RECT 523.750 2794.300 524.335 2794.310 ;
        RECT 526.510 2794.610 526.890 2794.620 ;
        RECT 527.685 2794.610 528.015 2794.625 ;
        RECT 526.510 2794.310 528.015 2794.610 ;
        RECT 526.510 2794.300 526.890 2794.310 ;
        RECT 524.005 2794.295 524.335 2794.300 ;
        RECT 527.685 2794.295 528.015 2794.310 ;
        RECT 530.190 2794.610 530.570 2794.620 ;
        RECT 530.905 2794.610 531.235 2794.625 ;
        RECT 530.190 2794.310 531.235 2794.610 ;
        RECT 530.190 2794.300 530.570 2794.310 ;
        RECT 530.905 2794.295 531.235 2794.310 ;
        RECT 535.710 2794.610 536.090 2794.620 ;
        RECT 537.345 2794.610 537.675 2794.625 ;
        RECT 542.405 2794.620 542.735 2794.625 ;
        RECT 542.150 2794.610 542.735 2794.620 ;
        RECT 535.710 2794.310 537.675 2794.610 ;
        RECT 541.950 2794.310 542.735 2794.610 ;
        RECT 535.710 2794.300 536.090 2794.310 ;
        RECT 537.345 2794.295 537.675 2794.310 ;
        RECT 542.150 2794.300 542.735 2794.310 ;
        RECT 547.670 2794.610 548.050 2794.620 ;
        RECT 551.605 2794.610 551.935 2794.625 ;
        RECT 547.670 2794.310 551.935 2794.610 ;
        RECT 547.670 2794.300 548.050 2794.310 ;
        RECT 542.405 2794.295 542.735 2794.300 ;
        RECT 551.605 2794.295 551.935 2794.310 ;
        RECT 979.865 2794.610 980.195 2794.625 ;
        RECT 980.990 2794.610 981.370 2794.620 ;
        RECT 979.865 2794.310 981.370 2794.610 ;
        RECT 979.865 2794.295 980.195 2794.310 ;
        RECT 980.990 2794.300 981.370 2794.310 ;
        RECT 986.765 2794.610 987.095 2794.625 ;
        RECT 987.430 2794.610 987.810 2794.620 ;
        RECT 986.765 2794.310 987.810 2794.610 ;
        RECT 986.765 2794.295 987.095 2794.310 ;
        RECT 987.430 2794.300 987.810 2794.310 ;
        RECT 1007.465 2794.610 1007.795 2794.625 ;
        RECT 1008.590 2794.610 1008.970 2794.620 ;
        RECT 1007.465 2794.310 1008.970 2794.610 ;
        RECT 1007.465 2794.295 1007.795 2794.310 ;
        RECT 1008.590 2794.300 1008.970 2794.310 ;
        RECT 1013.190 2794.610 1013.570 2794.620 ;
        RECT 1013.905 2794.610 1014.235 2794.625 ;
        RECT 1013.190 2794.310 1014.235 2794.610 ;
        RECT 1013.190 2794.300 1013.570 2794.310 ;
        RECT 1013.905 2794.295 1014.235 2794.310 ;
        RECT 1019.630 2794.610 1020.010 2794.620 ;
        RECT 1020.805 2794.610 1021.135 2794.625 ;
        RECT 1019.630 2794.310 1021.135 2794.610 ;
        RECT 1019.630 2794.300 1020.010 2794.310 ;
        RECT 1020.805 2794.295 1021.135 2794.310 ;
        RECT 1026.990 2794.610 1027.370 2794.620 ;
        RECT 1027.705 2794.610 1028.035 2794.625 ;
        RECT 1026.990 2794.310 1028.035 2794.610 ;
        RECT 1026.990 2794.300 1027.370 2794.310 ;
        RECT 1027.705 2794.295 1028.035 2794.310 ;
        RECT 1030.465 2794.620 1030.795 2794.625 ;
        RECT 1041.965 2794.620 1042.295 2794.625 ;
        RECT 1053.005 2794.620 1053.335 2794.625 ;
        RECT 1030.465 2794.610 1031.050 2794.620 ;
        RECT 1041.710 2794.610 1042.295 2794.620 ;
        RECT 1052.750 2794.610 1053.335 2794.620 ;
        RECT 1030.465 2794.310 1031.250 2794.610 ;
        RECT 1041.510 2794.310 1042.295 2794.610 ;
        RECT 1052.550 2794.310 1053.335 2794.610 ;
        RECT 1030.465 2794.300 1031.050 2794.310 ;
        RECT 1041.710 2794.300 1042.295 2794.310 ;
        RECT 1052.750 2794.300 1053.335 2794.310 ;
        RECT 1030.465 2794.295 1030.795 2794.300 ;
        RECT 1041.965 2794.295 1042.295 2794.300 ;
        RECT 1053.005 2794.295 1053.335 2794.300 ;
        RECT 1058.985 2794.620 1059.315 2794.625 ;
        RECT 1065.425 2794.620 1065.755 2794.625 ;
        RECT 1058.985 2794.610 1059.570 2794.620 ;
        RECT 1065.425 2794.610 1066.010 2794.620 ;
        RECT 1069.565 2794.610 1069.895 2794.625 ;
        RECT 1076.465 2794.620 1076.795 2794.625 ;
        RECT 1070.230 2794.610 1070.610 2794.620 ;
        RECT 1058.985 2794.310 1059.770 2794.610 ;
        RECT 1065.425 2794.310 1066.210 2794.610 ;
        RECT 1069.565 2794.310 1070.610 2794.610 ;
        RECT 1058.985 2794.300 1059.570 2794.310 ;
        RECT 1065.425 2794.300 1066.010 2794.310 ;
        RECT 1058.985 2794.295 1059.315 2794.300 ;
        RECT 1065.425 2794.295 1065.755 2794.300 ;
        RECT 1069.565 2794.295 1069.895 2794.310 ;
        RECT 1070.230 2794.300 1070.610 2794.310 ;
        RECT 1076.465 2794.610 1077.050 2794.620 ;
        RECT 1087.710 2794.610 1088.090 2794.620 ;
        RECT 1089.805 2794.610 1090.135 2794.625 ;
        RECT 1076.465 2794.310 1077.250 2794.610 ;
        RECT 1087.710 2794.310 1090.135 2794.610 ;
        RECT 1076.465 2794.300 1077.050 2794.310 ;
        RECT 1087.710 2794.300 1088.090 2794.310 ;
        RECT 1076.465 2794.295 1076.795 2794.300 ;
        RECT 1089.805 2794.295 1090.135 2794.310 ;
        RECT 1094.150 2794.610 1094.530 2794.620 ;
        RECT 1094.865 2794.610 1095.195 2794.625 ;
        RECT 1111.885 2794.620 1112.215 2794.625 ;
        RECT 1111.630 2794.610 1112.215 2794.620 ;
        RECT 1094.150 2794.310 1095.195 2794.610 ;
        RECT 1111.430 2794.310 1112.215 2794.610 ;
        RECT 1094.150 2794.300 1094.530 2794.310 ;
        RECT 1094.865 2794.295 1095.195 2794.310 ;
        RECT 1111.630 2794.300 1112.215 2794.310 ;
        RECT 1111.885 2794.295 1112.215 2794.300 ;
        RECT 1117.865 2794.620 1118.195 2794.625 ;
        RECT 1122.465 2794.620 1122.795 2794.625 ;
        RECT 1129.365 2794.620 1129.695 2794.625 ;
        RECT 1135.805 2794.620 1136.135 2794.625 ;
        RECT 1117.865 2794.610 1118.450 2794.620 ;
        RECT 1122.465 2794.610 1123.050 2794.620 ;
        RECT 1129.110 2794.610 1129.695 2794.620 ;
        RECT 1135.550 2794.610 1136.135 2794.620 ;
        RECT 1117.865 2794.310 1118.650 2794.610 ;
        RECT 1122.465 2794.310 1123.250 2794.610 ;
        RECT 1128.910 2794.310 1129.695 2794.610 ;
        RECT 1135.350 2794.310 1136.135 2794.610 ;
        RECT 1117.865 2794.300 1118.450 2794.310 ;
        RECT 1122.465 2794.300 1123.050 2794.310 ;
        RECT 1129.110 2794.300 1129.695 2794.310 ;
        RECT 1135.550 2794.300 1136.135 2794.310 ;
        RECT 1117.865 2794.295 1118.195 2794.300 ;
        RECT 1122.465 2794.295 1122.795 2794.300 ;
        RECT 1129.365 2794.295 1129.695 2794.300 ;
        RECT 1135.805 2794.295 1136.135 2794.300 ;
        RECT 1140.865 2794.620 1141.195 2794.625 ;
        RECT 1147.765 2794.620 1148.095 2794.625 ;
        RECT 1140.865 2794.610 1141.450 2794.620 ;
        RECT 1147.510 2794.610 1148.095 2794.620 ;
        RECT 1140.865 2794.310 1141.650 2794.610 ;
        RECT 1147.310 2794.310 1148.095 2794.610 ;
        RECT 1140.865 2794.300 1141.450 2794.310 ;
        RECT 1147.510 2794.300 1148.095 2794.310 ;
        RECT 1140.865 2794.295 1141.195 2794.300 ;
        RECT 1147.765 2794.295 1148.095 2794.300 ;
        RECT 1607.765 2794.610 1608.095 2794.625 ;
        RECT 1613.950 2794.610 1614.330 2794.620 ;
        RECT 1607.765 2794.310 1614.330 2794.610 ;
        RECT 1607.765 2794.295 1608.095 2794.310 ;
        RECT 1613.950 2794.300 1614.330 2794.310 ;
        RECT 1614.665 2794.610 1614.995 2794.625 ;
        RECT 1620.390 2794.610 1620.770 2794.620 ;
        RECT 1614.665 2794.310 1620.770 2794.610 ;
        RECT 1614.665 2794.295 1614.995 2794.310 ;
        RECT 1620.390 2794.300 1620.770 2794.310 ;
        RECT 1621.565 2794.610 1621.895 2794.625 ;
        RECT 1625.910 2794.610 1626.290 2794.620 ;
        RECT 1621.565 2794.310 1626.290 2794.610 ;
        RECT 1621.565 2794.295 1621.895 2794.310 ;
        RECT 1625.910 2794.300 1626.290 2794.310 ;
        RECT 1628.465 2794.610 1628.795 2794.625 ;
        RECT 1631.430 2794.610 1631.810 2794.620 ;
        RECT 1628.465 2794.310 1631.810 2794.610 ;
        RECT 1628.465 2794.295 1628.795 2794.310 ;
        RECT 1631.430 2794.300 1631.810 2794.310 ;
        RECT 1635.365 2794.610 1635.695 2794.625 ;
        RECT 1637.870 2794.610 1638.250 2794.620 ;
        RECT 1635.365 2794.310 1638.250 2794.610 ;
        RECT 1635.365 2794.295 1635.695 2794.310 ;
        RECT 1637.870 2794.300 1638.250 2794.310 ;
        RECT 1646.405 2794.610 1646.735 2794.625 ;
        RECT 1649.165 2794.620 1649.495 2794.625 ;
        RECT 1647.990 2794.610 1648.370 2794.620 ;
        RECT 1646.405 2794.310 1648.370 2794.610 ;
        RECT 1646.405 2794.295 1646.735 2794.310 ;
        RECT 1647.990 2794.300 1648.370 2794.310 ;
        RECT 1648.910 2794.610 1649.495 2794.620 ;
        RECT 1652.385 2794.620 1652.715 2794.625 ;
        RECT 1652.385 2794.610 1652.970 2794.620 ;
        RECT 1656.065 2794.610 1656.395 2794.625 ;
        RECT 1661.790 2794.610 1662.170 2794.620 ;
        RECT 1648.910 2794.310 1649.720 2794.610 ;
        RECT 1652.385 2794.310 1653.170 2794.610 ;
        RECT 1656.065 2794.310 1662.170 2794.610 ;
        RECT 1648.910 2794.300 1649.495 2794.310 ;
        RECT 1649.165 2794.295 1649.495 2794.300 ;
        RECT 1652.385 2794.300 1652.970 2794.310 ;
        RECT 1652.385 2794.295 1652.715 2794.300 ;
        RECT 1656.065 2794.295 1656.395 2794.310 ;
        RECT 1661.790 2794.300 1662.170 2794.310 ;
        RECT 1662.965 2794.610 1663.295 2794.625 ;
        RECT 1666.390 2794.610 1666.770 2794.620 ;
        RECT 1662.965 2794.310 1666.770 2794.610 ;
        RECT 1662.965 2794.295 1663.295 2794.310 ;
        RECT 1666.390 2794.300 1666.770 2794.310 ;
        RECT 1669.865 2794.610 1670.195 2794.625 ;
        RECT 1672.830 2794.610 1673.210 2794.620 ;
        RECT 1669.865 2794.310 1673.210 2794.610 ;
        RECT 1669.865 2794.295 1670.195 2794.310 ;
        RECT 1672.830 2794.300 1673.210 2794.310 ;
        RECT 1676.765 2794.610 1677.095 2794.625 ;
        RECT 1683.665 2794.620 1683.995 2794.625 ;
        RECT 1679.270 2794.610 1679.650 2794.620 ;
        RECT 1683.665 2794.610 1684.250 2794.620 ;
        RECT 1676.765 2794.310 1679.650 2794.610 ;
        RECT 1683.440 2794.310 1684.250 2794.610 ;
        RECT 1676.765 2794.295 1677.095 2794.310 ;
        RECT 1679.270 2794.300 1679.650 2794.310 ;
        RECT 1683.665 2794.300 1684.250 2794.310 ;
        RECT 1690.565 2794.610 1690.895 2794.625 ;
        RECT 1695.830 2794.610 1696.210 2794.620 ;
        RECT 1690.565 2794.310 1696.210 2794.610 ;
        RECT 1683.665 2794.295 1683.995 2794.300 ;
        RECT 1690.565 2794.295 1690.895 2794.310 ;
        RECT 1695.830 2794.300 1696.210 2794.310 ;
        RECT 1697.465 2794.610 1697.795 2794.625 ;
        RECT 1706.205 2794.620 1706.535 2794.625 ;
        RECT 1712.645 2794.620 1712.975 2794.625 ;
        RECT 1718.165 2794.620 1718.495 2794.625 ;
        RECT 1702.270 2794.610 1702.650 2794.620 ;
        RECT 1705.950 2794.610 1706.535 2794.620 ;
        RECT 1712.390 2794.610 1712.975 2794.620 ;
        RECT 1717.910 2794.610 1718.495 2794.620 ;
        RECT 1697.465 2794.310 1702.650 2794.610 ;
        RECT 1705.750 2794.310 1706.535 2794.610 ;
        RECT 1712.190 2794.310 1712.975 2794.610 ;
        RECT 1717.710 2794.310 1718.495 2794.610 ;
        RECT 1697.465 2794.295 1697.795 2794.310 ;
        RECT 1702.270 2794.300 1702.650 2794.310 ;
        RECT 1705.950 2794.300 1706.535 2794.310 ;
        RECT 1712.390 2794.300 1712.975 2794.310 ;
        RECT 1717.910 2794.300 1718.495 2794.310 ;
        RECT 1723.430 2794.610 1723.810 2794.620 ;
        RECT 1724.145 2794.610 1724.475 2794.625 ;
        RECT 1723.430 2794.310 1724.475 2794.610 ;
        RECT 1723.430 2794.300 1723.810 2794.310 ;
        RECT 1706.205 2794.295 1706.535 2794.300 ;
        RECT 1712.645 2794.295 1712.975 2794.300 ;
        RECT 1718.165 2794.295 1718.495 2794.300 ;
        RECT 1724.145 2794.295 1724.475 2794.310 ;
        RECT 1728.745 2794.620 1729.075 2794.625 ;
        RECT 1734.265 2794.620 1734.595 2794.625 ;
        RECT 1741.165 2794.620 1741.495 2794.625 ;
        RECT 1747.605 2794.620 1747.935 2794.625 ;
        RECT 1728.745 2794.610 1729.330 2794.620 ;
        RECT 1734.265 2794.610 1734.850 2794.620 ;
        RECT 1740.910 2794.610 1741.495 2794.620 ;
        RECT 1747.350 2794.610 1747.935 2794.620 ;
        RECT 1728.745 2794.310 1729.530 2794.610 ;
        RECT 1734.265 2794.310 1735.050 2794.610 ;
        RECT 1740.710 2794.310 1741.495 2794.610 ;
        RECT 1747.150 2794.310 1747.935 2794.610 ;
        RECT 1728.745 2794.300 1729.330 2794.310 ;
        RECT 1734.265 2794.300 1734.850 2794.310 ;
        RECT 1740.910 2794.300 1741.495 2794.310 ;
        RECT 1747.350 2794.300 1747.935 2794.310 ;
        RECT 1728.745 2794.295 1729.075 2794.300 ;
        RECT 1734.265 2794.295 1734.595 2794.300 ;
        RECT 1741.165 2794.295 1741.495 2794.300 ;
        RECT 1747.605 2794.295 1747.935 2794.300 ;
        RECT 1758.645 2794.610 1758.975 2794.625 ;
        RECT 1794.270 2794.610 1794.650 2794.620 ;
        RECT 1758.645 2794.310 1794.650 2794.610 ;
        RECT 1758.645 2794.295 1758.975 2794.310 ;
        RECT 1794.270 2794.300 1794.650 2794.310 ;
        RECT 1017.585 2793.930 1017.915 2793.945 ;
        RECT 1018.710 2793.930 1019.090 2793.940 ;
        RECT 1017.585 2793.630 1019.090 2793.930 ;
        RECT 1017.585 2793.615 1017.915 2793.630 ;
        RECT 1018.710 2793.620 1019.090 2793.630 ;
        RECT 1083.110 2793.930 1083.490 2793.940 ;
        RECT 1088.885 2793.930 1089.215 2793.945 ;
        RECT 1083.110 2793.630 1089.215 2793.930 ;
        RECT 1083.110 2793.620 1083.490 2793.630 ;
        RECT 1088.885 2793.615 1089.215 2793.630 ;
        RECT 1159.265 2793.930 1159.595 2793.945 ;
        RECT 1164.070 2793.930 1164.450 2793.940 ;
        RECT 1159.265 2793.630 1164.450 2793.930 ;
        RECT 1159.265 2793.615 1159.595 2793.630 ;
        RECT 1164.070 2793.620 1164.450 2793.630 ;
        RECT 1166.165 2793.930 1166.495 2793.945 ;
        RECT 1610.985 2793.940 1611.315 2793.945 ;
        RECT 1617.885 2793.940 1618.215 2793.945 ;
        RECT 1167.750 2793.930 1168.130 2793.940 ;
        RECT 1610.985 2793.930 1611.570 2793.940 ;
        RECT 1166.165 2793.630 1168.130 2793.930 ;
        RECT 1610.760 2793.630 1611.570 2793.930 ;
        RECT 1166.165 2793.615 1166.495 2793.630 ;
        RECT 1167.750 2793.620 1168.130 2793.630 ;
        RECT 1610.985 2793.620 1611.570 2793.630 ;
        RECT 1617.630 2793.930 1618.215 2793.940 ;
        RECT 1624.070 2793.930 1624.450 2793.940 ;
        RECT 1624.785 2793.930 1625.115 2793.945 ;
        RECT 1617.630 2793.630 1618.440 2793.930 ;
        RECT 1624.070 2793.630 1625.115 2793.930 ;
        RECT 1617.630 2793.620 1618.215 2793.630 ;
        RECT 1624.070 2793.620 1624.450 2793.630 ;
        RECT 1610.985 2793.615 1611.315 2793.620 ;
        RECT 1617.885 2793.615 1618.215 2793.620 ;
        RECT 1624.785 2793.615 1625.115 2793.630 ;
        RECT 1630.510 2793.930 1630.890 2793.940 ;
        RECT 1631.685 2793.930 1632.015 2793.945 ;
        RECT 1630.510 2793.630 1632.015 2793.930 ;
        RECT 1630.510 2793.620 1630.890 2793.630 ;
        RECT 1631.685 2793.615 1632.015 2793.630 ;
        RECT 1635.110 2793.930 1635.490 2793.940 ;
        RECT 1638.585 2793.930 1638.915 2793.945 ;
        RECT 1635.110 2793.630 1638.915 2793.930 ;
        RECT 1635.110 2793.620 1635.490 2793.630 ;
        RECT 1638.585 2793.615 1638.915 2793.630 ;
        RECT 1642.265 2793.615 1642.595 2793.945 ;
        RECT 1649.625 2793.930 1649.955 2793.945 ;
        RECT 1658.825 2793.940 1659.155 2793.945 ;
        RECT 1663.425 2793.940 1663.755 2793.945 ;
        RECT 1670.325 2793.940 1670.655 2793.945 ;
        RECT 1655.350 2793.930 1655.730 2793.940 ;
        RECT 1649.625 2793.630 1655.730 2793.930 ;
        RECT 1649.625 2793.615 1649.955 2793.630 ;
        RECT 1655.350 2793.620 1655.730 2793.630 ;
        RECT 1658.825 2793.930 1659.410 2793.940 ;
        RECT 1663.425 2793.930 1664.010 2793.940 ;
        RECT 1670.070 2793.930 1670.655 2793.940 ;
        RECT 1658.825 2793.630 1659.610 2793.930 ;
        RECT 1663.425 2793.630 1664.210 2793.930 ;
        RECT 1669.870 2793.630 1670.655 2793.930 ;
        RECT 1658.825 2793.620 1659.410 2793.630 ;
        RECT 1663.425 2793.620 1664.010 2793.630 ;
        RECT 1670.070 2793.620 1670.655 2793.630 ;
        RECT 1658.825 2793.615 1659.155 2793.620 ;
        RECT 1663.425 2793.615 1663.755 2793.620 ;
        RECT 1670.325 2793.615 1670.655 2793.620 ;
        RECT 1677.225 2793.940 1677.555 2793.945 ;
        RECT 1677.225 2793.930 1677.810 2793.940 ;
        RECT 1682.285 2793.930 1682.615 2793.945 ;
        RECT 1682.950 2793.930 1683.330 2793.940 ;
        RECT 1677.225 2793.630 1678.010 2793.930 ;
        RECT 1682.285 2793.630 1683.330 2793.930 ;
        RECT 1677.225 2793.620 1677.810 2793.630 ;
        RECT 1677.225 2793.615 1677.555 2793.620 ;
        RECT 1682.285 2793.615 1682.615 2793.630 ;
        RECT 1682.950 2793.620 1683.330 2793.630 ;
        RECT 1690.105 2793.615 1690.435 2793.945 ;
        RECT 1695.165 2793.940 1695.495 2793.945 ;
        RECT 1694.910 2793.930 1695.495 2793.940 ;
        RECT 1694.710 2793.630 1695.495 2793.930 ;
        RECT 1694.910 2793.620 1695.495 2793.630 ;
        RECT 1695.165 2793.615 1695.495 2793.620 ;
        RECT 1699.305 2793.940 1699.635 2793.945 ;
        RECT 1699.305 2793.930 1699.890 2793.940 ;
        RECT 1766.465 2793.930 1766.795 2793.945 ;
        RECT 1767.590 2793.930 1767.970 2793.940 ;
        RECT 1699.305 2793.630 1700.090 2793.930 ;
        RECT 1766.465 2793.630 1767.970 2793.930 ;
        RECT 1699.305 2793.620 1699.890 2793.630 ;
        RECT 1699.305 2793.615 1699.635 2793.620 ;
        RECT 1766.465 2793.615 1766.795 2793.630 ;
        RECT 1767.590 2793.620 1767.970 2793.630 ;
        RECT 1773.365 2793.930 1773.695 2793.945 ;
        RECT 1780.265 2793.940 1780.595 2793.945 ;
        RECT 1774.030 2793.930 1774.410 2793.940 ;
        RECT 1780.265 2793.930 1780.850 2793.940 ;
        RECT 1773.365 2793.630 1774.410 2793.930 ;
        RECT 1780.040 2793.630 1780.850 2793.930 ;
        RECT 1773.365 2793.615 1773.695 2793.630 ;
        RECT 1774.030 2793.620 1774.410 2793.630 ;
        RECT 1780.265 2793.620 1780.850 2793.630 ;
        RECT 1780.265 2793.615 1780.595 2793.620 ;
        RECT 348.950 2793.250 349.330 2793.260 ;
        RECT 351.045 2793.250 351.375 2793.265 ;
        RECT 348.950 2792.950 351.375 2793.250 ;
        RECT 348.950 2792.940 349.330 2792.950 ;
        RECT 351.045 2792.935 351.375 2792.950 ;
        RECT 396.790 2793.250 397.170 2793.260 ;
        RECT 397.965 2793.250 398.295 2793.265 ;
        RECT 396.790 2792.950 398.295 2793.250 ;
        RECT 396.790 2792.940 397.170 2792.950 ;
        RECT 397.965 2792.935 398.295 2792.950 ;
        RECT 414.065 2793.260 414.395 2793.265 ;
        RECT 414.065 2793.250 414.650 2793.260 ;
        RECT 426.025 2793.250 426.355 2793.265 ;
        RECT 427.150 2793.250 427.530 2793.260 ;
        RECT 414.065 2792.950 414.850 2793.250 ;
        RECT 426.025 2792.950 427.530 2793.250 ;
        RECT 414.065 2792.940 414.650 2792.950 ;
        RECT 414.065 2792.935 414.395 2792.940 ;
        RECT 426.025 2792.935 426.355 2792.950 ;
        RECT 427.150 2792.940 427.530 2792.950 ;
        RECT 430.830 2793.250 431.210 2793.260 ;
        RECT 433.845 2793.250 434.175 2793.265 ;
        RECT 430.830 2792.950 434.175 2793.250 ;
        RECT 430.830 2792.940 431.210 2792.950 ;
        RECT 433.845 2792.935 434.175 2792.950 ;
        RECT 455.465 2793.260 455.795 2793.265 ;
        RECT 466.505 2793.260 466.835 2793.265 ;
        RECT 468.805 2793.260 469.135 2793.265 ;
        RECT 455.465 2793.250 456.050 2793.260 ;
        RECT 466.505 2793.250 467.090 2793.260 ;
        RECT 468.550 2793.250 469.135 2793.260 ;
        RECT 455.465 2792.950 456.250 2793.250 ;
        RECT 466.505 2792.950 467.290 2793.250 ;
        RECT 468.350 2792.950 469.135 2793.250 ;
        RECT 455.465 2792.940 456.050 2792.950 ;
        RECT 466.505 2792.940 467.090 2792.950 ;
        RECT 468.550 2792.940 469.135 2792.950 ;
        RECT 455.465 2792.935 455.795 2792.940 ;
        RECT 466.505 2792.935 466.835 2792.940 ;
        RECT 468.805 2792.935 469.135 2792.940 ;
        RECT 500.085 2793.250 500.415 2793.265 ;
        RECT 509.745 2793.260 510.075 2793.265 ;
        RECT 513.885 2793.260 514.215 2793.265 ;
        RECT 501.670 2793.250 502.050 2793.260 ;
        RECT 500.085 2792.950 502.050 2793.250 ;
        RECT 500.085 2792.935 500.415 2792.950 ;
        RECT 501.670 2792.940 502.050 2792.950 ;
        RECT 509.745 2793.250 510.330 2793.260 ;
        RECT 513.630 2793.250 514.215 2793.260 ;
        RECT 519.405 2793.250 519.735 2793.265 ;
        RECT 520.070 2793.250 520.450 2793.260 ;
        RECT 509.745 2792.950 510.530 2793.250 ;
        RECT 513.630 2792.950 514.440 2793.250 ;
        RECT 519.405 2792.950 520.450 2793.250 ;
        RECT 509.745 2792.940 510.330 2792.950 ;
        RECT 513.630 2792.940 514.215 2792.950 ;
        RECT 509.745 2792.935 510.075 2792.940 ;
        RECT 513.885 2792.935 514.215 2792.940 ;
        RECT 519.405 2792.935 519.735 2792.950 ;
        RECT 520.070 2792.940 520.450 2792.950 ;
        RECT 531.110 2793.250 531.490 2793.260 ;
        RECT 534.585 2793.250 534.915 2793.265 ;
        RECT 538.725 2793.260 539.055 2793.265 ;
        RECT 538.470 2793.250 539.055 2793.260 ;
        RECT 531.110 2792.950 534.915 2793.250 ;
        RECT 538.270 2792.950 539.055 2793.250 ;
        RECT 531.110 2792.940 531.490 2792.950 ;
        RECT 534.585 2792.935 534.915 2792.950 ;
        RECT 538.470 2792.940 539.055 2792.950 ;
        RECT 538.725 2792.935 539.055 2792.940 ;
        RECT 541.485 2793.250 541.815 2793.265 ;
        RECT 543.070 2793.250 543.450 2793.260 ;
        RECT 541.485 2792.950 543.450 2793.250 ;
        RECT 541.485 2792.935 541.815 2792.950 ;
        RECT 543.070 2792.940 543.450 2792.950 ;
        RECT 1010.685 2793.250 1011.015 2793.265 ;
        RECT 1024.485 2793.260 1024.815 2793.265 ;
        RECT 1012.270 2793.250 1012.650 2793.260 ;
        RECT 1024.230 2793.250 1024.815 2793.260 ;
        RECT 1010.685 2792.950 1012.650 2793.250 ;
        RECT 1024.030 2792.950 1024.815 2793.250 ;
        RECT 1010.685 2792.935 1011.015 2792.950 ;
        RECT 1012.270 2792.940 1012.650 2792.950 ;
        RECT 1024.230 2792.940 1024.815 2792.950 ;
        RECT 1024.485 2792.935 1024.815 2792.940 ;
        RECT 1045.185 2793.250 1045.515 2793.265 ;
        RECT 1048.150 2793.250 1048.530 2793.260 ;
        RECT 1045.185 2792.950 1048.530 2793.250 ;
        RECT 1045.185 2792.935 1045.515 2792.950 ;
        RECT 1048.150 2792.940 1048.530 2792.950 ;
        RECT 1174.445 2793.250 1174.775 2793.265 ;
        RECT 1186.865 2793.260 1187.195 2793.265 ;
        RECT 1175.110 2793.250 1175.490 2793.260 ;
        RECT 1186.865 2793.250 1187.450 2793.260 ;
        RECT 1174.445 2792.950 1175.490 2793.250 ;
        RECT 1186.640 2792.950 1187.450 2793.250 ;
        RECT 1174.445 2792.935 1174.775 2792.950 ;
        RECT 1175.110 2792.940 1175.490 2792.950 ;
        RECT 1186.865 2792.940 1187.450 2792.950 ;
        RECT 1411.550 2793.250 1411.930 2793.260 ;
        RECT 1642.280 2793.250 1642.580 2793.615 ;
        RECT 1411.550 2792.950 1642.580 2793.250 ;
        RECT 1690.120 2793.250 1690.420 2793.615 ;
        RECT 1740.245 2793.250 1740.575 2793.265 ;
        RECT 1789.670 2793.250 1790.050 2793.260 ;
        RECT 1690.120 2792.950 1740.575 2793.250 ;
        RECT 1411.550 2792.940 1411.930 2792.950 ;
        RECT 1186.865 2792.935 1187.195 2792.940 ;
        RECT 1740.245 2792.935 1740.575 2792.950 ;
        RECT 1761.190 2792.950 1790.050 2793.250 ;
        RECT 1159.725 2792.570 1160.055 2792.585 ;
        RECT 1193.765 2792.580 1194.095 2792.585 ;
        RECT 1180.630 2792.570 1181.010 2792.580 ;
        RECT 1159.725 2792.270 1181.010 2792.570 ;
        RECT 1159.725 2792.255 1160.055 2792.270 ;
        RECT 1180.630 2792.260 1181.010 2792.270 ;
        RECT 1193.510 2792.570 1194.095 2792.580 ;
        RECT 1417.070 2792.570 1417.450 2792.580 ;
        RECT 1642.265 2792.570 1642.595 2792.585 ;
        RECT 1193.510 2792.270 1194.320 2792.570 ;
        RECT 1417.070 2792.270 1642.595 2792.570 ;
        RECT 1193.510 2792.260 1194.095 2792.270 ;
        RECT 1417.070 2792.260 1417.450 2792.270 ;
        RECT 1193.765 2792.255 1194.095 2792.260 ;
        RECT 1642.265 2792.255 1642.595 2792.270 ;
        RECT 1690.105 2792.570 1690.435 2792.585 ;
        RECT 1728.285 2792.570 1728.615 2792.585 ;
        RECT 1690.105 2792.270 1728.615 2792.570 ;
        RECT 1690.105 2792.255 1690.435 2792.270 ;
        RECT 1728.285 2792.255 1728.615 2792.270 ;
        RECT 1752.665 2792.580 1752.995 2792.585 ;
        RECT 1752.665 2792.570 1753.250 2792.580 ;
        RECT 1761.190 2792.570 1761.490 2792.950 ;
        RECT 1789.670 2792.940 1790.050 2792.950 ;
        RECT 1752.665 2792.270 1753.450 2792.570 ;
        RECT 1758.430 2792.270 1761.490 2792.570 ;
        RECT 1787.165 2792.570 1787.495 2792.585 ;
        RECT 1787.830 2792.570 1788.210 2792.580 ;
        RECT 1787.165 2792.270 1788.210 2792.570 ;
        RECT 1752.665 2792.260 1753.250 2792.270 ;
        RECT 1752.665 2792.255 1752.995 2792.260 ;
        RECT 390.350 2791.890 390.730 2791.900 ;
        RECT 392.905 2791.890 393.235 2791.905 ;
        RECT 390.350 2791.590 393.235 2791.890 ;
        RECT 390.350 2791.580 390.730 2791.590 ;
        RECT 392.905 2791.575 393.235 2791.590 ;
        RECT 460.270 2791.890 460.650 2791.900 ;
        RECT 461.905 2791.890 462.235 2791.905 ;
        RECT 460.270 2791.590 462.235 2791.890 ;
        RECT 460.270 2791.580 460.650 2791.590 ;
        RECT 461.905 2791.575 462.235 2791.590 ;
        RECT 489.965 2791.890 490.295 2791.905 ;
        RECT 506.985 2791.890 507.315 2791.905 ;
        RECT 508.110 2791.890 508.490 2791.900 ;
        RECT 489.965 2791.590 508.490 2791.890 ;
        RECT 489.965 2791.575 490.295 2791.590 ;
        RECT 506.985 2791.575 507.315 2791.590 ;
        RECT 508.110 2791.580 508.490 2791.590 ;
        RECT 1075.545 2791.890 1075.875 2791.905 ;
        RECT 1105.190 2791.890 1105.570 2791.900 ;
        RECT 1107.745 2791.890 1108.075 2791.905 ;
        RECT 1075.545 2791.590 1108.075 2791.890 ;
        RECT 1075.545 2791.575 1075.875 2791.590 ;
        RECT 1105.190 2791.580 1105.570 2791.590 ;
        RECT 1107.745 2791.575 1108.075 2791.590 ;
        RECT 1152.365 2791.890 1152.695 2791.905 ;
        RECT 1159.265 2791.900 1159.595 2791.905 ;
        RECT 1153.030 2791.890 1153.410 2791.900 ;
        RECT 1159.265 2791.890 1159.850 2791.900 ;
        RECT 1152.365 2791.590 1153.410 2791.890 ;
        RECT 1159.040 2791.590 1159.850 2791.890 ;
        RECT 1152.365 2791.575 1152.695 2791.590 ;
        RECT 1153.030 2791.580 1153.410 2791.590 ;
        RECT 1159.265 2791.580 1159.850 2791.590 ;
        RECT 1418.910 2791.890 1419.290 2791.900 ;
        RECT 1758.430 2791.890 1758.730 2792.270 ;
        RECT 1787.165 2792.255 1787.495 2792.270 ;
        RECT 1787.830 2792.260 1788.210 2792.270 ;
        RECT 1418.910 2791.590 1758.730 2791.890 ;
        RECT 1418.910 2791.580 1419.290 2791.590 ;
        RECT 1159.265 2791.575 1159.595 2791.580 ;
        RECT 378.390 2791.210 378.770 2791.220 ;
        RECT 379.105 2791.210 379.435 2791.225 ;
        RECT 378.390 2790.910 379.435 2791.210 ;
        RECT 378.390 2790.900 378.770 2790.910 ;
        RECT 379.105 2790.895 379.435 2790.910 ;
        RECT 1417.990 2791.210 1418.370 2791.220 ;
        RECT 1758.645 2791.210 1758.975 2791.225 ;
        RECT 1417.990 2790.910 1758.975 2791.210 ;
        RECT 1417.990 2790.900 1418.370 2790.910 ;
        RECT 1758.645 2790.895 1758.975 2790.910 ;
        RECT 1759.565 2791.210 1759.895 2791.225 ;
        RECT 1762.070 2791.210 1762.450 2791.220 ;
        RECT 1759.565 2790.910 1762.450 2791.210 ;
        RECT 1759.565 2790.895 1759.895 2790.910 ;
        RECT 1762.070 2790.900 1762.450 2790.910 ;
        RECT 1773.365 2791.210 1773.695 2791.225 ;
        RECT 1778.630 2791.210 1779.010 2791.220 ;
        RECT 1773.365 2790.910 1779.010 2791.210 ;
        RECT 1773.365 2790.895 1773.695 2790.910 ;
        RECT 1778.630 2790.900 1779.010 2790.910 ;
        RECT 1728.285 2790.530 1728.615 2790.545 ;
        RECT 1759.565 2790.530 1759.895 2790.545 ;
        RECT 1765.750 2790.530 1766.130 2790.540 ;
        RECT 1728.285 2790.230 1758.730 2790.530 ;
        RECT 1728.285 2790.215 1728.615 2790.230 ;
        RECT 1587.065 2789.860 1587.395 2789.865 ;
        RECT 1587.065 2789.850 1587.650 2789.860 ;
        RECT 1586.840 2789.550 1587.650 2789.850 ;
        RECT 1587.065 2789.540 1587.650 2789.550 ;
        RECT 1600.865 2789.850 1601.195 2789.865 ;
        RECT 1602.910 2789.850 1603.290 2789.860 ;
        RECT 1600.865 2789.550 1603.290 2789.850 ;
        RECT 1587.065 2789.535 1587.395 2789.540 ;
        RECT 1600.865 2789.535 1601.195 2789.550 ;
        RECT 1602.910 2789.540 1603.290 2789.550 ;
        RECT 1684.125 2789.850 1684.455 2789.865 ;
        RECT 1689.390 2789.850 1689.770 2789.860 ;
        RECT 1684.125 2789.550 1689.770 2789.850 ;
        RECT 1684.125 2789.535 1684.455 2789.550 ;
        RECT 1689.390 2789.540 1689.770 2789.550 ;
        RECT 1001.025 2789.180 1001.355 2789.185 ;
        RECT 1001.025 2789.170 1001.610 2789.180 ;
        RECT 1000.800 2788.870 1001.610 2789.170 ;
        RECT 1001.025 2788.860 1001.610 2788.870 ;
        RECT 1001.025 2788.855 1001.355 2788.860 ;
        RECT 993.665 2788.500 993.995 2788.505 ;
        RECT 993.665 2788.490 994.250 2788.500 ;
        RECT 993.440 2788.190 994.250 2788.490 ;
        RECT 993.665 2788.180 994.250 2788.190 ;
        RECT 1035.270 2788.490 1035.650 2788.500 ;
        RECT 1038.285 2788.490 1038.615 2788.505 ;
        RECT 1035.270 2788.190 1038.615 2788.490 ;
        RECT 1035.270 2788.180 1035.650 2788.190 ;
        RECT 993.665 2788.175 993.995 2788.180 ;
        RECT 1038.285 2788.175 1038.615 2788.190 ;
        RECT 1051.830 2788.490 1052.210 2788.500 ;
        RECT 1055.305 2788.490 1055.635 2788.505 ;
        RECT 1051.830 2788.190 1055.635 2788.490 ;
        RECT 1051.830 2788.180 1052.210 2788.190 ;
        RECT 1055.305 2788.175 1055.635 2788.190 ;
        RECT 1086.790 2788.490 1087.170 2788.500 ;
        RECT 1089.345 2788.490 1089.675 2788.505 ;
        RECT 1086.790 2788.190 1089.675 2788.490 ;
        RECT 1086.790 2788.180 1087.170 2788.190 ;
        RECT 1089.345 2788.175 1089.675 2788.190 ;
        RECT 1128.190 2788.490 1128.570 2788.500 ;
        RECT 1130.745 2788.490 1131.075 2788.505 ;
        RECT 1128.190 2788.190 1131.075 2788.490 ;
        RECT 1128.190 2788.180 1128.570 2788.190 ;
        RECT 1130.745 2788.175 1131.075 2788.190 ;
        RECT 1163.150 2788.490 1163.530 2788.500 ;
        RECT 1165.705 2788.490 1166.035 2788.505 ;
        RECT 1163.150 2788.190 1166.035 2788.490 ;
        RECT 1163.150 2788.180 1163.530 2788.190 ;
        RECT 1165.705 2788.175 1166.035 2788.190 ;
        RECT 1718.625 2788.490 1718.955 2788.505 ;
        RECT 1724.350 2788.490 1724.730 2788.500 ;
        RECT 1718.625 2788.190 1724.730 2788.490 ;
        RECT 1758.430 2788.490 1758.730 2790.230 ;
        RECT 1759.565 2790.230 1766.130 2790.530 ;
        RECT 1759.565 2790.215 1759.895 2790.230 ;
        RECT 1765.750 2790.220 1766.130 2790.230 ;
        RECT 1766.465 2789.850 1766.795 2789.865 ;
        RECT 1772.190 2789.850 1772.570 2789.860 ;
        RECT 1766.465 2789.550 1772.570 2789.850 ;
        RECT 1766.465 2789.535 1766.795 2789.550 ;
        RECT 1772.190 2789.540 1772.570 2789.550 ;
        RECT 1783.230 2788.490 1783.610 2788.500 ;
        RECT 1758.430 2788.190 1783.610 2788.490 ;
        RECT 1718.625 2788.175 1718.955 2788.190 ;
        RECT 1724.350 2788.180 1724.730 2788.190 ;
        RECT 1783.230 2788.180 1783.610 2788.190 ;
        RECT 1034.605 2787.820 1034.935 2787.825 ;
        RECT 1034.350 2787.810 1034.935 2787.820 ;
        RECT 1039.870 2787.810 1040.250 2787.820 ;
        RECT 1041.505 2787.810 1041.835 2787.825 ;
        RECT 1034.350 2787.510 1035.160 2787.810 ;
        RECT 1039.870 2787.510 1041.835 2787.810 ;
        RECT 1034.350 2787.500 1034.935 2787.510 ;
        RECT 1039.870 2787.500 1040.250 2787.510 ;
        RECT 1034.605 2787.495 1034.935 2787.500 ;
        RECT 1041.505 2787.495 1041.835 2787.510 ;
        RECT 1046.310 2787.810 1046.690 2787.820 ;
        RECT 1048.405 2787.810 1048.735 2787.825 ;
        RECT 1062.205 2787.820 1062.535 2787.825 ;
        RECT 1046.310 2787.510 1048.735 2787.810 ;
        RECT 1046.310 2787.500 1046.690 2787.510 ;
        RECT 1048.405 2787.495 1048.735 2787.510 ;
        RECT 1061.950 2787.810 1062.535 2787.820 ;
        RECT 1067.470 2787.810 1067.850 2787.820 ;
        RECT 1069.105 2787.810 1069.435 2787.825 ;
        RECT 1061.950 2787.510 1062.760 2787.810 ;
        RECT 1067.470 2787.510 1069.435 2787.810 ;
        RECT 1061.950 2787.500 1062.535 2787.510 ;
        RECT 1067.470 2787.500 1067.850 2787.510 ;
        RECT 1062.205 2787.495 1062.535 2787.500 ;
        RECT 1069.105 2787.495 1069.435 2787.510 ;
        RECT 1073.910 2787.810 1074.290 2787.820 ;
        RECT 1076.005 2787.810 1076.335 2787.825 ;
        RECT 1073.910 2787.510 1076.335 2787.810 ;
        RECT 1073.910 2787.500 1074.290 2787.510 ;
        RECT 1076.005 2787.495 1076.335 2787.510 ;
        RECT 1081.270 2787.810 1081.650 2787.820 ;
        RECT 1082.905 2787.810 1083.235 2787.825 ;
        RECT 1089.805 2787.820 1090.135 2787.825 ;
        RECT 1081.270 2787.510 1083.235 2787.810 ;
        RECT 1081.270 2787.500 1081.650 2787.510 ;
        RECT 1082.905 2787.495 1083.235 2787.510 ;
        RECT 1089.550 2787.810 1090.135 2787.820 ;
        RECT 1095.990 2787.810 1096.370 2787.820 ;
        RECT 1096.705 2787.810 1097.035 2787.825 ;
        RECT 1103.605 2787.820 1103.935 2787.825 ;
        RECT 1089.550 2787.510 1090.360 2787.810 ;
        RECT 1095.990 2787.510 1097.035 2787.810 ;
        RECT 1089.550 2787.500 1090.135 2787.510 ;
        RECT 1095.990 2787.500 1096.370 2787.510 ;
        RECT 1089.805 2787.495 1090.135 2787.500 ;
        RECT 1096.705 2787.495 1097.035 2787.510 ;
        RECT 1103.350 2787.810 1103.935 2787.820 ;
        RECT 1109.790 2787.810 1110.170 2787.820 ;
        RECT 1110.505 2787.810 1110.835 2787.825 ;
        RECT 1103.350 2787.510 1104.160 2787.810 ;
        RECT 1109.790 2787.510 1110.835 2787.810 ;
        RECT 1103.350 2787.500 1103.935 2787.510 ;
        RECT 1109.790 2787.500 1110.170 2787.510 ;
        RECT 1103.605 2787.495 1103.935 2787.500 ;
        RECT 1110.505 2787.495 1110.835 2787.510 ;
        RECT 1116.230 2787.810 1116.610 2787.820 ;
        RECT 1117.405 2787.810 1117.735 2787.825 ;
        RECT 1116.230 2787.510 1117.735 2787.810 ;
        RECT 1116.230 2787.500 1116.610 2787.510 ;
        RECT 1117.405 2787.495 1117.735 2787.510 ;
        RECT 1121.750 2787.810 1122.130 2787.820 ;
        RECT 1124.305 2787.810 1124.635 2787.825 ;
        RECT 1131.205 2787.820 1131.535 2787.825 ;
        RECT 1121.750 2787.510 1124.635 2787.810 ;
        RECT 1121.750 2787.500 1122.130 2787.510 ;
        RECT 1124.305 2787.495 1124.635 2787.510 ;
        RECT 1130.950 2787.810 1131.535 2787.820 ;
        RECT 1137.390 2787.810 1137.770 2787.820 ;
        RECT 1138.105 2787.810 1138.435 2787.825 ;
        RECT 1130.950 2787.510 1131.760 2787.810 ;
        RECT 1137.390 2787.510 1138.435 2787.810 ;
        RECT 1130.950 2787.500 1131.535 2787.510 ;
        RECT 1137.390 2787.500 1137.770 2787.510 ;
        RECT 1131.205 2787.495 1131.535 2787.500 ;
        RECT 1138.105 2787.495 1138.435 2787.510 ;
        RECT 1143.830 2787.810 1144.210 2787.820 ;
        RECT 1145.005 2787.810 1145.335 2787.825 ;
        RECT 1143.830 2787.510 1145.335 2787.810 ;
        RECT 1143.830 2787.500 1144.210 2787.510 ;
        RECT 1145.005 2787.495 1145.335 2787.510 ;
        RECT 1151.190 2787.810 1151.570 2787.820 ;
        RECT 1151.905 2787.810 1152.235 2787.825 ;
        RECT 1151.190 2787.510 1152.235 2787.810 ;
        RECT 1151.190 2787.500 1151.570 2787.510 ;
        RECT 1151.905 2787.495 1152.235 2787.510 ;
        RECT 1153.950 2787.810 1154.330 2787.820 ;
        RECT 1158.805 2787.810 1159.135 2787.825 ;
        RECT 1165.245 2787.820 1165.575 2787.825 ;
        RECT 1172.605 2787.820 1172.935 2787.825 ;
        RECT 1153.950 2787.510 1159.135 2787.810 ;
        RECT 1153.950 2787.500 1154.330 2787.510 ;
        RECT 1158.805 2787.495 1159.135 2787.510 ;
        RECT 1164.990 2787.810 1165.575 2787.820 ;
        RECT 1172.350 2787.810 1172.935 2787.820 ;
        RECT 1164.990 2787.510 1165.800 2787.810 ;
        RECT 1172.150 2787.510 1172.935 2787.810 ;
        RECT 1164.990 2787.500 1165.575 2787.510 ;
        RECT 1172.350 2787.500 1172.935 2787.510 ;
        RECT 1178.790 2787.810 1179.170 2787.820 ;
        RECT 1179.505 2787.810 1179.835 2787.825 ;
        RECT 1186.405 2787.820 1186.735 2787.825 ;
        RECT 1178.790 2787.510 1179.835 2787.810 ;
        RECT 1178.790 2787.500 1179.170 2787.510 ;
        RECT 1165.245 2787.495 1165.575 2787.500 ;
        RECT 1172.605 2787.495 1172.935 2787.500 ;
        RECT 1179.505 2787.495 1179.835 2787.510 ;
        RECT 1186.150 2787.810 1186.735 2787.820 ;
        RECT 1191.670 2787.810 1192.050 2787.820 ;
        RECT 1193.305 2787.810 1193.635 2787.825 ;
        RECT 1186.150 2787.510 1186.960 2787.810 ;
        RECT 1191.670 2787.510 1193.635 2787.810 ;
        RECT 1186.150 2787.500 1186.735 2787.510 ;
        RECT 1191.670 2787.500 1192.050 2787.510 ;
        RECT 1186.405 2787.495 1186.735 2787.500 ;
        RECT 1193.305 2787.495 1193.635 2787.510 ;
        RECT 1198.110 2787.810 1198.490 2787.820 ;
        RECT 1200.205 2787.810 1200.535 2787.825 ;
        RECT 1198.110 2787.510 1200.535 2787.810 ;
        RECT 1198.110 2787.500 1198.490 2787.510 ;
        RECT 1200.205 2787.495 1200.535 2787.510 ;
        RECT 1580.165 2787.810 1580.495 2787.825 ;
        RECT 1581.750 2787.810 1582.130 2787.820 ;
        RECT 1580.165 2787.510 1582.130 2787.810 ;
        RECT 1580.165 2787.495 1580.495 2787.510 ;
        RECT 1581.750 2787.500 1582.130 2787.510 ;
        RECT 1593.965 2787.810 1594.295 2787.825 ;
        RECT 1594.630 2787.810 1595.010 2787.820 ;
        RECT 1593.965 2787.510 1595.010 2787.810 ;
        RECT 1593.965 2787.495 1594.295 2787.510 ;
        RECT 1594.630 2787.500 1595.010 2787.510 ;
        RECT 1601.325 2787.810 1601.655 2787.825 ;
        RECT 1604.750 2787.810 1605.130 2787.820 ;
        RECT 1601.325 2787.510 1605.130 2787.810 ;
        RECT 1601.325 2787.495 1601.655 2787.510 ;
        RECT 1604.750 2787.500 1605.130 2787.510 ;
        RECT 1704.365 2787.810 1704.695 2787.825 ;
        RECT 1708.710 2787.810 1709.090 2787.820 ;
        RECT 1704.365 2787.510 1709.090 2787.810 ;
        RECT 1704.365 2787.495 1704.695 2787.510 ;
        RECT 1708.710 2787.500 1709.090 2787.510 ;
        RECT 1711.265 2787.810 1711.595 2787.825 ;
        RECT 1713.310 2787.810 1713.690 2787.820 ;
        RECT 1711.265 2787.510 1713.690 2787.810 ;
        RECT 1711.265 2787.495 1711.595 2787.510 ;
        RECT 1713.310 2787.500 1713.690 2787.510 ;
        RECT 1718.165 2787.810 1718.495 2787.825 ;
        RECT 1719.750 2787.810 1720.130 2787.820 ;
        RECT 1718.165 2787.510 1720.130 2787.810 ;
        RECT 1718.165 2787.495 1718.495 2787.510 ;
        RECT 1719.750 2787.500 1720.130 2787.510 ;
        RECT 1725.065 2787.810 1725.395 2787.825 ;
        RECT 1730.790 2787.810 1731.170 2787.820 ;
        RECT 1725.065 2787.510 1731.170 2787.810 ;
        RECT 1725.065 2787.495 1725.395 2787.510 ;
        RECT 1730.790 2787.500 1731.170 2787.510 ;
        RECT 1731.965 2787.810 1732.295 2787.825 ;
        RECT 1737.230 2787.810 1737.610 2787.820 ;
        RECT 1731.965 2787.510 1737.610 2787.810 ;
        RECT 1731.965 2787.495 1732.295 2787.510 ;
        RECT 1737.230 2787.500 1737.610 2787.510 ;
        RECT 1738.865 2787.810 1739.195 2787.825 ;
        RECT 1743.670 2787.810 1744.050 2787.820 ;
        RECT 1738.865 2787.510 1744.050 2787.810 ;
        RECT 1738.865 2787.495 1739.195 2787.510 ;
        RECT 1743.670 2787.500 1744.050 2787.510 ;
        RECT 1745.765 2787.810 1746.095 2787.825 ;
        RECT 1748.270 2787.810 1748.650 2787.820 ;
        RECT 1745.765 2787.510 1748.650 2787.810 ;
        RECT 1745.765 2787.495 1746.095 2787.510 ;
        RECT 1748.270 2787.500 1748.650 2787.510 ;
        RECT 1753.125 2787.810 1753.455 2787.825 ;
        RECT 1754.710 2787.810 1755.090 2787.820 ;
        RECT 1753.125 2787.510 1755.090 2787.810 ;
        RECT 1753.125 2787.495 1753.455 2787.510 ;
        RECT 1754.710 2787.500 1755.090 2787.510 ;
        RECT 1642.265 2785.770 1642.595 2785.785 ;
        RECT 1644.310 2785.770 1644.690 2785.780 ;
        RECT 1642.265 2785.470 1644.690 2785.770 ;
        RECT 1642.265 2785.455 1642.595 2785.470 ;
        RECT 1644.310 2785.460 1644.690 2785.470 ;
        RECT 460.525 2723.890 460.855 2723.905 ;
        RECT 942.605 2723.890 942.935 2723.905 ;
        RECT 460.525 2723.590 942.935 2723.890 ;
        RECT 460.525 2723.575 460.855 2723.590 ;
        RECT 942.605 2723.575 942.935 2723.590 ;
        RECT 439.825 2723.210 440.155 2723.225 ;
        RECT 943.525 2723.210 943.855 2723.225 ;
        RECT 439.825 2722.910 943.855 2723.210 ;
        RECT 439.825 2722.895 440.155 2722.910 ;
        RECT 943.525 2722.895 943.855 2722.910 ;
        RECT 429.245 2722.530 429.575 2722.545 ;
        RECT 944.445 2722.530 944.775 2722.545 ;
        RECT 429.245 2722.230 944.775 2722.530 ;
        RECT 429.245 2722.215 429.575 2722.230 ;
        RECT 944.445 2722.215 944.775 2722.230 ;
        RECT 419.125 2721.850 419.455 2721.865 ;
        RECT 941.225 2721.850 941.555 2721.865 ;
        RECT 419.125 2721.550 941.555 2721.850 ;
        RECT 419.125 2721.535 419.455 2721.550 ;
        RECT 941.225 2721.535 941.555 2721.550 ;
        RECT 707.545 2716.410 707.875 2716.425 ;
        RECT 1041.505 2716.410 1041.835 2716.425 ;
        RECT 707.545 2716.110 1041.835 2716.410 ;
        RECT 707.545 2716.095 707.875 2716.110 ;
        RECT 1041.505 2716.095 1041.835 2716.110 ;
        RECT 720.885 2715.730 721.215 2715.745 ;
        RECT 1052.085 2715.730 1052.415 2715.745 ;
        RECT 720.885 2715.430 1052.415 2715.730 ;
        RECT 720.885 2715.415 721.215 2715.430 ;
        RECT 1052.085 2715.415 1052.415 2715.430 ;
        RECT 530.905 2715.050 531.235 2715.065 ;
        RECT 1030.925 2715.050 1031.255 2715.065 ;
        RECT 530.905 2714.750 1031.255 2715.050 ;
        RECT 530.905 2714.735 531.235 2714.750 ;
        RECT 1030.925 2714.735 1031.255 2714.750 ;
      LAYER met3 ;
        RECT 300.065 2696.480 1395.600 2697.340 ;
      LAYER met3 ;
        RECT 1396.000 2696.880 1400.000 2697.480 ;
      LAYER met3 ;
        RECT 300.065 2695.840 1396.000 2696.480 ;
        RECT 304.400 2694.440 1396.000 2695.840 ;
        RECT 300.065 2693.120 1396.000 2694.440 ;
        RECT 300.065 2691.720 1395.600 2693.120 ;
      LAYER met3 ;
        RECT 1396.000 2692.120 1400.000 2692.720 ;
      LAYER met3 ;
        RECT 300.065 2687.680 1396.000 2691.720 ;
        RECT 300.065 2686.320 1395.600 2687.680 ;
      LAYER met3 ;
        RECT 1396.000 2686.680 1400.000 2687.280 ;
      LAYER met3 ;
        RECT 304.400 2686.280 1395.600 2686.320 ;
        RECT 304.400 2684.920 1396.000 2686.280 ;
        RECT 300.065 2682.920 1396.000 2684.920 ;
        RECT 300.065 2681.520 1395.600 2682.920 ;
      LAYER met3 ;
        RECT 1396.000 2681.920 1400.000 2682.520 ;
      LAYER met3 ;
        RECT 300.065 2677.480 1396.000 2681.520 ;
        RECT 300.065 2676.800 1395.600 2677.480 ;
        RECT 304.400 2676.080 1395.600 2676.800 ;
      LAYER met3 ;
        RECT 1396.000 2676.480 1400.000 2677.080 ;
      LAYER met3 ;
        RECT 304.400 2675.400 1396.000 2676.080 ;
        RECT 300.065 2672.720 1396.000 2675.400 ;
        RECT 300.065 2671.320 1395.600 2672.720 ;
      LAYER met3 ;
        RECT 1396.000 2671.720 1400.000 2672.320 ;
      LAYER met3 ;
        RECT 300.065 2667.960 1396.000 2671.320 ;
        RECT 300.065 2667.280 1395.600 2667.960 ;
        RECT 304.400 2666.560 1395.600 2667.280 ;
      LAYER met3 ;
        RECT 1396.000 2666.960 1400.000 2667.560 ;
      LAYER met3 ;
        RECT 304.400 2665.880 1396.000 2666.560 ;
        RECT 300.065 2662.520 1396.000 2665.880 ;
        RECT 300.065 2661.120 1395.600 2662.520 ;
      LAYER met3 ;
        RECT 1396.000 2661.520 1400.000 2662.120 ;
      LAYER met3 ;
        RECT 300.065 2657.760 1396.000 2661.120 ;
        RECT 304.400 2656.360 1395.600 2657.760 ;
      LAYER met3 ;
        RECT 1396.000 2656.760 1400.000 2657.360 ;
      LAYER met3 ;
        RECT 300.065 2652.320 1396.000 2656.360 ;
        RECT 300.065 2650.920 1395.600 2652.320 ;
      LAYER met3 ;
        RECT 1396.000 2651.320 1400.000 2651.920 ;
      LAYER met3 ;
        RECT 300.065 2647.560 1396.000 2650.920 ;
        RECT 304.400 2646.160 1395.600 2647.560 ;
      LAYER met3 ;
        RECT 1396.000 2646.560 1400.000 2647.160 ;
      LAYER met3 ;
        RECT 300.065 2642.120 1396.000 2646.160 ;
        RECT 300.065 2640.720 1395.600 2642.120 ;
      LAYER met3 ;
        RECT 1396.000 2641.120 1400.000 2641.720 ;
      LAYER met3 ;
        RECT 300.065 2638.040 1396.000 2640.720 ;
        RECT 304.400 2637.360 1396.000 2638.040 ;
        RECT 304.400 2636.640 1395.600 2637.360 ;
        RECT 300.065 2635.960 1395.600 2636.640 ;
      LAYER met3 ;
        RECT 1396.000 2636.360 1400.000 2636.960 ;
      LAYER met3 ;
        RECT 300.065 2632.600 1396.000 2635.960 ;
        RECT 300.065 2631.200 1395.600 2632.600 ;
      LAYER met3 ;
        RECT 1396.000 2631.600 1400.000 2632.200 ;
      LAYER met3 ;
        RECT 300.065 2628.520 1396.000 2631.200 ;
        RECT 304.400 2627.160 1396.000 2628.520 ;
        RECT 304.400 2627.120 1395.600 2627.160 ;
        RECT 300.065 2625.760 1395.600 2627.120 ;
      LAYER met3 ;
        RECT 1396.000 2626.160 1400.000 2626.760 ;
      LAYER met3 ;
        RECT 300.065 2622.400 1396.000 2625.760 ;
        RECT 300.065 2621.000 1395.600 2622.400 ;
      LAYER met3 ;
        RECT 1396.000 2621.400 1400.000 2622.000 ;
      LAYER met3 ;
        RECT 300.065 2619.000 1396.000 2621.000 ;
        RECT 304.400 2617.600 1396.000 2619.000 ;
        RECT 300.065 2616.960 1396.000 2617.600 ;
        RECT 300.065 2615.560 1395.600 2616.960 ;
      LAYER met3 ;
        RECT 1396.000 2615.960 1400.000 2616.560 ;
      LAYER met3 ;
        RECT 300.065 2612.200 1396.000 2615.560 ;
        RECT 300.065 2610.800 1395.600 2612.200 ;
      LAYER met3 ;
        RECT 1396.000 2611.200 1400.000 2611.800 ;
      LAYER met3 ;
        RECT 300.065 2609.480 1396.000 2610.800 ;
        RECT 304.400 2608.080 1396.000 2609.480 ;
        RECT 300.065 2606.760 1396.000 2608.080 ;
        RECT 300.065 2605.360 1395.600 2606.760 ;
      LAYER met3 ;
        RECT 1396.000 2605.760 1400.000 2606.360 ;
      LAYER met3 ;
        RECT 300.065 2602.000 1396.000 2605.360 ;
        RECT 300.065 2600.600 1395.600 2602.000 ;
      LAYER met3 ;
        RECT 1396.000 2601.000 1400.000 2601.600 ;
      LAYER met3 ;
        RECT 300.065 2599.280 1396.000 2600.600 ;
        RECT 304.400 2597.880 1396.000 2599.280 ;
        RECT 300.065 2597.240 1396.000 2597.880 ;
        RECT 300.065 2595.840 1395.600 2597.240 ;
      LAYER met3 ;
        RECT 1396.000 2596.240 1400.000 2596.840 ;
      LAYER met3 ;
        RECT 300.065 2591.800 1396.000 2595.840 ;
        RECT 300.065 2590.400 1395.600 2591.800 ;
      LAYER met3 ;
        RECT 1396.000 2590.800 1400.000 2591.400 ;
      LAYER met3 ;
        RECT 300.065 2589.760 1396.000 2590.400 ;
        RECT 304.400 2588.360 1396.000 2589.760 ;
        RECT 300.065 2587.040 1396.000 2588.360 ;
        RECT 300.065 2585.640 1395.600 2587.040 ;
      LAYER met3 ;
        RECT 1396.000 2586.040 1400.000 2586.640 ;
      LAYER met3 ;
        RECT 300.065 2581.600 1396.000 2585.640 ;
        RECT 300.065 2580.240 1395.600 2581.600 ;
      LAYER met3 ;
        RECT 1396.000 2580.600 1400.000 2581.200 ;
      LAYER met3 ;
        RECT 304.400 2580.200 1395.600 2580.240 ;
        RECT 304.400 2578.840 1396.000 2580.200 ;
        RECT 300.065 2576.840 1396.000 2578.840 ;
        RECT 300.065 2575.440 1395.600 2576.840 ;
      LAYER met3 ;
        RECT 1396.000 2575.840 1400.000 2576.440 ;
      LAYER met3 ;
        RECT 300.065 2572.080 1396.000 2575.440 ;
        RECT 300.065 2570.720 1395.600 2572.080 ;
      LAYER met3 ;
        RECT 1396.000 2571.080 1400.000 2571.680 ;
      LAYER met3 ;
        RECT 304.400 2570.680 1395.600 2570.720 ;
        RECT 304.400 2569.320 1396.000 2570.680 ;
        RECT 300.065 2566.640 1396.000 2569.320 ;
        RECT 300.065 2565.240 1395.600 2566.640 ;
      LAYER met3 ;
        RECT 1396.000 2565.640 1400.000 2566.240 ;
      LAYER met3 ;
        RECT 300.065 2561.880 1396.000 2565.240 ;
        RECT 300.065 2561.200 1395.600 2561.880 ;
        RECT 304.400 2560.480 1395.600 2561.200 ;
      LAYER met3 ;
        RECT 1396.000 2560.880 1400.000 2561.480 ;
      LAYER met3 ;
        RECT 304.400 2559.800 1396.000 2560.480 ;
        RECT 300.065 2556.440 1396.000 2559.800 ;
        RECT 300.065 2555.040 1395.600 2556.440 ;
      LAYER met3 ;
        RECT 1396.000 2555.440 1400.000 2556.040 ;
      LAYER met3 ;
        RECT 300.065 2551.680 1396.000 2555.040 ;
        RECT 300.065 2551.000 1395.600 2551.680 ;
        RECT 304.400 2550.280 1395.600 2551.000 ;
      LAYER met3 ;
        RECT 1396.000 2550.680 1400.000 2551.280 ;
      LAYER met3 ;
        RECT 304.400 2549.600 1396.000 2550.280 ;
        RECT 300.065 2546.240 1396.000 2549.600 ;
        RECT 300.065 2544.840 1395.600 2546.240 ;
      LAYER met3 ;
        RECT 1396.000 2545.240 1400.000 2545.840 ;
      LAYER met3 ;
        RECT 300.065 2541.480 1396.000 2544.840 ;
        RECT 304.400 2540.080 1395.600 2541.480 ;
      LAYER met3 ;
        RECT 1396.000 2540.480 1400.000 2541.080 ;
      LAYER met3 ;
        RECT 300.065 2536.720 1396.000 2540.080 ;
        RECT 300.065 2535.320 1395.600 2536.720 ;
      LAYER met3 ;
        RECT 1396.000 2535.720 1400.000 2536.320 ;
      LAYER met3 ;
        RECT 300.065 2531.960 1396.000 2535.320 ;
        RECT 304.400 2531.280 1396.000 2531.960 ;
        RECT 304.400 2530.560 1395.600 2531.280 ;
        RECT 300.065 2529.880 1395.600 2530.560 ;
      LAYER met3 ;
        RECT 1396.000 2530.280 1400.000 2530.880 ;
      LAYER met3 ;
        RECT 300.065 2526.520 1396.000 2529.880 ;
        RECT 300.065 2525.120 1395.600 2526.520 ;
      LAYER met3 ;
        RECT 1396.000 2525.520 1400.000 2526.120 ;
      LAYER met3 ;
        RECT 300.065 2522.440 1396.000 2525.120 ;
        RECT 304.400 2521.080 1396.000 2522.440 ;
        RECT 304.400 2521.040 1395.600 2521.080 ;
        RECT 300.065 2519.680 1395.600 2521.040 ;
      LAYER met3 ;
        RECT 1396.000 2520.080 1400.000 2520.680 ;
      LAYER met3 ;
        RECT 300.065 2516.320 1396.000 2519.680 ;
        RECT 300.065 2514.920 1395.600 2516.320 ;
      LAYER met3 ;
        RECT 1396.000 2515.320 1400.000 2515.920 ;
      LAYER met3 ;
        RECT 300.065 2512.920 1396.000 2514.920 ;
        RECT 304.400 2511.520 1396.000 2512.920 ;
        RECT 300.065 2510.880 1396.000 2511.520 ;
        RECT 300.065 2509.480 1395.600 2510.880 ;
      LAYER met3 ;
        RECT 1396.000 2509.880 1400.000 2510.480 ;
      LAYER met3 ;
        RECT 300.065 2506.120 1396.000 2509.480 ;
        RECT 300.065 2504.720 1395.600 2506.120 ;
      LAYER met3 ;
        RECT 1396.000 2505.120 1400.000 2505.720 ;
      LAYER met3 ;
        RECT 300.065 2502.720 1396.000 2504.720 ;
        RECT 304.400 2501.360 1396.000 2502.720 ;
        RECT 304.400 2501.320 1395.600 2501.360 ;
        RECT 300.065 2499.960 1395.600 2501.320 ;
      LAYER met3 ;
        RECT 1396.000 2500.360 1400.000 2500.960 ;
      LAYER met3 ;
        RECT 300.065 2495.920 1396.000 2499.960 ;
        RECT 300.065 2494.520 1395.600 2495.920 ;
      LAYER met3 ;
        RECT 1396.000 2494.920 1400.000 2495.520 ;
      LAYER met3 ;
        RECT 300.065 2493.200 1396.000 2494.520 ;
        RECT 304.400 2491.800 1396.000 2493.200 ;
        RECT 300.065 2491.160 1396.000 2491.800 ;
        RECT 300.065 2489.760 1395.600 2491.160 ;
      LAYER met3 ;
        RECT 1396.000 2490.160 1400.000 2490.760 ;
      LAYER met3 ;
        RECT 300.065 2485.720 1396.000 2489.760 ;
        RECT 300.065 2484.320 1395.600 2485.720 ;
      LAYER met3 ;
        RECT 1396.000 2484.720 1400.000 2485.320 ;
      LAYER met3 ;
        RECT 300.065 2483.680 1396.000 2484.320 ;
        RECT 304.400 2482.280 1396.000 2483.680 ;
        RECT 300.065 2480.960 1396.000 2482.280 ;
        RECT 300.065 2479.560 1395.600 2480.960 ;
      LAYER met3 ;
        RECT 1396.000 2479.960 1400.000 2480.560 ;
      LAYER met3 ;
        RECT 300.065 2476.200 1396.000 2479.560 ;
        RECT 300.065 2474.800 1395.600 2476.200 ;
      LAYER met3 ;
        RECT 1396.000 2475.200 1400.000 2475.800 ;
      LAYER met3 ;
        RECT 300.065 2474.160 1396.000 2474.800 ;
        RECT 304.400 2472.760 1396.000 2474.160 ;
        RECT 300.065 2470.760 1396.000 2472.760 ;
        RECT 300.065 2469.360 1395.600 2470.760 ;
      LAYER met3 ;
        RECT 1396.000 2469.760 1400.000 2470.360 ;
      LAYER met3 ;
        RECT 300.065 2466.000 1396.000 2469.360 ;
        RECT 300.065 2464.640 1395.600 2466.000 ;
      LAYER met3 ;
        RECT 1396.000 2465.000 1400.000 2465.600 ;
      LAYER met3 ;
        RECT 304.400 2464.600 1395.600 2464.640 ;
        RECT 304.400 2463.240 1396.000 2464.600 ;
        RECT 300.065 2460.560 1396.000 2463.240 ;
        RECT 300.065 2459.160 1395.600 2460.560 ;
      LAYER met3 ;
        RECT 1396.000 2459.560 1400.000 2460.160 ;
      LAYER met3 ;
        RECT 300.065 2455.800 1396.000 2459.160 ;
        RECT 300.065 2454.440 1395.600 2455.800 ;
      LAYER met3 ;
        RECT 1396.000 2454.800 1400.000 2455.400 ;
      LAYER met3 ;
        RECT 304.400 2454.400 1395.600 2454.440 ;
        RECT 304.400 2453.040 1396.000 2454.400 ;
        RECT 300.065 2450.360 1396.000 2453.040 ;
        RECT 300.065 2448.960 1395.600 2450.360 ;
      LAYER met3 ;
        RECT 1396.000 2449.360 1400.000 2449.960 ;
      LAYER met3 ;
        RECT 300.065 2445.600 1396.000 2448.960 ;
        RECT 300.065 2444.920 1395.600 2445.600 ;
        RECT 304.400 2444.200 1395.600 2444.920 ;
      LAYER met3 ;
        RECT 1396.000 2444.600 1400.000 2445.200 ;
      LAYER met3 ;
        RECT 304.400 2443.520 1396.000 2444.200 ;
        RECT 300.065 2440.840 1396.000 2443.520 ;
        RECT 300.065 2439.440 1395.600 2440.840 ;
      LAYER met3 ;
        RECT 1396.000 2439.840 1400.000 2440.440 ;
      LAYER met3 ;
        RECT 300.065 2435.400 1396.000 2439.440 ;
        RECT 304.400 2434.000 1395.600 2435.400 ;
      LAYER met3 ;
        RECT 1396.000 2434.400 1400.000 2435.000 ;
      LAYER met3 ;
        RECT 300.065 2430.640 1396.000 2434.000 ;
        RECT 300.065 2429.240 1395.600 2430.640 ;
      LAYER met3 ;
        RECT 1396.000 2429.640 1400.000 2430.240 ;
      LAYER met3 ;
        RECT 300.065 2425.880 1396.000 2429.240 ;
        RECT 304.400 2425.200 1396.000 2425.880 ;
        RECT 304.400 2424.480 1395.600 2425.200 ;
        RECT 300.065 2423.800 1395.600 2424.480 ;
      LAYER met3 ;
        RECT 1396.000 2424.200 1400.000 2424.800 ;
      LAYER met3 ;
        RECT 300.065 2420.440 1396.000 2423.800 ;
        RECT 300.065 2419.040 1395.600 2420.440 ;
      LAYER met3 ;
        RECT 1396.000 2419.440 1400.000 2420.040 ;
      LAYER met3 ;
        RECT 300.065 2416.360 1396.000 2419.040 ;
        RECT 304.400 2415.000 1396.000 2416.360 ;
        RECT 304.400 2414.960 1395.600 2415.000 ;
        RECT 300.065 2413.600 1395.600 2414.960 ;
      LAYER met3 ;
        RECT 1396.000 2414.000 1400.000 2414.600 ;
      LAYER met3 ;
        RECT 300.065 2410.240 1396.000 2413.600 ;
        RECT 300.065 2408.840 1395.600 2410.240 ;
      LAYER met3 ;
        RECT 1396.000 2409.240 1400.000 2409.840 ;
      LAYER met3 ;
        RECT 300.065 2406.840 1396.000 2408.840 ;
        RECT 304.400 2405.480 1396.000 2406.840 ;
        RECT 304.400 2405.440 1395.600 2405.480 ;
        RECT 300.065 2404.080 1395.600 2405.440 ;
      LAYER met3 ;
        RECT 1396.000 2404.480 1400.000 2405.080 ;
      LAYER met3 ;
        RECT 300.065 2400.040 1396.000 2404.080 ;
        RECT 300.065 2398.640 1395.600 2400.040 ;
      LAYER met3 ;
        RECT 1396.000 2399.040 1400.000 2399.640 ;
      LAYER met3 ;
        RECT 300.065 2396.640 1396.000 2398.640 ;
        RECT 304.400 2395.280 1396.000 2396.640 ;
        RECT 304.400 2395.240 1395.600 2395.280 ;
        RECT 300.065 2393.880 1395.600 2395.240 ;
      LAYER met3 ;
        RECT 1396.000 2394.280 1400.000 2394.880 ;
      LAYER met3 ;
        RECT 300.065 2389.840 1396.000 2393.880 ;
        RECT 300.065 2388.440 1395.600 2389.840 ;
      LAYER met3 ;
        RECT 1396.000 2388.840 1400.000 2389.440 ;
      LAYER met3 ;
        RECT 300.065 2387.120 1396.000 2388.440 ;
        RECT 304.400 2385.720 1396.000 2387.120 ;
        RECT 300.065 2385.080 1396.000 2385.720 ;
        RECT 300.065 2383.680 1395.600 2385.080 ;
      LAYER met3 ;
        RECT 1396.000 2384.080 1400.000 2384.680 ;
      LAYER met3 ;
        RECT 300.065 2379.640 1396.000 2383.680 ;
        RECT 300.065 2378.240 1395.600 2379.640 ;
      LAYER met3 ;
        RECT 1396.000 2378.640 1400.000 2379.240 ;
      LAYER met3 ;
        RECT 300.065 2377.600 1396.000 2378.240 ;
        RECT 304.400 2376.200 1396.000 2377.600 ;
        RECT 300.065 2374.880 1396.000 2376.200 ;
        RECT 300.065 2373.480 1395.600 2374.880 ;
      LAYER met3 ;
        RECT 1396.000 2373.880 1400.000 2374.480 ;
      LAYER met3 ;
        RECT 300.065 2370.120 1396.000 2373.480 ;
        RECT 300.065 2368.720 1395.600 2370.120 ;
      LAYER met3 ;
        RECT 1396.000 2369.120 1400.000 2369.720 ;
      LAYER met3 ;
        RECT 300.065 2368.080 1396.000 2368.720 ;
        RECT 304.400 2366.680 1396.000 2368.080 ;
        RECT 300.065 2364.680 1396.000 2366.680 ;
        RECT 300.065 2363.280 1395.600 2364.680 ;
      LAYER met3 ;
        RECT 1396.000 2363.680 1400.000 2364.280 ;
      LAYER met3 ;
        RECT 300.065 2359.920 1396.000 2363.280 ;
        RECT 300.065 2358.560 1395.600 2359.920 ;
      LAYER met3 ;
        RECT 1396.000 2358.920 1400.000 2359.520 ;
      LAYER met3 ;
        RECT 304.400 2358.520 1395.600 2358.560 ;
        RECT 304.400 2357.160 1396.000 2358.520 ;
        RECT 300.065 2354.480 1396.000 2357.160 ;
        RECT 300.065 2353.080 1395.600 2354.480 ;
      LAYER met3 ;
        RECT 1396.000 2353.480 1400.000 2354.080 ;
      LAYER met3 ;
        RECT 300.065 2349.720 1396.000 2353.080 ;
        RECT 300.065 2348.360 1395.600 2349.720 ;
      LAYER met3 ;
        RECT 1396.000 2348.720 1400.000 2349.320 ;
      LAYER met3 ;
        RECT 304.400 2348.320 1395.600 2348.360 ;
        RECT 304.400 2346.960 1396.000 2348.320 ;
        RECT 300.065 2344.960 1396.000 2346.960 ;
        RECT 300.065 2343.560 1395.600 2344.960 ;
      LAYER met3 ;
        RECT 1396.000 2343.960 1400.000 2344.560 ;
      LAYER met3 ;
        RECT 300.065 2339.520 1396.000 2343.560 ;
        RECT 300.065 2338.840 1395.600 2339.520 ;
        RECT 304.400 2338.120 1395.600 2338.840 ;
      LAYER met3 ;
        RECT 1396.000 2338.520 1400.000 2339.120 ;
      LAYER met3 ;
        RECT 304.400 2337.440 1396.000 2338.120 ;
        RECT 300.065 2334.760 1396.000 2337.440 ;
        RECT 300.065 2333.360 1395.600 2334.760 ;
      LAYER met3 ;
        RECT 1396.000 2333.760 1400.000 2334.360 ;
      LAYER met3 ;
        RECT 300.065 2329.320 1396.000 2333.360 ;
        RECT 304.400 2327.920 1395.600 2329.320 ;
      LAYER met3 ;
        RECT 1396.000 2328.320 1400.000 2328.920 ;
      LAYER met3 ;
        RECT 300.065 2324.560 1396.000 2327.920 ;
        RECT 300.065 2323.160 1395.600 2324.560 ;
      LAYER met3 ;
        RECT 1396.000 2323.560 1400.000 2324.160 ;
      LAYER met3 ;
        RECT 300.065 2319.800 1396.000 2323.160 ;
        RECT 304.400 2319.120 1396.000 2319.800 ;
        RECT 304.400 2318.400 1395.600 2319.120 ;
        RECT 300.065 2317.720 1395.600 2318.400 ;
      LAYER met3 ;
        RECT 1396.000 2318.120 1400.000 2318.720 ;
      LAYER met3 ;
        RECT 300.065 2314.360 1396.000 2317.720 ;
        RECT 300.065 2312.960 1395.600 2314.360 ;
      LAYER met3 ;
        RECT 1396.000 2313.360 1400.000 2313.960 ;
      LAYER met3 ;
        RECT 300.065 2310.280 1396.000 2312.960 ;
        RECT 304.400 2309.600 1396.000 2310.280 ;
        RECT 304.400 2308.880 1395.600 2309.600 ;
        RECT 300.065 2308.200 1395.600 2308.880 ;
      LAYER met3 ;
        RECT 1396.000 2308.600 1400.000 2309.200 ;
      LAYER met3 ;
        RECT 300.065 2304.160 1396.000 2308.200 ;
        RECT 300.065 2302.760 1395.600 2304.160 ;
      LAYER met3 ;
        RECT 1396.000 2303.160 1400.000 2303.760 ;
      LAYER met3 ;
        RECT 300.065 2300.080 1396.000 2302.760 ;
        RECT 304.400 2299.400 1396.000 2300.080 ;
        RECT 304.400 2298.680 1395.600 2299.400 ;
        RECT 300.065 2298.000 1395.600 2298.680 ;
      LAYER met3 ;
        RECT 1396.000 2298.400 1400.000 2299.000 ;
      LAYER met3 ;
        RECT 300.065 2293.960 1396.000 2298.000 ;
        RECT 300.065 2292.560 1395.600 2293.960 ;
      LAYER met3 ;
        RECT 1396.000 2292.960 1400.000 2293.560 ;
      LAYER met3 ;
        RECT 300.065 2290.560 1396.000 2292.560 ;
        RECT 304.400 2289.200 1396.000 2290.560 ;
        RECT 304.400 2289.160 1395.600 2289.200 ;
        RECT 300.065 2287.800 1395.600 2289.160 ;
      LAYER met3 ;
        RECT 1396.000 2288.200 1400.000 2288.800 ;
      LAYER met3 ;
        RECT 300.065 2283.760 1396.000 2287.800 ;
        RECT 300.065 2282.360 1395.600 2283.760 ;
      LAYER met3 ;
        RECT 1396.000 2282.760 1400.000 2283.360 ;
      LAYER met3 ;
        RECT 300.065 2281.040 1396.000 2282.360 ;
        RECT 304.400 2279.640 1396.000 2281.040 ;
        RECT 300.065 2279.000 1396.000 2279.640 ;
        RECT 300.065 2277.600 1395.600 2279.000 ;
      LAYER met3 ;
        RECT 1396.000 2278.000 1400.000 2278.600 ;
      LAYER met3 ;
        RECT 300.065 2274.240 1396.000 2277.600 ;
        RECT 300.065 2272.840 1395.600 2274.240 ;
      LAYER met3 ;
        RECT 1396.000 2273.240 1400.000 2273.840 ;
      LAYER met3 ;
        RECT 300.065 2271.520 1396.000 2272.840 ;
        RECT 304.400 2270.120 1396.000 2271.520 ;
        RECT 300.065 2268.800 1396.000 2270.120 ;
        RECT 300.065 2267.400 1395.600 2268.800 ;
      LAYER met3 ;
        RECT 1396.000 2267.800 1400.000 2268.400 ;
      LAYER met3 ;
        RECT 300.065 2264.040 1396.000 2267.400 ;
        RECT 300.065 2262.640 1395.600 2264.040 ;
      LAYER met3 ;
        RECT 1396.000 2263.040 1400.000 2263.640 ;
      LAYER met3 ;
        RECT 300.065 2262.000 1396.000 2262.640 ;
        RECT 304.400 2260.600 1396.000 2262.000 ;
        RECT 300.065 2258.600 1396.000 2260.600 ;
        RECT 300.065 2257.200 1395.600 2258.600 ;
      LAYER met3 ;
        RECT 1396.000 2257.600 1400.000 2258.200 ;
      LAYER met3 ;
        RECT 300.065 2253.840 1396.000 2257.200 ;
        RECT 300.065 2252.440 1395.600 2253.840 ;
      LAYER met3 ;
        RECT 1396.000 2252.840 1400.000 2253.440 ;
      LAYER met3 ;
        RECT 300.065 2251.800 1396.000 2252.440 ;
        RECT 304.400 2250.400 1396.000 2251.800 ;
        RECT 300.065 2249.080 1396.000 2250.400 ;
        RECT 300.065 2247.680 1395.600 2249.080 ;
      LAYER met3 ;
        RECT 1396.000 2248.080 1400.000 2248.680 ;
      LAYER met3 ;
        RECT 300.065 2243.640 1396.000 2247.680 ;
        RECT 300.065 2242.280 1395.600 2243.640 ;
      LAYER met3 ;
        RECT 1396.000 2242.640 1400.000 2243.240 ;
      LAYER met3 ;
        RECT 304.400 2242.240 1395.600 2242.280 ;
        RECT 304.400 2240.880 1396.000 2242.240 ;
        RECT 300.065 2238.880 1396.000 2240.880 ;
        RECT 300.065 2237.480 1395.600 2238.880 ;
      LAYER met3 ;
        RECT 1396.000 2237.880 1400.000 2238.480 ;
      LAYER met3 ;
        RECT 300.065 2233.440 1396.000 2237.480 ;
        RECT 300.065 2232.760 1395.600 2233.440 ;
        RECT 304.400 2232.040 1395.600 2232.760 ;
      LAYER met3 ;
        RECT 1396.000 2232.440 1400.000 2233.040 ;
      LAYER met3 ;
        RECT 304.400 2231.360 1396.000 2232.040 ;
        RECT 300.065 2228.680 1396.000 2231.360 ;
        RECT 300.065 2227.280 1395.600 2228.680 ;
      LAYER met3 ;
        RECT 1396.000 2227.680 1400.000 2228.280 ;
      LAYER met3 ;
        RECT 300.065 2223.240 1396.000 2227.280 ;
        RECT 304.400 2221.840 1395.600 2223.240 ;
      LAYER met3 ;
        RECT 1396.000 2222.240 1400.000 2222.840 ;
      LAYER met3 ;
        RECT 300.065 2218.480 1396.000 2221.840 ;
        RECT 300.065 2217.080 1395.600 2218.480 ;
      LAYER met3 ;
        RECT 1396.000 2217.480 1400.000 2218.080 ;
      LAYER met3 ;
        RECT 300.065 2213.720 1396.000 2217.080 ;
        RECT 304.400 2212.320 1395.600 2213.720 ;
      LAYER met3 ;
        RECT 1396.000 2212.720 1400.000 2213.320 ;
      LAYER met3 ;
        RECT 300.065 2208.280 1396.000 2212.320 ;
        RECT 300.065 2206.880 1395.600 2208.280 ;
      LAYER met3 ;
        RECT 1396.000 2207.280 1400.000 2207.880 ;
      LAYER met3 ;
        RECT 300.065 2203.520 1396.000 2206.880 ;
        RECT 304.400 2202.120 1395.600 2203.520 ;
      LAYER met3 ;
        RECT 1396.000 2202.520 1400.000 2203.120 ;
      LAYER met3 ;
        RECT 300.065 2198.080 1396.000 2202.120 ;
        RECT 300.065 2196.680 1395.600 2198.080 ;
      LAYER met3 ;
        RECT 1396.000 2197.080 1400.000 2197.680 ;
      LAYER met3 ;
        RECT 300.065 2194.000 1396.000 2196.680 ;
        RECT 304.400 2193.320 1396.000 2194.000 ;
        RECT 304.400 2192.600 1395.600 2193.320 ;
        RECT 300.065 2191.920 1395.600 2192.600 ;
      LAYER met3 ;
        RECT 1396.000 2192.320 1400.000 2192.920 ;
      LAYER met3 ;
        RECT 300.065 2187.880 1396.000 2191.920 ;
        RECT 300.065 2186.480 1395.600 2187.880 ;
      LAYER met3 ;
        RECT 1396.000 2186.880 1400.000 2187.480 ;
      LAYER met3 ;
        RECT 300.065 2184.480 1396.000 2186.480 ;
        RECT 304.400 2183.120 1396.000 2184.480 ;
        RECT 304.400 2183.080 1395.600 2183.120 ;
        RECT 300.065 2181.720 1395.600 2183.080 ;
      LAYER met3 ;
        RECT 1396.000 2182.120 1400.000 2182.720 ;
      LAYER met3 ;
        RECT 300.065 2178.360 1396.000 2181.720 ;
        RECT 300.065 2176.960 1395.600 2178.360 ;
      LAYER met3 ;
        RECT 1396.000 2177.360 1400.000 2177.960 ;
      LAYER met3 ;
        RECT 300.065 2174.960 1396.000 2176.960 ;
        RECT 304.400 2173.560 1396.000 2174.960 ;
        RECT 300.065 2172.920 1396.000 2173.560 ;
        RECT 300.065 2171.520 1395.600 2172.920 ;
      LAYER met3 ;
        RECT 1396.000 2171.920 1400.000 2172.520 ;
      LAYER met3 ;
        RECT 300.065 2168.160 1396.000 2171.520 ;
        RECT 300.065 2166.760 1395.600 2168.160 ;
      LAYER met3 ;
        RECT 1396.000 2167.160 1400.000 2167.760 ;
      LAYER met3 ;
        RECT 300.065 2165.440 1396.000 2166.760 ;
        RECT 304.400 2164.040 1396.000 2165.440 ;
        RECT 300.065 2162.720 1396.000 2164.040 ;
        RECT 300.065 2161.320 1395.600 2162.720 ;
      LAYER met3 ;
        RECT 1396.000 2161.720 1400.000 2162.320 ;
      LAYER met3 ;
        RECT 300.065 2157.960 1396.000 2161.320 ;
        RECT 300.065 2156.560 1395.600 2157.960 ;
      LAYER met3 ;
        RECT 1396.000 2156.960 1400.000 2157.560 ;
      LAYER met3 ;
        RECT 300.065 2155.920 1396.000 2156.560 ;
        RECT 304.400 2154.520 1396.000 2155.920 ;
        RECT 300.065 2153.200 1396.000 2154.520 ;
        RECT 300.065 2151.800 1395.600 2153.200 ;
      LAYER met3 ;
        RECT 1396.000 2152.200 1400.000 2152.800 ;
      LAYER met3 ;
        RECT 300.065 2147.760 1396.000 2151.800 ;
        RECT 300.065 2146.360 1395.600 2147.760 ;
      LAYER met3 ;
        RECT 1396.000 2147.250 1400.000 2147.360 ;
        RECT 1407.665 2147.250 1407.995 2147.265 ;
        RECT 1396.000 2146.950 1407.995 2147.250 ;
        RECT 1396.000 2146.760 1400.000 2146.950 ;
        RECT 1407.665 2146.935 1407.995 2146.950 ;
      LAYER met3 ;
        RECT 300.065 2145.720 1396.000 2146.360 ;
        RECT 304.400 2144.320 1396.000 2145.720 ;
        RECT 300.065 2143.000 1396.000 2144.320 ;
        RECT 300.065 2141.600 1395.600 2143.000 ;
      LAYER met3 ;
        RECT 1396.000 2142.490 1400.000 2142.600 ;
        RECT 1407.665 2142.490 1407.995 2142.505 ;
        RECT 1396.000 2142.190 1407.995 2142.490 ;
        RECT 1396.000 2142.000 1400.000 2142.190 ;
        RECT 1407.665 2142.175 1407.995 2142.190 ;
      LAYER met3 ;
        RECT 300.065 2137.560 1396.000 2141.600 ;
        RECT 300.065 2136.200 1395.600 2137.560 ;
      LAYER met3 ;
        RECT 1396.000 2137.050 1400.000 2137.160 ;
        RECT 1408.125 2137.050 1408.455 2137.065 ;
        RECT 1396.000 2136.750 1408.455 2137.050 ;
        RECT 1396.000 2136.560 1400.000 2136.750 ;
        RECT 1408.125 2136.735 1408.455 2136.750 ;
      LAYER met3 ;
        RECT 304.400 2136.160 1395.600 2136.200 ;
        RECT 304.400 2134.800 1396.000 2136.160 ;
        RECT 300.065 2132.800 1396.000 2134.800 ;
        RECT 300.065 2131.400 1395.600 2132.800 ;
      LAYER met3 ;
        RECT 1396.000 2132.290 1400.000 2132.400 ;
        RECT 1407.665 2132.290 1407.995 2132.305 ;
        RECT 1396.000 2131.990 1407.995 2132.290 ;
        RECT 1396.000 2131.800 1400.000 2131.990 ;
        RECT 1407.665 2131.975 1407.995 2131.990 ;
      LAYER met3 ;
        RECT 300.065 2127.360 1396.000 2131.400 ;
        RECT 300.065 2126.680 1395.600 2127.360 ;
        RECT 304.400 2125.960 1395.600 2126.680 ;
      LAYER met3 ;
        RECT 1396.000 2126.850 1400.000 2126.960 ;
        RECT 1407.665 2126.850 1407.995 2126.865 ;
        RECT 1396.000 2126.550 1407.995 2126.850 ;
        RECT 1396.000 2126.360 1400.000 2126.550 ;
        RECT 1407.665 2126.535 1407.995 2126.550 ;
      LAYER met3 ;
        RECT 304.400 2125.280 1396.000 2125.960 ;
        RECT 300.065 2122.600 1396.000 2125.280 ;
        RECT 300.065 2121.200 1395.600 2122.600 ;
      LAYER met3 ;
        RECT 1396.000 2122.090 1400.000 2122.200 ;
        RECT 1407.665 2122.090 1407.995 2122.105 ;
        RECT 1396.000 2121.790 1407.995 2122.090 ;
        RECT 1396.000 2121.600 1400.000 2121.790 ;
        RECT 1407.665 2121.775 1407.995 2121.790 ;
      LAYER met3 ;
        RECT 300.065 2117.840 1396.000 2121.200 ;
        RECT 300.065 2117.160 1395.600 2117.840 ;
        RECT 304.400 2116.440 1395.600 2117.160 ;
      LAYER met3 ;
        RECT 1396.000 2117.330 1400.000 2117.440 ;
        RECT 1408.125 2117.330 1408.455 2117.345 ;
        RECT 1396.000 2117.030 1408.455 2117.330 ;
        RECT 1396.000 2116.840 1400.000 2117.030 ;
        RECT 1408.125 2117.015 1408.455 2117.030 ;
      LAYER met3 ;
        RECT 304.400 2115.760 1396.000 2116.440 ;
        RECT 300.065 2112.400 1396.000 2115.760 ;
        RECT 300.065 2111.000 1395.600 2112.400 ;
      LAYER met3 ;
        RECT 1396.000 2111.890 1400.000 2112.000 ;
        RECT 1407.665 2111.890 1407.995 2111.905 ;
        RECT 1396.000 2111.590 1407.995 2111.890 ;
        RECT 1396.000 2111.400 1400.000 2111.590 ;
        RECT 1407.665 2111.575 1407.995 2111.590 ;
      LAYER met3 ;
        RECT 300.065 2107.640 1396.000 2111.000 ;
        RECT 304.400 2106.240 1395.600 2107.640 ;
      LAYER met3 ;
        RECT 1396.000 2107.130 1400.000 2107.240 ;
        RECT 1407.665 2107.130 1407.995 2107.145 ;
        RECT 1396.000 2106.830 1407.995 2107.130 ;
        RECT 1396.000 2106.640 1400.000 2106.830 ;
        RECT 1407.665 2106.815 1407.995 2106.830 ;
      LAYER met3 ;
        RECT 300.065 2102.200 1396.000 2106.240 ;
        RECT 300.065 2100.800 1395.600 2102.200 ;
      LAYER met3 ;
        RECT 1396.000 2101.690 1400.000 2101.800 ;
        RECT 1407.665 2101.690 1407.995 2101.705 ;
        RECT 1396.000 2101.390 1407.995 2101.690 ;
        RECT 1396.000 2101.200 1400.000 2101.390 ;
        RECT 1407.665 2101.375 1407.995 2101.390 ;
      LAYER met3 ;
        RECT 300.065 2097.440 1396.000 2100.800 ;
        RECT 304.400 2096.040 1395.600 2097.440 ;
      LAYER met3 ;
        RECT 1396.000 2096.930 1400.000 2097.040 ;
        RECT 1408.125 2096.930 1408.455 2096.945 ;
        RECT 1396.000 2096.630 1408.455 2096.930 ;
        RECT 1396.000 2096.440 1400.000 2096.630 ;
        RECT 1408.125 2096.615 1408.455 2096.630 ;
      LAYER met3 ;
        RECT 300.065 2092.000 1396.000 2096.040 ;
        RECT 300.065 2090.600 1395.600 2092.000 ;
      LAYER met3 ;
        RECT 1396.000 2091.490 1400.000 2091.600 ;
        RECT 1407.665 2091.490 1407.995 2091.505 ;
        RECT 1396.000 2091.190 1407.995 2091.490 ;
        RECT 1396.000 2091.000 1400.000 2091.190 ;
        RECT 1407.665 2091.175 1407.995 2091.190 ;
      LAYER met3 ;
        RECT 300.065 2087.920 1396.000 2090.600 ;
        RECT 304.400 2087.240 1396.000 2087.920 ;
        RECT 304.400 2086.520 1395.600 2087.240 ;
        RECT 300.065 2085.840 1395.600 2086.520 ;
      LAYER met3 ;
        RECT 1396.000 2086.730 1400.000 2086.840 ;
        RECT 1414.105 2086.730 1414.435 2086.745 ;
        RECT 1396.000 2086.430 1414.435 2086.730 ;
        RECT 1396.000 2086.240 1400.000 2086.430 ;
        RECT 1414.105 2086.415 1414.435 2086.430 ;
      LAYER met3 ;
        RECT 300.065 2082.480 1396.000 2085.840 ;
        RECT 300.065 2081.080 1395.600 2082.480 ;
      LAYER met3 ;
        RECT 1396.000 2081.970 1400.000 2082.080 ;
        RECT 1411.345 2081.970 1411.675 2081.985 ;
        RECT 1396.000 2081.670 1411.675 2081.970 ;
        RECT 1396.000 2081.480 1400.000 2081.670 ;
        RECT 1411.345 2081.655 1411.675 2081.670 ;
      LAYER met3 ;
        RECT 300.065 2078.400 1396.000 2081.080 ;
        RECT 304.400 2077.040 1396.000 2078.400 ;
        RECT 304.400 2077.000 1395.600 2077.040 ;
        RECT 300.065 2075.640 1395.600 2077.000 ;
      LAYER met3 ;
        RECT 1396.000 2076.530 1400.000 2076.640 ;
        RECT 1408.585 2076.530 1408.915 2076.545 ;
        RECT 1396.000 2076.230 1408.915 2076.530 ;
        RECT 1396.000 2076.040 1400.000 2076.230 ;
        RECT 1408.585 2076.215 1408.915 2076.230 ;
      LAYER met3 ;
        RECT 300.065 2072.280 1396.000 2075.640 ;
        RECT 300.065 2070.880 1395.600 2072.280 ;
      LAYER met3 ;
        RECT 1396.000 2071.770 1400.000 2071.880 ;
        RECT 1410.425 2071.770 1410.755 2071.785 ;
        RECT 1396.000 2071.470 1410.755 2071.770 ;
        RECT 1396.000 2071.280 1400.000 2071.470 ;
        RECT 1410.425 2071.455 1410.755 2071.470 ;
      LAYER met3 ;
        RECT 300.065 2068.880 1396.000 2070.880 ;
      LAYER met3 ;
        RECT 1835.465 2069.730 1835.795 2069.745 ;
        RECT 1838.430 2069.730 1838.810 2069.740 ;
        RECT 1835.465 2069.430 1838.810 2069.730 ;
        RECT 1835.465 2069.415 1835.795 2069.430 ;
        RECT 1838.430 2069.420 1838.810 2069.430 ;
        RECT 1842.365 2069.730 1842.695 2069.745 ;
        RECT 1844.870 2069.730 1845.250 2069.740 ;
        RECT 1842.365 2069.430 1845.250 2069.730 ;
        RECT 1842.365 2069.415 1842.695 2069.430 ;
        RECT 1844.870 2069.420 1845.250 2069.430 ;
        RECT 1849.265 2069.730 1849.595 2069.745 ;
        RECT 1851.310 2069.730 1851.690 2069.740 ;
        RECT 1849.265 2069.430 1851.690 2069.730 ;
        RECT 1849.265 2069.415 1849.595 2069.430 ;
        RECT 1851.310 2069.420 1851.690 2069.430 ;
        RECT 1856.165 2069.730 1856.495 2069.745 ;
        RECT 1863.065 2069.740 1863.395 2069.745 ;
        RECT 1869.965 2069.740 1870.295 2069.745 ;
        RECT 1857.750 2069.730 1858.130 2069.740 ;
        RECT 1863.065 2069.730 1863.650 2069.740 ;
        RECT 1856.165 2069.430 1858.130 2069.730 ;
        RECT 1862.840 2069.430 1863.650 2069.730 ;
        RECT 1856.165 2069.415 1856.495 2069.430 ;
        RECT 1857.750 2069.420 1858.130 2069.430 ;
        RECT 1863.065 2069.420 1863.650 2069.430 ;
        RECT 1869.710 2069.730 1870.295 2069.740 ;
        RECT 1876.865 2069.730 1877.195 2069.745 ;
        RECT 1879.830 2069.730 1880.210 2069.740 ;
        RECT 1869.710 2069.430 1870.520 2069.730 ;
        RECT 1876.865 2069.430 1880.210 2069.730 ;
        RECT 1869.710 2069.420 1870.295 2069.430 ;
        RECT 1863.065 2069.415 1863.395 2069.420 ;
        RECT 1869.965 2069.415 1870.295 2069.420 ;
        RECT 1876.865 2069.415 1877.195 2069.430 ;
        RECT 1879.830 2069.420 1880.210 2069.430 ;
        RECT 1883.765 2069.730 1884.095 2069.745 ;
        RECT 1886.270 2069.730 1886.650 2069.740 ;
        RECT 1883.765 2069.430 1886.650 2069.730 ;
        RECT 1883.765 2069.415 1884.095 2069.430 ;
        RECT 1886.270 2069.420 1886.650 2069.430 ;
        RECT 1890.665 2069.730 1890.995 2069.745 ;
        RECT 1891.790 2069.730 1892.170 2069.740 ;
        RECT 1890.665 2069.430 1892.170 2069.730 ;
        RECT 1890.665 2069.415 1890.995 2069.430 ;
        RECT 1891.790 2069.420 1892.170 2069.430 ;
        RECT 1897.565 2069.730 1897.895 2069.745 ;
        RECT 1904.465 2069.740 1904.795 2069.745 ;
        RECT 1911.365 2069.740 1911.695 2069.745 ;
        RECT 1898.230 2069.730 1898.610 2069.740 ;
        RECT 1904.465 2069.730 1905.050 2069.740 ;
        RECT 1897.565 2069.430 1898.610 2069.730 ;
        RECT 1904.240 2069.430 1905.050 2069.730 ;
        RECT 1897.565 2069.415 1897.895 2069.430 ;
        RECT 1898.230 2069.420 1898.610 2069.430 ;
        RECT 1904.465 2069.420 1905.050 2069.430 ;
        RECT 1911.110 2069.730 1911.695 2069.740 ;
        RECT 1925.165 2069.730 1925.495 2069.745 ;
        RECT 1925.830 2069.730 1926.210 2069.740 ;
        RECT 1911.110 2069.430 1911.920 2069.730 ;
        RECT 1925.165 2069.430 1926.210 2069.730 ;
        RECT 1911.110 2069.420 1911.695 2069.430 ;
        RECT 1904.465 2069.415 1904.795 2069.420 ;
        RECT 1911.365 2069.415 1911.695 2069.420 ;
        RECT 1925.165 2069.415 1925.495 2069.430 ;
        RECT 1925.830 2069.420 1926.210 2069.430 ;
      LAYER met3 ;
        RECT 304.400 2067.480 1396.000 2068.880 ;
      LAYER met3 ;
        RECT 1870.425 2069.050 1870.755 2069.065 ;
        RECT 1873.390 2069.050 1873.770 2069.060 ;
        RECT 1870.425 2068.750 1873.770 2069.050 ;
        RECT 1870.425 2068.735 1870.755 2068.750 ;
        RECT 1873.390 2068.740 1873.770 2068.750 ;
        RECT 1911.825 2069.050 1912.155 2069.065 ;
        RECT 1914.790 2069.050 1915.170 2069.060 ;
        RECT 1911.825 2068.750 1915.170 2069.050 ;
        RECT 1911.825 2068.735 1912.155 2068.750 ;
        RECT 1914.790 2068.740 1915.170 2068.750 ;
        RECT 1919.185 2069.050 1919.515 2069.065 ;
        RECT 1920.310 2069.050 1920.690 2069.060 ;
        RECT 1919.185 2068.750 1920.690 2069.050 ;
        RECT 1919.185 2068.735 1919.515 2068.750 ;
        RECT 1920.310 2068.740 1920.690 2068.750 ;
        RECT 1980.365 2068.370 1980.695 2068.385 ;
        RECT 1987.265 2068.380 1987.595 2068.385 ;
        RECT 1981.950 2068.370 1982.330 2068.380 ;
        RECT 1987.265 2068.370 1987.850 2068.380 ;
        RECT 1980.365 2068.070 1982.330 2068.370 ;
        RECT 1987.040 2068.070 1987.850 2068.370 ;
        RECT 1980.365 2068.055 1980.695 2068.070 ;
        RECT 1981.950 2068.060 1982.330 2068.070 ;
        RECT 1987.265 2068.060 1987.850 2068.070 ;
        RECT 1987.265 2068.055 1987.595 2068.060 ;
        RECT 2028.665 2067.700 2028.995 2067.705 ;
        RECT 2028.665 2067.690 2029.250 2067.700 ;
      LAYER met3 ;
        RECT 300.065 2066.840 1396.000 2067.480 ;
      LAYER met3 ;
        RECT 2028.440 2067.390 2029.250 2067.690 ;
        RECT 2028.665 2067.380 2029.250 2067.390 ;
        RECT 2028.665 2067.375 2028.995 2067.380 ;
        RECT 1841.445 2067.020 1841.775 2067.025 ;
        RECT 1841.190 2067.010 1841.775 2067.020 ;
      LAYER met3 ;
        RECT 300.065 2065.440 1395.600 2066.840 ;
      LAYER met3 ;
        RECT 1840.990 2066.710 1841.775 2067.010 ;
        RECT 1841.190 2066.700 1841.775 2066.710 ;
        RECT 1841.445 2066.695 1841.775 2066.700 ;
        RECT 1843.745 2067.010 1844.075 2067.025 ;
        RECT 1848.805 2067.020 1849.135 2067.025 ;
        RECT 1890.205 2067.020 1890.535 2067.025 ;
        RECT 1941.725 2067.020 1942.055 2067.025 ;
        RECT 1848.550 2067.010 1849.135 2067.020 ;
        RECT 1889.950 2067.010 1890.535 2067.020 ;
        RECT 1941.470 2067.010 1942.055 2067.020 ;
        RECT 1843.745 2066.710 1849.540 2067.010 ;
        RECT 1889.750 2066.710 1890.535 2067.010 ;
        RECT 1941.270 2066.710 1942.055 2067.010 ;
        RECT 1843.745 2066.695 1844.075 2066.710 ;
        RECT 1848.550 2066.700 1849.135 2066.710 ;
        RECT 1889.950 2066.700 1890.535 2066.710 ;
        RECT 1941.470 2066.700 1942.055 2066.710 ;
        RECT 1848.805 2066.695 1849.135 2066.700 ;
        RECT 1890.205 2066.695 1890.535 2066.700 ;
        RECT 1941.725 2066.695 1942.055 2066.700 ;
        RECT 2021.765 2067.010 2022.095 2067.025 ;
        RECT 2023.350 2067.010 2023.730 2067.020 ;
        RECT 2021.765 2066.710 2023.730 2067.010 ;
        RECT 2021.765 2066.695 2022.095 2066.710 ;
        RECT 2023.350 2066.700 2023.730 2066.710 ;
        RECT 1396.000 2066.330 1400.000 2066.440 ;
        RECT 1414.105 2066.330 1414.435 2066.345 ;
        RECT 1396.000 2066.030 1414.435 2066.330 ;
        RECT 1396.000 2065.840 1400.000 2066.030 ;
        RECT 1414.105 2066.015 1414.435 2066.030 ;
        RECT 1849.265 2066.330 1849.595 2066.345 ;
        RECT 1854.990 2066.330 1855.370 2066.340 ;
        RECT 1849.265 2066.030 1855.370 2066.330 ;
        RECT 1849.265 2066.015 1849.595 2066.030 ;
        RECT 1854.990 2066.020 1855.370 2066.030 ;
        RECT 1898.025 2066.330 1898.355 2066.345 ;
        RECT 1900.990 2066.330 1901.370 2066.340 ;
        RECT 1898.025 2066.030 1901.370 2066.330 ;
        RECT 1898.025 2066.015 1898.355 2066.030 ;
        RECT 1900.990 2066.020 1901.370 2066.030 ;
        RECT 1932.065 2066.330 1932.395 2066.345 ;
        RECT 1934.110 2066.330 1934.490 2066.340 ;
        RECT 1932.065 2066.030 1934.490 2066.330 ;
        RECT 1932.065 2066.015 1932.395 2066.030 ;
        RECT 1934.110 2066.020 1934.490 2066.030 ;
        RECT 2007.965 2066.330 2008.295 2066.345 ;
        RECT 2011.390 2066.330 2011.770 2066.340 ;
        RECT 2007.965 2066.030 2011.770 2066.330 ;
        RECT 2007.965 2066.015 2008.295 2066.030 ;
        RECT 2011.390 2066.020 2011.770 2066.030 ;
        RECT 2015.785 2066.330 2016.115 2066.345 ;
        RECT 2016.910 2066.330 2017.290 2066.340 ;
        RECT 2015.785 2066.030 2017.290 2066.330 ;
        RECT 2015.785 2066.015 2016.115 2066.030 ;
        RECT 2016.910 2066.020 2017.290 2066.030 ;
        RECT 2035.565 2066.330 2035.895 2066.345 ;
        RECT 2037.150 2066.330 2037.530 2066.340 ;
        RECT 2035.565 2066.030 2037.530 2066.330 ;
        RECT 2035.565 2066.015 2035.895 2066.030 ;
        RECT 2037.150 2066.020 2037.530 2066.030 ;
        RECT 1859.845 2065.660 1860.175 2065.665 ;
        RECT 1859.590 2065.650 1860.175 2065.660 ;
      LAYER met3 ;
        RECT 300.065 2062.080 1396.000 2065.440 ;
      LAYER met3 ;
        RECT 1859.390 2065.350 1860.175 2065.650 ;
        RECT 1859.590 2065.340 1860.175 2065.350 ;
        RECT 1859.845 2065.335 1860.175 2065.340 ;
        RECT 1864.905 2065.660 1865.235 2065.665 ;
        RECT 1864.905 2065.650 1865.490 2065.660 ;
        RECT 1893.885 2065.650 1894.215 2065.665 ;
        RECT 1907.685 2065.660 1908.015 2065.665 ;
        RECT 1894.550 2065.650 1894.930 2065.660 ;
        RECT 1907.430 2065.650 1908.015 2065.660 ;
        RECT 1864.905 2065.350 1865.690 2065.650 ;
        RECT 1893.885 2065.350 1894.930 2065.650 ;
        RECT 1907.230 2065.350 1908.015 2065.650 ;
        RECT 1864.905 2065.340 1865.490 2065.350 ;
        RECT 1864.905 2065.335 1865.235 2065.340 ;
        RECT 1893.885 2065.335 1894.215 2065.350 ;
        RECT 1894.550 2065.340 1894.930 2065.350 ;
        RECT 1907.430 2065.340 1908.015 2065.350 ;
        RECT 1907.685 2065.335 1908.015 2065.340 ;
        RECT 1911.365 2065.650 1911.695 2065.665 ;
        RECT 1912.030 2065.650 1912.410 2065.660 ;
        RECT 1911.365 2065.350 1912.410 2065.650 ;
        RECT 1911.365 2065.335 1911.695 2065.350 ;
        RECT 1912.030 2065.340 1912.410 2065.350 ;
        RECT 1935.950 2065.650 1936.330 2065.660 ;
        RECT 1936.665 2065.650 1936.995 2065.665 ;
        RECT 1935.950 2065.350 1936.995 2065.650 ;
        RECT 1935.950 2065.340 1936.330 2065.350 ;
        RECT 1936.665 2065.335 1936.995 2065.350 ;
        RECT 1994.165 2065.650 1994.495 2065.665 ;
        RECT 1999.430 2065.650 1999.810 2065.660 ;
        RECT 1994.165 2065.350 1999.810 2065.650 ;
        RECT 1994.165 2065.335 1994.495 2065.350 ;
        RECT 1999.430 2065.340 1999.810 2065.350 ;
        RECT 2042.465 2065.650 2042.795 2065.665 ;
        RECT 2043.590 2065.650 2043.970 2065.660 ;
        RECT 2042.465 2065.350 2043.970 2065.650 ;
        RECT 2042.465 2065.335 2042.795 2065.350 ;
        RECT 2043.590 2065.340 2043.970 2065.350 ;
        RECT 1871.805 2064.980 1872.135 2064.985 ;
        RECT 1917.805 2064.980 1918.135 2064.985 ;
        RECT 1871.550 2064.970 1872.135 2064.980 ;
        RECT 1917.550 2064.970 1918.135 2064.980 ;
        RECT 1871.350 2064.670 1872.135 2064.970 ;
        RECT 1917.350 2064.670 1918.135 2064.970 ;
        RECT 1871.550 2064.660 1872.135 2064.670 ;
        RECT 1917.550 2064.660 1918.135 2064.670 ;
        RECT 1923.990 2064.970 1924.370 2064.980 ;
        RECT 1924.705 2064.970 1925.035 2064.985 ;
        RECT 1923.990 2064.670 1925.035 2064.970 ;
        RECT 1923.990 2064.660 1924.370 2064.670 ;
        RECT 1871.805 2064.655 1872.135 2064.660 ;
        RECT 1917.805 2064.655 1918.135 2064.660 ;
        RECT 1924.705 2064.655 1925.035 2064.670 ;
        RECT 1929.510 2064.970 1929.890 2064.980 ;
        RECT 1930.225 2064.970 1930.555 2064.985 ;
        RECT 1929.510 2064.670 1930.555 2064.970 ;
        RECT 1929.510 2064.660 1929.890 2064.670 ;
        RECT 1930.225 2064.655 1930.555 2064.670 ;
        RECT 2001.065 2064.970 2001.395 2064.985 ;
        RECT 2005.870 2064.970 2006.250 2064.980 ;
        RECT 2001.065 2064.670 2006.250 2064.970 ;
        RECT 2001.065 2064.655 2001.395 2064.670 ;
        RECT 2005.870 2064.660 2006.250 2064.670 ;
        RECT 1877.325 2064.300 1877.655 2064.305 ;
        RECT 1882.845 2064.300 1883.175 2064.305 ;
        RECT 1877.070 2064.290 1877.655 2064.300 ;
        RECT 1882.590 2064.290 1883.175 2064.300 ;
        RECT 1876.870 2063.990 1877.655 2064.290 ;
        RECT 1882.390 2063.990 1883.175 2064.290 ;
        RECT 1877.070 2063.980 1877.655 2063.990 ;
        RECT 1882.590 2063.980 1883.175 2063.990 ;
        RECT 1877.325 2063.975 1877.655 2063.980 ;
        RECT 1882.845 2063.975 1883.175 2063.980 ;
        RECT 1966.565 2064.290 1966.895 2064.305 ;
        RECT 1967.230 2064.290 1967.610 2064.300 ;
        RECT 1966.565 2063.990 1967.610 2064.290 ;
        RECT 1966.565 2063.975 1966.895 2063.990 ;
        RECT 1967.230 2063.980 1967.610 2063.990 ;
        RECT 1987.265 2064.290 1987.595 2064.305 ;
        RECT 1992.990 2064.290 1993.370 2064.300 ;
        RECT 1987.265 2063.990 1993.370 2064.290 ;
        RECT 1987.265 2063.975 1987.595 2063.990 ;
        RECT 1992.990 2063.980 1993.370 2063.990 ;
        RECT 1948.165 2063.620 1948.495 2063.625 ;
        RECT 1954.605 2063.620 1954.935 2063.625 ;
        RECT 1947.910 2063.610 1948.495 2063.620 ;
        RECT 1954.350 2063.610 1954.935 2063.620 ;
        RECT 1947.710 2063.310 1948.495 2063.610 ;
        RECT 1954.150 2063.310 1954.935 2063.610 ;
        RECT 1947.910 2063.300 1948.495 2063.310 ;
        RECT 1954.350 2063.300 1954.935 2063.310 ;
        RECT 1948.165 2063.295 1948.495 2063.300 ;
        RECT 1954.605 2063.295 1954.935 2063.300 ;
        RECT 1958.745 2063.620 1959.075 2063.625 ;
        RECT 1965.645 2063.620 1965.975 2063.625 ;
        RECT 1958.745 2063.610 1959.330 2063.620 ;
        RECT 1965.390 2063.610 1965.975 2063.620 ;
        RECT 1958.745 2063.310 1959.530 2063.610 ;
        RECT 1965.190 2063.310 1965.975 2063.610 ;
        RECT 1958.745 2063.300 1959.330 2063.310 ;
        RECT 1965.390 2063.300 1965.975 2063.310 ;
        RECT 1958.745 2063.295 1959.075 2063.300 ;
        RECT 1965.645 2063.295 1965.975 2063.300 ;
        RECT 1969.785 2063.620 1970.115 2063.625 ;
        RECT 1973.465 2063.620 1973.795 2063.625 ;
        RECT 1976.685 2063.620 1977.015 2063.625 ;
        RECT 1980.365 2063.620 1980.695 2063.625 ;
        RECT 1969.785 2063.610 1970.370 2063.620 ;
        RECT 1973.465 2063.610 1974.050 2063.620 ;
        RECT 1976.430 2063.610 1977.015 2063.620 ;
        RECT 1969.785 2063.310 1970.570 2063.610 ;
        RECT 1973.240 2063.310 1974.050 2063.610 ;
        RECT 1976.230 2063.310 1977.015 2063.610 ;
        RECT 1969.785 2063.300 1970.370 2063.310 ;
        RECT 1973.465 2063.300 1974.050 2063.310 ;
        RECT 1976.430 2063.300 1977.015 2063.310 ;
        RECT 1980.110 2063.610 1980.695 2063.620 ;
        RECT 2028.665 2063.610 2028.995 2063.625 ;
        RECT 2031.630 2063.610 2032.010 2063.620 ;
        RECT 1980.110 2063.310 1980.920 2063.610 ;
        RECT 2028.665 2063.310 2032.010 2063.610 ;
        RECT 1980.110 2063.300 1980.695 2063.310 ;
        RECT 1969.785 2063.295 1970.115 2063.300 ;
        RECT 1973.465 2063.295 1973.795 2063.300 ;
        RECT 1976.685 2063.295 1977.015 2063.300 ;
        RECT 1980.365 2063.295 1980.695 2063.300 ;
        RECT 2028.665 2063.295 2028.995 2063.310 ;
        RECT 2031.630 2063.300 2032.010 2063.310 ;
      LAYER met3 ;
        RECT 300.065 2060.680 1395.600 2062.080 ;
      LAYER met3 ;
        RECT 1396.000 2061.570 1400.000 2061.680 ;
        RECT 1410.425 2061.570 1410.755 2061.585 ;
        RECT 1396.000 2061.270 1410.755 2061.570 ;
        RECT 1396.000 2061.080 1400.000 2061.270 ;
        RECT 1410.425 2061.255 1410.755 2061.270 ;
      LAYER met3 ;
        RECT 300.065 2059.360 1396.000 2060.680 ;
        RECT 304.400 2057.960 1396.000 2059.360 ;
      LAYER met3 ;
        RECT 1940.345 2058.860 1940.675 2058.865 ;
        RECT 1940.345 2058.850 1940.930 2058.860 ;
        RECT 1940.120 2058.550 1940.930 2058.850 ;
        RECT 1940.345 2058.540 1940.930 2058.550 ;
        RECT 1940.345 2058.535 1940.675 2058.540 ;
        RECT 1955.065 2058.180 1955.395 2058.185 ;
        RECT 1987.265 2058.180 1987.595 2058.185 ;
        RECT 1995.545 2058.180 1995.875 2058.185 ;
        RECT 1955.065 2058.170 1955.650 2058.180 ;
        RECT 1987.265 2058.170 1987.650 2058.180 ;
        RECT 1995.545 2058.170 1996.130 2058.180 ;
      LAYER met3 ;
        RECT 300.065 2056.640 1396.000 2057.960 ;
      LAYER met3 ;
        RECT 1954.840 2057.870 1955.650 2058.170 ;
        RECT 1986.840 2057.870 1987.650 2058.170 ;
        RECT 1995.320 2057.870 1996.130 2058.170 ;
        RECT 1955.065 2057.860 1955.650 2057.870 ;
        RECT 1987.265 2057.860 1987.650 2057.870 ;
        RECT 1995.545 2057.860 1996.130 2057.870 ;
        RECT 1955.065 2057.855 1955.395 2057.860 ;
        RECT 1987.265 2057.855 1987.595 2057.860 ;
        RECT 1995.545 2057.855 1995.875 2057.860 ;
        RECT 1946.325 2057.500 1946.655 2057.505 ;
        RECT 1990.025 2057.500 1990.355 2057.505 ;
        RECT 2004.745 2057.500 2005.075 2057.505 ;
        RECT 2016.245 2057.500 2016.575 2057.505 ;
        RECT 1946.325 2057.490 1946.770 2057.500 ;
        RECT 1990.025 2057.490 1990.610 2057.500 ;
        RECT 2004.745 2057.490 2005.170 2057.500 ;
        RECT 2016.245 2057.490 2016.850 2057.500 ;
        RECT 1945.960 2057.190 1946.770 2057.490 ;
        RECT 1989.800 2057.190 1990.610 2057.490 ;
        RECT 2004.360 2057.190 2005.170 2057.490 ;
        RECT 2016.040 2057.190 2016.850 2057.490 ;
        RECT 1946.325 2057.180 1946.770 2057.190 ;
        RECT 1990.025 2057.180 1990.610 2057.190 ;
        RECT 2004.745 2057.180 2005.170 2057.190 ;
        RECT 2016.245 2057.180 2016.850 2057.190 ;
        RECT 1946.325 2057.175 1946.655 2057.180 ;
        RECT 1990.025 2057.175 1990.355 2057.180 ;
        RECT 2004.745 2057.175 2005.075 2057.180 ;
        RECT 2016.245 2057.175 2016.575 2057.180 ;
        RECT 2008.425 2056.820 2008.755 2056.825 ;
        RECT 2021.765 2056.820 2022.095 2056.825 ;
        RECT 2008.425 2056.810 2009.010 2056.820 ;
      LAYER met3 ;
        RECT 300.065 2055.240 1395.600 2056.640 ;
      LAYER met3 ;
        RECT 2008.200 2056.510 2009.010 2056.810 ;
        RECT 2008.425 2056.500 2009.010 2056.510 ;
        RECT 2021.510 2056.810 2022.095 2056.820 ;
        RECT 2021.510 2056.510 2022.320 2056.810 ;
        RECT 2021.510 2056.500 2022.095 2056.510 ;
        RECT 2008.425 2056.495 2008.755 2056.500 ;
        RECT 2021.765 2056.495 2022.095 2056.500 ;
        RECT 1396.000 2056.130 1400.000 2056.240 ;
        RECT 1414.105 2056.130 1414.435 2056.145 ;
        RECT 1396.000 2055.830 1414.435 2056.130 ;
        RECT 1396.000 2055.640 1400.000 2055.830 ;
        RECT 1414.105 2055.815 1414.435 2055.830 ;
        RECT 1948.625 2055.460 1948.955 2055.465 ;
        RECT 1948.625 2055.450 1949.210 2055.460 ;
      LAYER met3 ;
        RECT 300.065 2051.880 1396.000 2055.240 ;
      LAYER met3 ;
        RECT 1948.400 2055.150 1949.210 2055.450 ;
        RECT 1948.625 2055.140 1949.210 2055.150 ;
        RECT 1948.625 2055.135 1948.955 2055.140 ;
        RECT 1961.505 2052.060 1961.835 2052.065 ;
        RECT 2049.825 2052.060 2050.155 2052.065 ;
        RECT 1961.480 2052.050 1961.860 2052.060 ;
        RECT 2049.825 2052.050 2050.410 2052.060 ;
      LAYER met3 ;
        RECT 300.065 2050.480 1395.600 2051.880 ;
      LAYER met3 ;
        RECT 1961.050 2051.750 1961.860 2052.050 ;
        RECT 2049.600 2051.750 2050.410 2052.050 ;
        RECT 1961.480 2051.740 1961.860 2051.750 ;
        RECT 2049.825 2051.740 2050.410 2051.750 ;
        RECT 1961.505 2051.735 1961.835 2051.740 ;
        RECT 2049.825 2051.735 2050.155 2051.740 ;
        RECT 1396.000 2051.370 1400.000 2051.480 ;
        RECT 1409.505 2051.370 1409.835 2051.385 ;
        RECT 1396.000 2051.070 1409.835 2051.370 ;
        RECT 1396.000 2050.880 1400.000 2051.070 ;
        RECT 1409.505 2051.055 1409.835 2051.070 ;
      LAYER met3 ;
        RECT 300.065 2049.160 1396.000 2050.480 ;
        RECT 304.400 2047.760 1396.000 2049.160 ;
        RECT 300.065 2047.120 1396.000 2047.760 ;
        RECT 300.065 2045.720 1395.600 2047.120 ;
      LAYER met3 ;
        RECT 1396.000 2046.610 1400.000 2046.720 ;
        RECT 1415.025 2046.610 1415.355 2046.625 ;
        RECT 1396.000 2046.310 1415.355 2046.610 ;
        RECT 1396.000 2046.120 1400.000 2046.310 ;
        RECT 1415.025 2046.295 1415.355 2046.310 ;
      LAYER met3 ;
        RECT 300.065 2041.680 1396.000 2045.720 ;
      LAYER met3 ;
        RECT 1414.565 2042.530 1414.895 2042.545 ;
        RECT 1399.630 2042.230 1414.895 2042.530 ;
      LAYER met3 ;
        RECT 300.065 2040.280 1395.600 2041.680 ;
      LAYER met3 ;
        RECT 1399.630 2041.280 1399.930 2042.230 ;
        RECT 1414.565 2042.215 1414.895 2042.230 ;
        RECT 1396.000 2040.680 1400.000 2041.280 ;
      LAYER met3 ;
        RECT 300.065 2039.640 1396.000 2040.280 ;
      LAYER met3 ;
        RECT 1412.265 2039.810 1412.595 2039.825 ;
      LAYER met3 ;
        RECT 304.400 2038.240 1396.000 2039.640 ;
        RECT 300.065 2036.920 1396.000 2038.240 ;
      LAYER met3 ;
        RECT 1399.630 2039.510 1412.595 2039.810 ;
      LAYER met3 ;
        RECT 300.065 2035.520 1395.600 2036.920 ;
      LAYER met3 ;
        RECT 1399.630 2036.520 1399.930 2039.510 ;
        RECT 1412.265 2039.495 1412.595 2039.510 ;
        RECT 1396.000 2035.920 1400.000 2036.520 ;
      LAYER met3 ;
        RECT 300.065 2031.480 1396.000 2035.520 ;
        RECT 300.065 2030.120 1395.600 2031.480 ;
      LAYER met3 ;
        RECT 1396.000 2030.970 1400.000 2031.080 ;
        RECT 1409.045 2030.970 1409.375 2030.985 ;
        RECT 1396.000 2030.670 1409.375 2030.970 ;
        RECT 1396.000 2030.480 1400.000 2030.670 ;
        RECT 1409.045 2030.655 1409.375 2030.670 ;
      LAYER met3 ;
        RECT 304.400 2030.080 1395.600 2030.120 ;
        RECT 304.400 2028.720 1396.000 2030.080 ;
        RECT 300.065 2026.720 1396.000 2028.720 ;
        RECT 300.065 2025.320 1395.600 2026.720 ;
      LAYER met3 ;
        RECT 1396.000 2026.210 1400.000 2026.320 ;
        RECT 1408.585 2026.210 1408.915 2026.225 ;
        RECT 1396.000 2025.910 1408.915 2026.210 ;
        RECT 1396.000 2025.720 1400.000 2025.910 ;
        RECT 1408.585 2025.895 1408.915 2025.910 ;
      LAYER met3 ;
        RECT 300.065 2021.960 1396.000 2025.320 ;
        RECT 300.065 2020.600 1395.600 2021.960 ;
      LAYER met3 ;
        RECT 1396.000 2021.450 1400.000 2021.560 ;
        RECT 1414.105 2021.450 1414.435 2021.465 ;
        RECT 1396.000 2021.150 1414.435 2021.450 ;
        RECT 1396.000 2020.960 1400.000 2021.150 ;
        RECT 1414.105 2021.135 1414.435 2021.150 ;
      LAYER met3 ;
        RECT 304.400 2020.560 1395.600 2020.600 ;
        RECT 304.400 2019.200 1396.000 2020.560 ;
        RECT 300.065 2016.520 1396.000 2019.200 ;
        RECT 300.065 2015.120 1395.600 2016.520 ;
      LAYER met3 ;
        RECT 1396.000 2016.010 1400.000 2016.120 ;
        RECT 1409.505 2016.010 1409.835 2016.025 ;
        RECT 1396.000 2015.710 1409.835 2016.010 ;
        RECT 1396.000 2015.520 1400.000 2015.710 ;
        RECT 1409.505 2015.695 1409.835 2015.710 ;
      LAYER met3 ;
        RECT 300.065 2011.760 1396.000 2015.120 ;
        RECT 300.065 2011.080 1395.600 2011.760 ;
        RECT 304.400 2010.360 1395.600 2011.080 ;
      LAYER met3 ;
        RECT 1396.000 2011.250 1400.000 2011.360 ;
        RECT 1410.885 2011.250 1411.215 2011.265 ;
        RECT 1396.000 2010.950 1411.215 2011.250 ;
        RECT 1396.000 2010.760 1400.000 2010.950 ;
        RECT 1410.885 2010.935 1411.215 2010.950 ;
      LAYER met3 ;
        RECT 304.400 2009.680 1396.000 2010.360 ;
        RECT 300.065 2006.320 1396.000 2009.680 ;
        RECT 300.065 2004.920 1395.600 2006.320 ;
      LAYER met3 ;
        RECT 1396.000 2005.810 1400.000 2005.920 ;
        RECT 1408.125 2005.810 1408.455 2005.825 ;
        RECT 1396.000 2005.510 1408.455 2005.810 ;
        RECT 1396.000 2005.320 1400.000 2005.510 ;
        RECT 1408.125 2005.495 1408.455 2005.510 ;
      LAYER met3 ;
        RECT 300.065 2001.560 1396.000 2004.920 ;
        RECT 300.065 2000.880 1395.600 2001.560 ;
        RECT 304.400 2000.160 1395.600 2000.880 ;
      LAYER met3 ;
        RECT 1396.000 2001.050 1400.000 2001.160 ;
        RECT 1408.125 2001.050 1408.455 2001.065 ;
        RECT 1396.000 2000.750 1408.455 2001.050 ;
        RECT 1396.000 2000.560 1400.000 2000.750 ;
        RECT 1408.125 2000.735 1408.455 2000.750 ;
      LAYER met3 ;
        RECT 304.400 1999.480 1396.000 2000.160 ;
        RECT 300.065 1996.120 1396.000 1999.480 ;
        RECT 300.065 1994.720 1395.600 1996.120 ;
      LAYER met3 ;
        RECT 1396.000 1995.610 1400.000 1995.720 ;
        RECT 1408.125 1995.610 1408.455 1995.625 ;
        RECT 1396.000 1995.310 1408.455 1995.610 ;
        RECT 1396.000 1995.120 1400.000 1995.310 ;
        RECT 1408.125 1995.295 1408.455 1995.310 ;
      LAYER met3 ;
        RECT 300.065 1991.360 1396.000 1994.720 ;
        RECT 304.400 1989.960 1395.600 1991.360 ;
      LAYER met3 ;
        RECT 1396.000 1990.850 1400.000 1990.960 ;
        RECT 1410.885 1990.850 1411.215 1990.865 ;
        RECT 1396.000 1990.550 1411.215 1990.850 ;
        RECT 1396.000 1990.360 1400.000 1990.550 ;
        RECT 1410.885 1990.535 1411.215 1990.550 ;
      LAYER met3 ;
        RECT 300.065 1986.600 1396.000 1989.960 ;
        RECT 300.065 1985.200 1395.600 1986.600 ;
      LAYER met3 ;
        RECT 1396.000 1986.090 1400.000 1986.200 ;
        RECT 1417.990 1986.090 1418.370 1986.100 ;
        RECT 1396.000 1985.790 1418.370 1986.090 ;
        RECT 1396.000 1985.600 1400.000 1985.790 ;
        RECT 1417.990 1985.780 1418.370 1985.790 ;
      LAYER met3 ;
        RECT 300.065 1981.840 1396.000 1985.200 ;
        RECT 304.400 1981.160 1396.000 1981.840 ;
        RECT 304.400 1980.440 1395.600 1981.160 ;
        RECT 300.065 1979.760 1395.600 1980.440 ;
      LAYER met3 ;
        RECT 1396.000 1980.650 1400.000 1980.760 ;
        RECT 1418.910 1980.650 1419.290 1980.660 ;
        RECT 1396.000 1980.350 1419.290 1980.650 ;
        RECT 1396.000 1980.160 1400.000 1980.350 ;
        RECT 1418.910 1980.340 1419.290 1980.350 ;
      LAYER met3 ;
        RECT 300.065 1976.400 1396.000 1979.760 ;
        RECT 300.065 1975.000 1395.600 1976.400 ;
      LAYER met3 ;
        RECT 1396.000 1975.890 1400.000 1976.000 ;
        RECT 1417.070 1975.890 1417.450 1975.900 ;
        RECT 1396.000 1975.590 1417.450 1975.890 ;
        RECT 1396.000 1975.400 1400.000 1975.590 ;
        RECT 1417.070 1975.580 1417.450 1975.590 ;
      LAYER met3 ;
        RECT 300.065 1972.320 1396.000 1975.000 ;
        RECT 304.400 1970.960 1396.000 1972.320 ;
        RECT 304.400 1970.920 1395.600 1970.960 ;
        RECT 300.065 1969.560 1395.600 1970.920 ;
      LAYER met3 ;
        RECT 1396.000 1970.450 1400.000 1970.560 ;
        RECT 1408.125 1970.450 1408.455 1970.465 ;
        RECT 1396.000 1970.150 1408.455 1970.450 ;
        RECT 1396.000 1969.960 1400.000 1970.150 ;
        RECT 1408.125 1970.135 1408.455 1970.150 ;
      LAYER met3 ;
        RECT 300.065 1966.200 1396.000 1969.560 ;
      LAYER met3 ;
        RECT 1408.585 1966.370 1408.915 1966.385 ;
        RECT 1412.265 1966.370 1412.595 1966.385 ;
      LAYER met3 ;
        RECT 300.065 1964.800 1395.600 1966.200 ;
      LAYER met3 ;
        RECT 1408.585 1966.070 1412.595 1966.370 ;
        RECT 1408.585 1966.055 1408.915 1966.070 ;
        RECT 1412.265 1966.055 1412.595 1966.070 ;
        RECT 1396.000 1965.690 1400.000 1965.800 ;
        RECT 1408.125 1965.690 1408.455 1965.705 ;
        RECT 1396.000 1965.390 1408.455 1965.690 ;
        RECT 1396.000 1965.200 1400.000 1965.390 ;
        RECT 1408.125 1965.375 1408.455 1965.390 ;
      LAYER met3 ;
        RECT 300.065 1962.800 1396.000 1964.800 ;
        RECT 304.400 1961.400 1396.000 1962.800 ;
        RECT 300.065 1960.760 1396.000 1961.400 ;
        RECT 300.065 1959.360 1395.600 1960.760 ;
      LAYER met3 ;
        RECT 1396.000 1960.250 1400.000 1960.360 ;
        RECT 1408.125 1960.250 1408.455 1960.265 ;
        RECT 1396.000 1959.950 1408.455 1960.250 ;
        RECT 1396.000 1959.760 1400.000 1959.950 ;
        RECT 1408.125 1959.935 1408.455 1959.950 ;
      LAYER met3 ;
        RECT 300.065 1956.000 1396.000 1959.360 ;
        RECT 300.065 1954.600 1395.600 1956.000 ;
      LAYER met3 ;
        RECT 1396.000 1955.490 1400.000 1955.600 ;
        RECT 1411.550 1955.490 1411.930 1955.500 ;
        RECT 1396.000 1955.190 1411.930 1955.490 ;
        RECT 1396.000 1955.000 1400.000 1955.190 ;
        RECT 1411.550 1955.180 1411.930 1955.190 ;
      LAYER met3 ;
        RECT 300.065 1952.600 1396.000 1954.600 ;
        RECT 304.400 1951.240 1396.000 1952.600 ;
      LAYER met3 ;
        RECT 1700.000 1951.445 1704.600 1951.745 ;
      LAYER met3 ;
        RECT 304.400 1951.200 1395.600 1951.240 ;
        RECT 300.065 1949.840 1395.600 1951.200 ;
      LAYER met3 ;
        RECT 1396.000 1950.730 1400.000 1950.840 ;
        RECT 1409.505 1950.730 1409.835 1950.745 ;
        RECT 1396.000 1950.430 1409.835 1950.730 ;
        RECT 1396.000 1950.240 1400.000 1950.430 ;
        RECT 1409.505 1950.415 1409.835 1950.430 ;
      LAYER met3 ;
        RECT 300.065 1945.800 1396.000 1949.840 ;
      LAYER met3 ;
        RECT 1690.105 1949.370 1690.435 1949.385 ;
        RECT 1700.470 1949.370 1700.770 1951.445 ;
        RECT 1690.105 1949.070 1700.770 1949.370 ;
        RECT 1690.105 1949.055 1690.435 1949.070 ;
        RECT 1700.470 1946.105 1700.770 1949.070 ;
        RECT 1700.000 1945.805 1704.600 1946.105 ;
      LAYER met3 ;
        RECT 300.065 1944.400 1395.600 1945.800 ;
      LAYER met3 ;
        RECT 1396.000 1945.290 1400.000 1945.400 ;
        RECT 1414.105 1945.290 1414.435 1945.305 ;
        RECT 1396.000 1944.990 1414.435 1945.290 ;
        RECT 1396.000 1944.800 1400.000 1944.990 ;
        RECT 1414.105 1944.975 1414.435 1944.990 ;
      LAYER met3 ;
        RECT 300.065 1943.080 1396.000 1944.400 ;
        RECT 304.400 1941.680 1396.000 1943.080 ;
        RECT 300.065 1941.040 1396.000 1941.680 ;
        RECT 300.065 1939.640 1395.600 1941.040 ;
      LAYER met3 ;
        RECT 1396.000 1940.530 1400.000 1940.640 ;
        RECT 1408.125 1940.530 1408.455 1940.545 ;
        RECT 1396.000 1940.230 1408.455 1940.530 ;
        RECT 1396.000 1940.040 1400.000 1940.230 ;
        RECT 1408.125 1940.215 1408.455 1940.230 ;
      LAYER met3 ;
        RECT 300.065 1935.600 1396.000 1939.640 ;
      LAYER met3 ;
        RECT 1700.470 1937.605 1700.770 1945.805 ;
        RECT 1700.000 1937.305 1704.600 1937.605 ;
      LAYER met3 ;
        RECT 300.065 1934.200 1395.600 1935.600 ;
      LAYER met3 ;
        RECT 1396.000 1935.090 1400.000 1935.200 ;
        RECT 1408.125 1935.090 1408.455 1935.105 ;
        RECT 1396.000 1934.790 1408.455 1935.090 ;
        RECT 1396.000 1934.600 1400.000 1934.790 ;
        RECT 1408.125 1934.775 1408.455 1934.790 ;
      LAYER met3 ;
        RECT 300.065 1933.560 1396.000 1934.200 ;
        RECT 304.400 1932.160 1396.000 1933.560 ;
        RECT 300.065 1930.840 1396.000 1932.160 ;
      LAYER met3 ;
        RECT 1700.470 1931.965 1700.770 1937.305 ;
        RECT 1700.000 1931.665 1704.600 1931.965 ;
      LAYER met3 ;
        RECT 300.065 1929.440 1395.600 1930.840 ;
      LAYER met3 ;
        RECT 1396.000 1930.330 1400.000 1930.440 ;
        RECT 1408.585 1930.330 1408.915 1930.345 ;
        RECT 1396.000 1930.030 1408.915 1930.330 ;
        RECT 1396.000 1929.840 1400.000 1930.030 ;
        RECT 1408.585 1930.015 1408.915 1930.030 ;
      LAYER met3 ;
        RECT 300.065 1926.080 1396.000 1929.440 ;
        RECT 300.065 1924.680 1395.600 1926.080 ;
      LAYER met3 ;
        RECT 1396.000 1925.570 1400.000 1925.680 ;
        RECT 1408.125 1925.570 1408.455 1925.585 ;
        RECT 1396.000 1925.270 1408.455 1925.570 ;
        RECT 1396.000 1925.080 1400.000 1925.270 ;
        RECT 1408.125 1925.255 1408.455 1925.270 ;
      LAYER met3 ;
        RECT 300.065 1924.040 1396.000 1924.680 ;
        RECT 304.400 1922.640 1396.000 1924.040 ;
      LAYER met3 ;
        RECT 1700.470 1923.465 1700.770 1931.665 ;
        RECT 1700.000 1923.165 1704.600 1923.465 ;
      LAYER met3 ;
        RECT 300.065 1920.640 1396.000 1922.640 ;
        RECT 300.065 1919.240 1395.600 1920.640 ;
      LAYER met3 ;
        RECT 1396.000 1920.130 1400.000 1920.240 ;
        RECT 1408.125 1920.130 1408.455 1920.145 ;
        RECT 1396.000 1919.830 1408.455 1920.130 ;
        RECT 1396.000 1919.640 1400.000 1919.830 ;
        RECT 1408.125 1919.815 1408.455 1919.830 ;
      LAYER met3 ;
        RECT 300.065 1915.880 1396.000 1919.240 ;
      LAYER met3 ;
        RECT 1700.470 1917.825 1700.770 1923.165 ;
        RECT 1700.000 1917.525 1704.600 1917.825 ;
      LAYER met3 ;
        RECT 300.065 1914.520 1395.600 1915.880 ;
      LAYER met3 ;
        RECT 1396.000 1915.370 1400.000 1915.480 ;
        RECT 1414.105 1915.370 1414.435 1915.385 ;
        RECT 1396.000 1915.070 1414.435 1915.370 ;
        RECT 1396.000 1914.880 1400.000 1915.070 ;
        RECT 1414.105 1915.055 1414.435 1915.070 ;
      LAYER met3 ;
        RECT 304.400 1914.480 1395.600 1914.520 ;
        RECT 304.400 1913.120 1396.000 1914.480 ;
        RECT 300.065 1910.440 1396.000 1913.120 ;
        RECT 300.065 1909.040 1395.600 1910.440 ;
      LAYER met3 ;
        RECT 1396.000 1909.930 1400.000 1910.040 ;
        RECT 1408.125 1909.930 1408.455 1909.945 ;
        RECT 1396.000 1909.630 1408.455 1909.930 ;
        RECT 1396.000 1909.440 1400.000 1909.630 ;
        RECT 1408.125 1909.615 1408.455 1909.630 ;
        RECT 1700.470 1909.325 1700.770 1917.525 ;
      LAYER met3 ;
        RECT 300.065 1905.680 1396.000 1909.040 ;
      LAYER met3 ;
        RECT 1700.000 1909.025 1704.600 1909.325 ;
        RECT 1686.885 1906.530 1687.215 1906.545 ;
        RECT 1700.470 1906.530 1700.770 1909.025 ;
        RECT 1686.885 1906.230 1700.770 1906.530 ;
        RECT 1686.885 1906.215 1687.215 1906.230 ;
      LAYER met3 ;
        RECT 300.065 1904.320 1395.600 1905.680 ;
      LAYER met3 ;
        RECT 1396.000 1905.170 1400.000 1905.280 ;
        RECT 1408.585 1905.170 1408.915 1905.185 ;
        RECT 1396.000 1904.870 1408.915 1905.170 ;
        RECT 1396.000 1904.680 1400.000 1904.870 ;
        RECT 1408.585 1904.855 1408.915 1904.870 ;
      LAYER met3 ;
        RECT 304.400 1904.280 1395.600 1904.320 ;
        RECT 304.400 1902.920 1396.000 1904.280 ;
        RECT 300.065 1900.240 1396.000 1902.920 ;
        RECT 300.065 1898.840 1395.600 1900.240 ;
      LAYER met3 ;
        RECT 1396.000 1899.730 1400.000 1899.840 ;
        RECT 1414.105 1899.730 1414.435 1899.745 ;
        RECT 1396.000 1899.430 1414.435 1899.730 ;
        RECT 1396.000 1899.240 1400.000 1899.430 ;
        RECT 1414.105 1899.415 1414.435 1899.430 ;
      LAYER met3 ;
        RECT 300.065 1895.480 1396.000 1898.840 ;
        RECT 300.065 1894.800 1395.600 1895.480 ;
        RECT 304.400 1894.080 1395.600 1894.800 ;
      LAYER met3 ;
        RECT 1396.000 1894.970 1400.000 1895.080 ;
        RECT 1414.105 1894.970 1414.435 1894.985 ;
        RECT 1396.000 1894.670 1414.435 1894.970 ;
        RECT 1396.000 1894.480 1400.000 1894.670 ;
        RECT 1414.105 1894.655 1414.435 1894.670 ;
      LAYER met3 ;
        RECT 304.400 1893.400 1396.000 1894.080 ;
        RECT 300.065 1890.720 1396.000 1893.400 ;
        RECT 300.065 1889.320 1395.600 1890.720 ;
      LAYER met3 ;
        RECT 1396.000 1890.210 1400.000 1890.320 ;
        RECT 1414.105 1890.210 1414.435 1890.225 ;
        RECT 1396.000 1889.910 1414.435 1890.210 ;
        RECT 1396.000 1889.720 1400.000 1889.910 ;
        RECT 1414.105 1889.895 1414.435 1889.910 ;
      LAYER met3 ;
        RECT 300.065 1885.280 1396.000 1889.320 ;
        RECT 304.400 1883.880 1395.600 1885.280 ;
      LAYER met3 ;
        RECT 1396.000 1884.770 1400.000 1884.880 ;
        RECT 1410.885 1884.770 1411.215 1884.785 ;
        RECT 1396.000 1884.470 1411.215 1884.770 ;
        RECT 1396.000 1884.280 1400.000 1884.470 ;
        RECT 1410.885 1884.455 1411.215 1884.470 ;
      LAYER met3 ;
        RECT 300.065 1880.520 1396.000 1883.880 ;
        RECT 300.065 1879.120 1395.600 1880.520 ;
      LAYER met3 ;
        RECT 1396.000 1880.010 1400.000 1880.120 ;
        RECT 1414.105 1880.010 1414.435 1880.025 ;
        RECT 1396.000 1879.710 1414.435 1880.010 ;
        RECT 1396.000 1879.520 1400.000 1879.710 ;
        RECT 1414.105 1879.695 1414.435 1879.710 ;
      LAYER met3 ;
        RECT 300.065 1875.760 1396.000 1879.120 ;
        RECT 304.400 1875.080 1396.000 1875.760 ;
        RECT 304.400 1874.360 1395.600 1875.080 ;
        RECT 300.065 1873.680 1395.600 1874.360 ;
      LAYER met3 ;
        RECT 1396.000 1874.570 1400.000 1874.680 ;
        RECT 1414.105 1874.570 1414.435 1874.585 ;
        RECT 1396.000 1874.270 1414.435 1874.570 ;
        RECT 1396.000 1874.080 1400.000 1874.270 ;
        RECT 1414.105 1874.255 1414.435 1874.270 ;
      LAYER met3 ;
        RECT 300.065 1870.320 1396.000 1873.680 ;
        RECT 300.065 1868.920 1395.600 1870.320 ;
      LAYER met3 ;
        RECT 1396.000 1869.810 1400.000 1869.920 ;
        RECT 1414.105 1869.810 1414.435 1869.825 ;
        RECT 1396.000 1869.510 1414.435 1869.810 ;
        RECT 1396.000 1869.320 1400.000 1869.510 ;
        RECT 1414.105 1869.495 1414.435 1869.510 ;
      LAYER met3 ;
        RECT 300.065 1866.240 1396.000 1868.920 ;
        RECT 304.400 1864.880 1396.000 1866.240 ;
        RECT 304.400 1864.840 1395.600 1864.880 ;
        RECT 300.065 1863.480 1395.600 1864.840 ;
      LAYER met3 ;
        RECT 1396.000 1864.370 1400.000 1864.480 ;
        RECT 1410.885 1864.370 1411.215 1864.385 ;
        RECT 1396.000 1864.070 1411.215 1864.370 ;
        RECT 1396.000 1863.880 1400.000 1864.070 ;
        RECT 1410.885 1864.055 1411.215 1864.070 ;
      LAYER met3 ;
        RECT 300.065 1860.120 1396.000 1863.480 ;
        RECT 300.065 1858.720 1395.600 1860.120 ;
      LAYER met3 ;
        RECT 1396.000 1859.610 1400.000 1859.720 ;
        RECT 1414.105 1859.610 1414.435 1859.625 ;
        RECT 1396.000 1859.310 1414.435 1859.610 ;
        RECT 1396.000 1859.120 1400.000 1859.310 ;
        RECT 1414.105 1859.295 1414.435 1859.310 ;
      LAYER met3 ;
        RECT 300.065 1856.720 1396.000 1858.720 ;
        RECT 304.400 1855.360 1396.000 1856.720 ;
        RECT 304.400 1855.320 1395.600 1855.360 ;
        RECT 300.065 1853.960 1395.600 1855.320 ;
      LAYER met3 ;
        RECT 1396.000 1854.850 1400.000 1854.960 ;
        RECT 1414.105 1854.850 1414.435 1854.865 ;
        RECT 1396.000 1854.550 1414.435 1854.850 ;
        RECT 1396.000 1854.360 1400.000 1854.550 ;
        RECT 1414.105 1854.535 1414.435 1854.550 ;
      LAYER met3 ;
        RECT 300.065 1849.920 1396.000 1853.960 ;
        RECT 300.065 1848.520 1395.600 1849.920 ;
      LAYER met3 ;
        RECT 1396.000 1849.410 1400.000 1849.520 ;
        RECT 1410.885 1849.410 1411.215 1849.425 ;
        RECT 1396.000 1849.110 1411.215 1849.410 ;
        RECT 1396.000 1848.920 1400.000 1849.110 ;
        RECT 1410.885 1849.095 1411.215 1849.110 ;
      LAYER met3 ;
        RECT 300.065 1846.520 1396.000 1848.520 ;
        RECT 304.400 1845.160 1396.000 1846.520 ;
        RECT 304.400 1845.120 1395.600 1845.160 ;
        RECT 300.065 1843.760 1395.600 1845.120 ;
      LAYER met3 ;
        RECT 1396.000 1844.650 1400.000 1844.760 ;
        RECT 1414.105 1844.650 1414.435 1844.665 ;
        RECT 1396.000 1844.350 1414.435 1844.650 ;
        RECT 1396.000 1844.160 1400.000 1844.350 ;
        RECT 1414.105 1844.335 1414.435 1844.350 ;
      LAYER met3 ;
        RECT 300.065 1839.720 1396.000 1843.760 ;
        RECT 300.065 1838.320 1395.600 1839.720 ;
      LAYER met3 ;
        RECT 1396.000 1839.210 1400.000 1839.320 ;
        RECT 1414.105 1839.210 1414.435 1839.225 ;
        RECT 1396.000 1838.910 1414.435 1839.210 ;
        RECT 1396.000 1838.720 1400.000 1838.910 ;
        RECT 1414.105 1838.895 1414.435 1838.910 ;
      LAYER met3 ;
        RECT 300.065 1837.000 1396.000 1838.320 ;
        RECT 304.400 1835.600 1396.000 1837.000 ;
        RECT 300.065 1834.960 1396.000 1835.600 ;
        RECT 300.065 1833.560 1395.600 1834.960 ;
      LAYER met3 ;
        RECT 1396.000 1834.450 1400.000 1834.560 ;
        RECT 1414.105 1834.450 1414.435 1834.465 ;
        RECT 1396.000 1834.150 1414.435 1834.450 ;
        RECT 1396.000 1833.960 1400.000 1834.150 ;
        RECT 1414.105 1834.135 1414.435 1834.150 ;
      LAYER met3 ;
        RECT 300.065 1829.520 1396.000 1833.560 ;
        RECT 300.065 1828.120 1395.600 1829.520 ;
      LAYER met3 ;
        RECT 1396.000 1829.010 1400.000 1829.120 ;
        RECT 1410.885 1829.010 1411.215 1829.025 ;
        RECT 1396.000 1828.710 1411.215 1829.010 ;
        RECT 1396.000 1828.520 1400.000 1828.710 ;
        RECT 1410.885 1828.695 1411.215 1828.710 ;
      LAYER met3 ;
        RECT 300.065 1827.480 1396.000 1828.120 ;
        RECT 304.400 1826.080 1396.000 1827.480 ;
        RECT 300.065 1824.760 1396.000 1826.080 ;
        RECT 300.065 1823.360 1395.600 1824.760 ;
      LAYER met3 ;
        RECT 1396.000 1824.250 1400.000 1824.360 ;
        RECT 1414.105 1824.250 1414.435 1824.265 ;
        RECT 1396.000 1823.950 1414.435 1824.250 ;
        RECT 1396.000 1823.760 1400.000 1823.950 ;
        RECT 1414.105 1823.935 1414.435 1823.950 ;
      LAYER met3 ;
        RECT 300.065 1820.000 1396.000 1823.360 ;
        RECT 300.065 1818.600 1395.600 1820.000 ;
      LAYER met3 ;
        RECT 1396.000 1819.490 1400.000 1819.600 ;
        RECT 1414.105 1819.490 1414.435 1819.505 ;
        RECT 1396.000 1819.190 1414.435 1819.490 ;
        RECT 1396.000 1819.000 1400.000 1819.190 ;
        RECT 1414.105 1819.175 1414.435 1819.190 ;
      LAYER met3 ;
        RECT 300.065 1817.960 1396.000 1818.600 ;
        RECT 304.400 1816.560 1396.000 1817.960 ;
        RECT 300.065 1814.560 1396.000 1816.560 ;
        RECT 300.065 1813.160 1395.600 1814.560 ;
      LAYER met3 ;
        RECT 1396.000 1814.050 1400.000 1814.160 ;
        RECT 1414.105 1814.050 1414.435 1814.065 ;
        RECT 1396.000 1813.750 1414.435 1814.050 ;
        RECT 1396.000 1813.560 1400.000 1813.750 ;
        RECT 1414.105 1813.735 1414.435 1813.750 ;
      LAYER met3 ;
        RECT 300.065 1809.800 1396.000 1813.160 ;
        RECT 300.065 1808.440 1395.600 1809.800 ;
      LAYER met3 ;
        RECT 1396.000 1809.290 1400.000 1809.400 ;
        RECT 1413.645 1809.290 1413.975 1809.305 ;
        RECT 1396.000 1808.990 1413.975 1809.290 ;
        RECT 1396.000 1808.800 1400.000 1808.990 ;
        RECT 1413.645 1808.975 1413.975 1808.990 ;
      LAYER met3 ;
        RECT 304.400 1808.400 1395.600 1808.440 ;
        RECT 304.400 1807.040 1396.000 1808.400 ;
        RECT 300.065 1804.360 1396.000 1807.040 ;
        RECT 300.065 1802.960 1395.600 1804.360 ;
      LAYER met3 ;
        RECT 1396.000 1803.850 1400.000 1803.960 ;
        RECT 1408.585 1803.850 1408.915 1803.865 ;
        RECT 1396.000 1803.550 1408.915 1803.850 ;
        RECT 1396.000 1803.360 1400.000 1803.550 ;
        RECT 1408.585 1803.535 1408.915 1803.550 ;
      LAYER met3 ;
        RECT 300.065 1799.600 1396.000 1802.960 ;
        RECT 300.065 1798.240 1395.600 1799.600 ;
      LAYER met3 ;
        RECT 1396.000 1799.090 1400.000 1799.200 ;
        RECT 1414.105 1799.090 1414.435 1799.105 ;
        RECT 1396.000 1798.790 1414.435 1799.090 ;
        RECT 1396.000 1798.600 1400.000 1798.790 ;
        RECT 1414.105 1798.775 1414.435 1798.790 ;
      LAYER met3 ;
        RECT 304.400 1798.200 1395.600 1798.240 ;
        RECT 304.400 1796.840 1396.000 1798.200 ;
        RECT 300.065 1794.840 1396.000 1796.840 ;
        RECT 300.065 1793.440 1395.600 1794.840 ;
      LAYER met3 ;
        RECT 1396.000 1794.330 1400.000 1794.440 ;
        RECT 1413.645 1794.330 1413.975 1794.345 ;
        RECT 1396.000 1794.030 1413.975 1794.330 ;
        RECT 1396.000 1793.840 1400.000 1794.030 ;
        RECT 1413.645 1794.015 1413.975 1794.030 ;
      LAYER met3 ;
        RECT 300.065 1789.400 1396.000 1793.440 ;
        RECT 300.065 1788.720 1395.600 1789.400 ;
        RECT 304.400 1788.000 1395.600 1788.720 ;
      LAYER met3 ;
        RECT 1396.000 1788.890 1400.000 1789.000 ;
        RECT 1409.505 1788.890 1409.835 1788.905 ;
        RECT 1396.000 1788.590 1409.835 1788.890 ;
        RECT 1396.000 1788.400 1400.000 1788.590 ;
        RECT 1409.505 1788.575 1409.835 1788.590 ;
      LAYER met3 ;
        RECT 304.400 1787.320 1396.000 1788.000 ;
        RECT 300.065 1784.640 1396.000 1787.320 ;
        RECT 300.065 1783.240 1395.600 1784.640 ;
      LAYER met3 ;
        RECT 1396.000 1784.130 1400.000 1784.240 ;
        RECT 1409.965 1784.130 1410.295 1784.145 ;
        RECT 1396.000 1783.830 1410.295 1784.130 ;
        RECT 1396.000 1783.640 1400.000 1783.830 ;
        RECT 1409.965 1783.815 1410.295 1783.830 ;
      LAYER met3 ;
        RECT 300.065 1779.200 1396.000 1783.240 ;
        RECT 304.400 1777.800 1395.600 1779.200 ;
      LAYER met3 ;
        RECT 1396.000 1778.690 1400.000 1778.800 ;
        RECT 1410.425 1778.690 1410.755 1778.705 ;
        RECT 1396.000 1778.390 1410.755 1778.690 ;
        RECT 1396.000 1778.200 1400.000 1778.390 ;
        RECT 1410.425 1778.375 1410.755 1778.390 ;
      LAYER met3 ;
        RECT 300.065 1774.440 1396.000 1777.800 ;
        RECT 300.065 1773.040 1395.600 1774.440 ;
      LAYER met3 ;
        RECT 1396.000 1773.930 1400.000 1774.040 ;
        RECT 1410.885 1773.930 1411.215 1773.945 ;
        RECT 1396.000 1773.630 1411.215 1773.930 ;
        RECT 1396.000 1773.440 1400.000 1773.630 ;
        RECT 1410.885 1773.615 1411.215 1773.630 ;
        RECT 1409.965 1773.250 1410.295 1773.265 ;
        RECT 1411.805 1773.250 1412.135 1773.265 ;
      LAYER met3 ;
        RECT 300.065 1769.680 1396.000 1773.040 ;
      LAYER met3 ;
        RECT 1409.965 1772.950 1412.135 1773.250 ;
        RECT 1409.965 1772.935 1410.295 1772.950 ;
        RECT 1411.805 1772.935 1412.135 1772.950 ;
      LAYER met3 ;
        RECT 304.400 1769.000 1396.000 1769.680 ;
        RECT 304.400 1768.280 1395.600 1769.000 ;
        RECT 300.065 1767.600 1395.600 1768.280 ;
      LAYER met3 ;
        RECT 1396.000 1768.490 1400.000 1768.600 ;
        RECT 1413.185 1768.490 1413.515 1768.505 ;
        RECT 1396.000 1768.190 1413.515 1768.490 ;
        RECT 1396.000 1768.000 1400.000 1768.190 ;
        RECT 1413.185 1768.175 1413.515 1768.190 ;
      LAYER met3 ;
        RECT 300.065 1764.240 1396.000 1767.600 ;
        RECT 300.065 1762.840 1395.600 1764.240 ;
      LAYER met3 ;
        RECT 1396.000 1763.730 1400.000 1763.840 ;
        RECT 1410.425 1763.730 1410.755 1763.745 ;
        RECT 1396.000 1763.430 1410.755 1763.730 ;
        RECT 1396.000 1763.240 1400.000 1763.430 ;
        RECT 1410.425 1763.415 1410.755 1763.430 ;
      LAYER met3 ;
        RECT 300.065 1760.160 1396.000 1762.840 ;
        RECT 304.400 1759.480 1396.000 1760.160 ;
        RECT 304.400 1758.760 1395.600 1759.480 ;
        RECT 300.065 1758.080 1395.600 1758.760 ;
      LAYER met3 ;
        RECT 1396.000 1758.970 1400.000 1759.080 ;
        RECT 1409.965 1758.970 1410.295 1758.985 ;
        RECT 1396.000 1758.670 1410.295 1758.970 ;
        RECT 1396.000 1758.480 1400.000 1758.670 ;
        RECT 1409.965 1758.655 1410.295 1758.670 ;
      LAYER met3 ;
        RECT 300.065 1754.040 1396.000 1758.080 ;
        RECT 300.065 1752.640 1395.600 1754.040 ;
      LAYER met3 ;
        RECT 1396.000 1753.530 1400.000 1753.640 ;
        RECT 1412.725 1753.530 1413.055 1753.545 ;
        RECT 1396.000 1753.230 1413.055 1753.530 ;
        RECT 1396.000 1753.040 1400.000 1753.230 ;
        RECT 1412.725 1753.215 1413.055 1753.230 ;
      LAYER met3 ;
        RECT 300.065 1749.960 1396.000 1752.640 ;
        RECT 304.400 1749.280 1396.000 1749.960 ;
        RECT 304.400 1748.560 1395.600 1749.280 ;
        RECT 300.065 1747.880 1395.600 1748.560 ;
      LAYER met3 ;
        RECT 1396.000 1748.770 1400.000 1748.880 ;
        RECT 1411.345 1748.770 1411.675 1748.785 ;
        RECT 1396.000 1748.470 1411.675 1748.770 ;
        RECT 1396.000 1748.280 1400.000 1748.470 ;
        RECT 1411.345 1748.455 1411.675 1748.470 ;
      LAYER met3 ;
        RECT 300.065 1743.840 1396.000 1747.880 ;
        RECT 300.065 1742.440 1395.600 1743.840 ;
      LAYER met3 ;
        RECT 1396.000 1743.330 1400.000 1743.440 ;
        RECT 1414.105 1743.330 1414.435 1743.345 ;
        RECT 1396.000 1743.030 1414.435 1743.330 ;
        RECT 1396.000 1742.840 1400.000 1743.030 ;
        RECT 1414.105 1743.015 1414.435 1743.030 ;
      LAYER met3 ;
        RECT 300.065 1740.440 1396.000 1742.440 ;
        RECT 304.400 1739.080 1396.000 1740.440 ;
        RECT 304.400 1739.040 1395.600 1739.080 ;
        RECT 300.065 1737.680 1395.600 1739.040 ;
      LAYER met3 ;
        RECT 1396.000 1738.570 1400.000 1738.680 ;
        RECT 1414.105 1738.570 1414.435 1738.585 ;
        RECT 1396.000 1738.270 1414.435 1738.570 ;
        RECT 1396.000 1738.080 1400.000 1738.270 ;
        RECT 1414.105 1738.255 1414.435 1738.270 ;
      LAYER met3 ;
        RECT 300.065 1733.640 1396.000 1737.680 ;
        RECT 300.065 1732.240 1395.600 1733.640 ;
      LAYER met3 ;
        RECT 1396.000 1733.130 1400.000 1733.240 ;
        RECT 1411.345 1733.130 1411.675 1733.145 ;
        RECT 1396.000 1732.830 1411.675 1733.130 ;
        RECT 1396.000 1732.640 1400.000 1732.830 ;
        RECT 1411.345 1732.815 1411.675 1732.830 ;
      LAYER met3 ;
        RECT 300.065 1730.920 1396.000 1732.240 ;
        RECT 304.400 1729.520 1396.000 1730.920 ;
        RECT 300.065 1728.880 1396.000 1729.520 ;
        RECT 300.065 1727.480 1395.600 1728.880 ;
      LAYER met3 ;
        RECT 1396.000 1728.370 1400.000 1728.480 ;
        RECT 1410.425 1728.370 1410.755 1728.385 ;
        RECT 1396.000 1728.070 1410.755 1728.370 ;
        RECT 1396.000 1727.880 1400.000 1728.070 ;
        RECT 1410.425 1728.055 1410.755 1728.070 ;
      LAYER met3 ;
        RECT 300.065 1724.120 1396.000 1727.480 ;
        RECT 300.065 1722.720 1395.600 1724.120 ;
      LAYER met3 ;
        RECT 1396.000 1723.610 1400.000 1723.720 ;
        RECT 1414.105 1723.610 1414.435 1723.625 ;
        RECT 1396.000 1723.310 1414.435 1723.610 ;
        RECT 1396.000 1723.120 1400.000 1723.310 ;
        RECT 1414.105 1723.295 1414.435 1723.310 ;
      LAYER met3 ;
        RECT 300.065 1721.400 1396.000 1722.720 ;
        RECT 304.400 1720.000 1396.000 1721.400 ;
        RECT 300.065 1718.680 1396.000 1720.000 ;
        RECT 300.065 1717.280 1395.600 1718.680 ;
      LAYER met3 ;
        RECT 1396.000 1718.170 1400.000 1718.280 ;
        RECT 1413.645 1718.170 1413.975 1718.185 ;
        RECT 1396.000 1717.870 1413.975 1718.170 ;
        RECT 1396.000 1717.680 1400.000 1717.870 ;
        RECT 1413.645 1717.855 1413.975 1717.870 ;
      LAYER met3 ;
        RECT 300.065 1713.920 1396.000 1717.280 ;
        RECT 300.065 1712.520 1395.600 1713.920 ;
      LAYER met3 ;
        RECT 1396.000 1713.410 1400.000 1713.520 ;
        RECT 1412.725 1713.410 1413.055 1713.425 ;
        RECT 1396.000 1713.110 1413.055 1713.410 ;
        RECT 1396.000 1712.920 1400.000 1713.110 ;
        RECT 1412.725 1713.095 1413.055 1713.110 ;
      LAYER met3 ;
        RECT 300.065 1711.880 1396.000 1712.520 ;
        RECT 304.400 1710.480 1396.000 1711.880 ;
        RECT 300.065 1708.480 1396.000 1710.480 ;
        RECT 300.065 1707.080 1395.600 1708.480 ;
      LAYER met3 ;
        RECT 1396.000 1707.970 1400.000 1708.080 ;
        RECT 1414.105 1707.970 1414.435 1707.985 ;
        RECT 1396.000 1707.670 1414.435 1707.970 ;
        RECT 1396.000 1707.480 1400.000 1707.670 ;
        RECT 1414.105 1707.655 1414.435 1707.670 ;
      LAYER met3 ;
        RECT 300.065 1703.720 1396.000 1707.080 ;
        RECT 300.065 1702.320 1395.600 1703.720 ;
      LAYER met3 ;
        RECT 1396.000 1703.210 1400.000 1703.320 ;
        RECT 1412.265 1703.210 1412.595 1703.225 ;
        RECT 1396.000 1702.910 1412.595 1703.210 ;
        RECT 1396.000 1702.720 1400.000 1702.910 ;
        RECT 1412.265 1702.895 1412.595 1702.910 ;
      LAYER met3 ;
        RECT 300.065 1701.680 1396.000 1702.320 ;
        RECT 304.400 1700.280 1396.000 1701.680 ;
        RECT 300.065 1698.960 1396.000 1700.280 ;
        RECT 300.065 1697.560 1395.600 1698.960 ;
      LAYER met3 ;
        RECT 1396.000 1698.450 1400.000 1698.560 ;
        RECT 1410.425 1698.450 1410.755 1698.465 ;
        RECT 1396.000 1698.150 1410.755 1698.450 ;
        RECT 1396.000 1697.960 1400.000 1698.150 ;
        RECT 1410.425 1698.135 1410.755 1698.150 ;
      LAYER met3 ;
        RECT 300.065 1693.520 1396.000 1697.560 ;
        RECT 300.065 1692.160 1395.600 1693.520 ;
      LAYER met3 ;
        RECT 1396.000 1693.010 1400.000 1693.120 ;
        RECT 1411.805 1693.010 1412.135 1693.025 ;
        RECT 1396.000 1692.710 1412.135 1693.010 ;
        RECT 1396.000 1692.520 1400.000 1692.710 ;
        RECT 1411.805 1692.695 1412.135 1692.710 ;
      LAYER met3 ;
        RECT 304.400 1692.120 1395.600 1692.160 ;
        RECT 304.400 1690.760 1396.000 1692.120 ;
        RECT 300.065 1688.760 1396.000 1690.760 ;
        RECT 300.065 1687.360 1395.600 1688.760 ;
      LAYER met3 ;
        RECT 1396.000 1688.250 1400.000 1688.360 ;
        RECT 1412.725 1688.250 1413.055 1688.265 ;
        RECT 1396.000 1687.950 1413.055 1688.250 ;
        RECT 1396.000 1687.760 1400.000 1687.950 ;
        RECT 1412.725 1687.935 1413.055 1687.950 ;
      LAYER met3 ;
        RECT 300.065 1683.320 1396.000 1687.360 ;
        RECT 300.065 1682.640 1395.600 1683.320 ;
        RECT 304.400 1681.920 1395.600 1682.640 ;
      LAYER met3 ;
        RECT 1396.000 1682.810 1400.000 1682.920 ;
        RECT 1409.965 1682.810 1410.295 1682.825 ;
        RECT 1396.000 1682.510 1410.295 1682.810 ;
        RECT 1396.000 1682.320 1400.000 1682.510 ;
        RECT 1409.965 1682.495 1410.295 1682.510 ;
      LAYER met3 ;
        RECT 304.400 1681.240 1396.000 1681.920 ;
        RECT 300.065 1678.560 1396.000 1681.240 ;
        RECT 300.065 1677.160 1395.600 1678.560 ;
      LAYER met3 ;
        RECT 1396.000 1678.050 1400.000 1678.160 ;
        RECT 1413.185 1678.050 1413.515 1678.065 ;
        RECT 1396.000 1677.750 1413.515 1678.050 ;
        RECT 1396.000 1677.560 1400.000 1677.750 ;
        RECT 1413.185 1677.735 1413.515 1677.750 ;
      LAYER met3 ;
        RECT 300.065 1673.120 1396.000 1677.160 ;
        RECT 304.400 1671.720 1395.600 1673.120 ;
      LAYER met3 ;
        RECT 1396.000 1672.610 1400.000 1672.720 ;
        RECT 1409.045 1672.610 1409.375 1672.625 ;
        RECT 1396.000 1672.310 1409.375 1672.610 ;
        RECT 1396.000 1672.120 1400.000 1672.310 ;
        RECT 1409.045 1672.295 1409.375 1672.310 ;
      LAYER met3 ;
        RECT 300.065 1668.360 1396.000 1671.720 ;
        RECT 300.065 1666.960 1395.600 1668.360 ;
      LAYER met3 ;
        RECT 1396.000 1667.850 1400.000 1667.960 ;
        RECT 1408.125 1667.850 1408.455 1667.865 ;
        RECT 1396.000 1667.550 1408.455 1667.850 ;
        RECT 1396.000 1667.360 1400.000 1667.550 ;
        RECT 1408.125 1667.535 1408.455 1667.550 ;
      LAYER met3 ;
        RECT 300.065 1663.600 1396.000 1666.960 ;
        RECT 304.400 1662.200 1395.600 1663.600 ;
      LAYER met3 ;
        RECT 1396.000 1663.090 1400.000 1663.200 ;
        RECT 1410.885 1663.090 1411.215 1663.105 ;
        RECT 1396.000 1662.790 1411.215 1663.090 ;
        RECT 1396.000 1662.600 1400.000 1662.790 ;
        RECT 1410.885 1662.775 1411.215 1662.790 ;
      LAYER met3 ;
        RECT 300.065 1658.160 1396.000 1662.200 ;
        RECT 300.065 1656.760 1395.600 1658.160 ;
      LAYER met3 ;
        RECT 1396.000 1657.650 1400.000 1657.760 ;
        RECT 1409.505 1657.650 1409.835 1657.665 ;
        RECT 1396.000 1657.350 1409.835 1657.650 ;
        RECT 1396.000 1657.160 1400.000 1657.350 ;
        RECT 1409.505 1657.335 1409.835 1657.350 ;
      LAYER met3 ;
        RECT 300.065 1653.400 1396.000 1656.760 ;
        RECT 304.400 1652.000 1395.600 1653.400 ;
      LAYER met3 ;
        RECT 1396.000 1652.890 1400.000 1653.000 ;
        RECT 1408.125 1652.890 1408.455 1652.905 ;
        RECT 1396.000 1652.590 1408.455 1652.890 ;
        RECT 1396.000 1652.400 1400.000 1652.590 ;
        RECT 1408.125 1652.575 1408.455 1652.590 ;
      LAYER met3 ;
        RECT 300.065 1647.960 1396.000 1652.000 ;
        RECT 300.065 1646.560 1395.600 1647.960 ;
      LAYER met3 ;
        RECT 1396.000 1647.450 1400.000 1647.560 ;
        RECT 1407.665 1647.450 1407.995 1647.465 ;
        RECT 1396.000 1647.150 1407.995 1647.450 ;
        RECT 1396.000 1646.960 1400.000 1647.150 ;
        RECT 1407.665 1647.135 1407.995 1647.150 ;
      LAYER met3 ;
        RECT 300.065 1643.880 1396.000 1646.560 ;
        RECT 304.400 1643.200 1396.000 1643.880 ;
        RECT 304.400 1642.480 1395.600 1643.200 ;
        RECT 300.065 1641.800 1395.600 1642.480 ;
      LAYER met3 ;
        RECT 1396.000 1642.690 1400.000 1642.800 ;
        RECT 1408.125 1642.690 1408.455 1642.705 ;
        RECT 1396.000 1642.390 1408.455 1642.690 ;
        RECT 1396.000 1642.200 1400.000 1642.390 ;
        RECT 1408.125 1642.375 1408.455 1642.390 ;
      LAYER met3 ;
        RECT 300.065 1637.760 1396.000 1641.800 ;
        RECT 300.065 1636.360 1395.600 1637.760 ;
      LAYER met3 ;
        RECT 1396.000 1637.250 1400.000 1637.360 ;
        RECT 1407.665 1637.250 1407.995 1637.265 ;
        RECT 1396.000 1636.950 1407.995 1637.250 ;
        RECT 1396.000 1636.760 1400.000 1636.950 ;
        RECT 1407.665 1636.935 1407.995 1636.950 ;
      LAYER met3 ;
        RECT 300.065 1634.360 1396.000 1636.360 ;
        RECT 304.400 1633.000 1396.000 1634.360 ;
        RECT 304.400 1632.960 1395.600 1633.000 ;
        RECT 300.065 1631.600 1395.600 1632.960 ;
      LAYER met3 ;
        RECT 1396.000 1632.490 1400.000 1632.600 ;
        RECT 1407.665 1632.490 1407.995 1632.505 ;
        RECT 1396.000 1632.190 1407.995 1632.490 ;
        RECT 1396.000 1632.000 1400.000 1632.190 ;
        RECT 1407.665 1632.175 1407.995 1632.190 ;
      LAYER met3 ;
        RECT 300.065 1628.240 1396.000 1631.600 ;
        RECT 300.065 1626.840 1395.600 1628.240 ;
      LAYER met3 ;
        RECT 1396.000 1627.730 1400.000 1627.840 ;
        RECT 1408.585 1627.730 1408.915 1627.745 ;
        RECT 1396.000 1627.430 1408.915 1627.730 ;
        RECT 1396.000 1627.240 1400.000 1627.430 ;
        RECT 1408.585 1627.415 1408.915 1627.430 ;
      LAYER met3 ;
        RECT 300.065 1624.840 1396.000 1626.840 ;
        RECT 304.400 1623.440 1396.000 1624.840 ;
        RECT 300.065 1622.800 1396.000 1623.440 ;
        RECT 300.065 1621.400 1395.600 1622.800 ;
      LAYER met3 ;
        RECT 1396.000 1622.290 1400.000 1622.400 ;
        RECT 1407.665 1622.290 1407.995 1622.305 ;
        RECT 1396.000 1621.990 1407.995 1622.290 ;
        RECT 1396.000 1621.800 1400.000 1621.990 ;
        RECT 1407.665 1621.975 1407.995 1621.990 ;
      LAYER met3 ;
        RECT 300.065 1618.040 1396.000 1621.400 ;
        RECT 300.065 1616.640 1395.600 1618.040 ;
      LAYER met3 ;
        RECT 1396.000 1617.530 1400.000 1617.640 ;
        RECT 1407.665 1617.530 1407.995 1617.545 ;
        RECT 1396.000 1617.230 1407.995 1617.530 ;
        RECT 1396.000 1617.040 1400.000 1617.230 ;
        RECT 1407.665 1617.215 1407.995 1617.230 ;
      LAYER met3 ;
        RECT 300.065 1615.320 1396.000 1616.640 ;
        RECT 304.400 1613.920 1396.000 1615.320 ;
        RECT 300.065 1612.600 1396.000 1613.920 ;
        RECT 300.065 1611.200 1395.600 1612.600 ;
      LAYER met3 ;
        RECT 1396.000 1612.090 1400.000 1612.200 ;
        RECT 1407.665 1612.090 1407.995 1612.105 ;
        RECT 1396.000 1611.790 1407.995 1612.090 ;
        RECT 1396.000 1611.600 1400.000 1611.790 ;
        RECT 1407.665 1611.775 1407.995 1611.790 ;
      LAYER met3 ;
        RECT 300.065 1607.840 1396.000 1611.200 ;
      LAYER met3 ;
        RECT 1688.725 1610.050 1689.055 1610.065 ;
        RECT 1688.725 1609.750 1700.770 1610.050 ;
        RECT 1688.725 1609.735 1689.055 1609.750 ;
        RECT 1700.470 1607.970 1700.770 1609.750 ;
      LAYER met3 ;
        RECT 300.065 1606.440 1395.600 1607.840 ;
      LAYER met3 ;
        RECT 1700.000 1607.670 1704.600 1607.970 ;
        RECT 1396.000 1607.330 1400.000 1607.440 ;
        RECT 1414.105 1607.330 1414.435 1607.345 ;
        RECT 1396.000 1607.030 1414.435 1607.330 ;
        RECT 1396.000 1606.840 1400.000 1607.030 ;
        RECT 1414.105 1607.015 1414.435 1607.030 ;
      LAYER met3 ;
        RECT 300.065 1605.800 1396.000 1606.440 ;
        RECT 304.400 1604.400 1396.000 1605.800 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met3 ;
        RECT 2097.665 1965.010 2097.995 1965.025 ;
        RECT 2085.950 1964.710 2097.995 1965.010 ;
        RECT 2085.950 1963.610 2086.250 1964.710 ;
        RECT 2097.665 1964.695 2097.995 1964.710 ;
        RECT 2081.880 1963.310 2086.480 1963.610 ;
        RECT 2081.880 1954.810 2086.480 1955.110 ;
        RECT 2085.950 1953.450 2086.250 1954.810 ;
        RECT 2097.665 1953.450 2097.995 1953.465 ;
        RECT 2085.950 1953.150 2097.995 1953.450 ;
        RECT 2097.665 1953.135 2097.995 1953.150 ;
        RECT 2081.880 1665.570 2086.480 1665.870 ;
        RECT 2085.950 1663.090 2086.250 1665.570 ;
        RECT 2099.505 1663.090 2099.835 1663.105 ;
        RECT 2085.950 1662.790 2099.835 1663.090 ;
        RECT 2099.505 1662.775 2099.835 1662.790 ;
        RECT 2081.880 1657.070 2086.480 1657.370 ;
        RECT 2085.950 1656.290 2086.250 1657.070 ;
        RECT 2100.885 1656.290 2101.215 1656.305 ;
        RECT 2085.950 1655.990 2101.215 1656.290 ;
        RECT 2100.885 1655.975 2101.215 1655.990 ;
        RECT 2081.880 1651.430 2086.480 1651.730 ;
        RECT 2085.950 1649.490 2086.250 1651.430 ;
        RECT 2099.965 1649.490 2100.295 1649.505 ;
        RECT 2085.950 1649.190 2100.295 1649.490 ;
        RECT 2099.965 1649.175 2100.295 1649.190 ;
        RECT 2099.045 1643.370 2099.375 1643.385 ;
        RECT 2085.950 1643.230 2099.375 1643.370 ;
        RECT 2081.880 1643.070 2099.375 1643.230 ;
        RECT 2081.880 1642.930 2086.480 1643.070 ;
        RECT 2099.045 1643.055 2099.375 1643.070 ;
        RECT 2081.880 1637.290 2086.480 1637.590 ;
        RECT 2085.950 1635.890 2086.250 1637.290 ;
        RECT 2098.585 1635.890 2098.915 1635.905 ;
        RECT 2085.950 1635.590 2098.915 1635.890 ;
        RECT 2098.585 1635.575 2098.915 1635.590 ;
        RECT 2098.125 1629.090 2098.455 1629.105 ;
        RECT 2081.880 1628.790 2098.455 1629.090 ;
        RECT 2098.125 1628.775 2098.455 1628.790 ;
        RECT 2081.880 1623.150 2086.480 1623.450 ;
        RECT 2082.270 1620.265 2082.570 1623.150 ;
        RECT 2082.025 1619.950 2082.570 1620.265 ;
        RECT 2082.025 1619.935 2082.355 1619.950 ;
      LAYER met3 ;
        RECT 300.065 1603.080 1396.000 1604.400 ;
      LAYER met3 ;
        RECT 1725.460 1604.095 1727.200 1605.000 ;
        RECT 1414.105 1603.930 1414.435 1603.945 ;
        RECT 1399.630 1603.630 1414.435 1603.930 ;
      LAYER met3 ;
        RECT 300.065 1602.215 1395.600 1603.080 ;
      LAYER met3 ;
        RECT 1399.630 1602.680 1399.930 1603.630 ;
        RECT 1414.105 1603.615 1414.435 1603.630 ;
        RECT 1396.000 1602.080 1400.000 1602.680 ;
        RECT 1720.005 1593.740 1720.335 1593.745 ;
        RECT 1719.750 1593.730 1720.335 1593.740 ;
        RECT 1719.550 1593.430 1720.335 1593.730 ;
        RECT 1719.750 1593.420 1720.335 1593.430 ;
        RECT 1720.005 1593.415 1720.335 1593.420 ;
        RECT 1738.865 1592.370 1739.195 1592.385 ;
        RECT 1739.990 1592.370 1740.370 1592.380 ;
        RECT 1738.865 1592.070 1740.370 1592.370 ;
        RECT 1738.865 1592.055 1739.195 1592.070 ;
        RECT 1739.990 1592.060 1740.370 1592.070 ;
      LAYER via3 ;
        RECT 646.140 3264.180 646.460 3264.500 ;
        RECT 668.220 3264.180 668.540 3264.500 ;
        RECT 1292.900 3264.180 1293.220 3264.500 ;
        RECT 1890.900 3264.180 1891.220 3264.500 ;
        RECT 1917.580 3264.180 1917.900 3264.500 ;
        RECT 1317.855 3258.060 1318.175 3258.380 ;
        RECT 1055.540 2799.740 1055.860 2800.060 ;
        RECT 1642.400 2799.060 1642.720 2799.380 ;
        RECT 1688.500 2799.060 1688.820 2799.380 ;
        RECT 1794.240 2799.060 1794.560 2799.380 ;
        RECT 1794.300 2798.380 1794.620 2798.700 ;
        RECT 1797.060 2798.380 1797.380 2798.700 ;
        RECT 1759.340 2796.340 1759.660 2796.660 ;
        RECT 1761.180 2795.660 1761.500 2795.980 ;
        RECT 1100.620 2794.980 1100.940 2795.300 ;
        RECT 337.020 2794.300 337.340 2794.620 ;
        RECT 342.540 2794.300 342.860 2794.620 ;
        RECT 350.820 2794.300 351.140 2794.620 ;
        RECT 358.180 2794.300 358.500 2794.620 ;
        RECT 361.860 2794.300 362.180 2794.620 ;
        RECT 364.620 2794.300 364.940 2794.620 ;
        RECT 368.300 2794.300 368.620 2794.620 ;
        RECT 371.060 2794.300 371.380 2794.620 ;
        RECT 374.740 2794.300 375.060 2794.620 ;
        RECT 379.340 2794.300 379.660 2794.620 ;
        RECT 383.940 2794.300 384.260 2794.620 ;
        RECT 386.700 2794.300 387.020 2794.620 ;
        RECT 392.220 2794.300 392.540 2794.620 ;
        RECT 395.900 2794.300 396.220 2794.620 ;
        RECT 399.580 2794.300 399.900 2794.620 ;
        RECT 403.260 2794.300 403.580 2794.620 ;
        RECT 406.020 2794.300 406.340 2794.620 ;
        RECT 409.700 2794.300 410.020 2794.620 ;
        RECT 413.380 2794.300 413.700 2794.620 ;
        RECT 418.900 2794.300 419.220 2794.620 ;
        RECT 420.740 2794.300 421.060 2794.620 ;
        RECT 425.340 2794.300 425.660 2794.620 ;
        RECT 431.780 2794.300 432.100 2794.620 ;
        RECT 433.620 2794.300 433.940 2794.620 ;
        RECT 439.140 2794.300 439.460 2794.620 ;
        RECT 440.980 2794.300 441.300 2794.620 ;
        RECT 444.660 2794.300 444.980 2794.620 ;
        RECT 445.580 2794.300 445.900 2794.620 ;
        RECT 449.260 2794.300 449.580 2794.620 ;
        RECT 454.780 2794.300 455.100 2794.620 ;
        RECT 462.140 2794.300 462.460 2794.620 ;
        RECT 465.820 2794.300 466.140 2794.620 ;
        RECT 474.100 2794.300 474.420 2794.620 ;
        RECT 475.020 2794.300 475.340 2794.620 ;
        RECT 478.700 2794.300 479.020 2794.620 ;
        RECT 482.380 2794.300 482.700 2794.620 ;
        RECT 485.140 2794.300 485.460 2794.620 ;
        RECT 488.820 2794.300 489.140 2794.620 ;
        RECT 490.660 2794.300 490.980 2794.620 ;
        RECT 495.260 2794.300 495.580 2794.620 ;
        RECT 498.020 2794.300 498.340 2794.620 ;
        RECT 500.780 2794.300 501.100 2794.620 ;
        RECT 507.220 2794.300 507.540 2794.620 ;
        RECT 516.420 2794.300 516.740 2794.620 ;
        RECT 523.780 2794.300 524.100 2794.620 ;
        RECT 526.540 2794.300 526.860 2794.620 ;
        RECT 530.220 2794.300 530.540 2794.620 ;
        RECT 535.740 2794.300 536.060 2794.620 ;
        RECT 542.180 2794.300 542.500 2794.620 ;
        RECT 547.700 2794.300 548.020 2794.620 ;
        RECT 981.020 2794.300 981.340 2794.620 ;
        RECT 987.460 2794.300 987.780 2794.620 ;
        RECT 1008.620 2794.300 1008.940 2794.620 ;
        RECT 1013.220 2794.300 1013.540 2794.620 ;
        RECT 1019.660 2794.300 1019.980 2794.620 ;
        RECT 1027.020 2794.300 1027.340 2794.620 ;
        RECT 1030.700 2794.300 1031.020 2794.620 ;
        RECT 1041.740 2794.300 1042.060 2794.620 ;
        RECT 1052.780 2794.300 1053.100 2794.620 ;
        RECT 1059.220 2794.300 1059.540 2794.620 ;
        RECT 1065.660 2794.300 1065.980 2794.620 ;
        RECT 1070.260 2794.300 1070.580 2794.620 ;
        RECT 1076.700 2794.300 1077.020 2794.620 ;
        RECT 1087.740 2794.300 1088.060 2794.620 ;
        RECT 1094.180 2794.300 1094.500 2794.620 ;
        RECT 1111.660 2794.300 1111.980 2794.620 ;
        RECT 1118.100 2794.300 1118.420 2794.620 ;
        RECT 1122.700 2794.300 1123.020 2794.620 ;
        RECT 1129.140 2794.300 1129.460 2794.620 ;
        RECT 1135.580 2794.300 1135.900 2794.620 ;
        RECT 1141.100 2794.300 1141.420 2794.620 ;
        RECT 1147.540 2794.300 1147.860 2794.620 ;
        RECT 1613.980 2794.300 1614.300 2794.620 ;
        RECT 1620.420 2794.300 1620.740 2794.620 ;
        RECT 1625.940 2794.300 1626.260 2794.620 ;
        RECT 1631.460 2794.300 1631.780 2794.620 ;
        RECT 1637.900 2794.300 1638.220 2794.620 ;
        RECT 1648.020 2794.300 1648.340 2794.620 ;
        RECT 1648.940 2794.300 1649.260 2794.620 ;
        RECT 1652.620 2794.300 1652.940 2794.620 ;
        RECT 1661.820 2794.300 1662.140 2794.620 ;
        RECT 1666.420 2794.300 1666.740 2794.620 ;
        RECT 1672.860 2794.300 1673.180 2794.620 ;
        RECT 1679.300 2794.300 1679.620 2794.620 ;
        RECT 1683.900 2794.300 1684.220 2794.620 ;
        RECT 1695.860 2794.300 1696.180 2794.620 ;
        RECT 1702.300 2794.300 1702.620 2794.620 ;
        RECT 1705.980 2794.300 1706.300 2794.620 ;
        RECT 1712.420 2794.300 1712.740 2794.620 ;
        RECT 1717.940 2794.300 1718.260 2794.620 ;
        RECT 1723.460 2794.300 1723.780 2794.620 ;
        RECT 1728.980 2794.300 1729.300 2794.620 ;
        RECT 1734.500 2794.300 1734.820 2794.620 ;
        RECT 1740.940 2794.300 1741.260 2794.620 ;
        RECT 1747.380 2794.300 1747.700 2794.620 ;
        RECT 1794.300 2794.300 1794.620 2794.620 ;
        RECT 1018.740 2793.620 1019.060 2793.940 ;
        RECT 1083.140 2793.620 1083.460 2793.940 ;
        RECT 1164.100 2793.620 1164.420 2793.940 ;
        RECT 1167.780 2793.620 1168.100 2793.940 ;
        RECT 1611.220 2793.620 1611.540 2793.940 ;
        RECT 1617.660 2793.620 1617.980 2793.940 ;
        RECT 1624.100 2793.620 1624.420 2793.940 ;
        RECT 1630.540 2793.620 1630.860 2793.940 ;
        RECT 1635.140 2793.620 1635.460 2793.940 ;
        RECT 1655.380 2793.620 1655.700 2793.940 ;
        RECT 1659.060 2793.620 1659.380 2793.940 ;
        RECT 1663.660 2793.620 1663.980 2793.940 ;
        RECT 1670.100 2793.620 1670.420 2793.940 ;
        RECT 1677.460 2793.620 1677.780 2793.940 ;
        RECT 1682.980 2793.620 1683.300 2793.940 ;
        RECT 1694.940 2793.620 1695.260 2793.940 ;
        RECT 1699.540 2793.620 1699.860 2793.940 ;
        RECT 1767.620 2793.620 1767.940 2793.940 ;
        RECT 1774.060 2793.620 1774.380 2793.940 ;
        RECT 1780.500 2793.620 1780.820 2793.940 ;
        RECT 348.980 2792.940 349.300 2793.260 ;
        RECT 396.820 2792.940 397.140 2793.260 ;
        RECT 414.300 2792.940 414.620 2793.260 ;
        RECT 427.180 2792.940 427.500 2793.260 ;
        RECT 430.860 2792.940 431.180 2793.260 ;
        RECT 455.700 2792.940 456.020 2793.260 ;
        RECT 466.740 2792.940 467.060 2793.260 ;
        RECT 468.580 2792.940 468.900 2793.260 ;
        RECT 501.700 2792.940 502.020 2793.260 ;
        RECT 509.980 2792.940 510.300 2793.260 ;
        RECT 513.660 2792.940 513.980 2793.260 ;
        RECT 520.100 2792.940 520.420 2793.260 ;
        RECT 531.140 2792.940 531.460 2793.260 ;
        RECT 538.500 2792.940 538.820 2793.260 ;
        RECT 543.100 2792.940 543.420 2793.260 ;
        RECT 1012.300 2792.940 1012.620 2793.260 ;
        RECT 1024.260 2792.940 1024.580 2793.260 ;
        RECT 1048.180 2792.940 1048.500 2793.260 ;
        RECT 1175.140 2792.940 1175.460 2793.260 ;
        RECT 1187.100 2792.940 1187.420 2793.260 ;
        RECT 1411.580 2792.940 1411.900 2793.260 ;
        RECT 1180.660 2792.260 1180.980 2792.580 ;
        RECT 1193.540 2792.260 1193.860 2792.580 ;
        RECT 1417.100 2792.260 1417.420 2792.580 ;
        RECT 1752.900 2792.260 1753.220 2792.580 ;
        RECT 1789.700 2792.940 1790.020 2793.260 ;
        RECT 390.380 2791.580 390.700 2791.900 ;
        RECT 460.300 2791.580 460.620 2791.900 ;
        RECT 508.140 2791.580 508.460 2791.900 ;
        RECT 1105.220 2791.580 1105.540 2791.900 ;
        RECT 1153.060 2791.580 1153.380 2791.900 ;
        RECT 1159.500 2791.580 1159.820 2791.900 ;
        RECT 1418.940 2791.580 1419.260 2791.900 ;
        RECT 1787.860 2792.260 1788.180 2792.580 ;
        RECT 378.420 2790.900 378.740 2791.220 ;
        RECT 1418.020 2790.900 1418.340 2791.220 ;
        RECT 1762.100 2790.900 1762.420 2791.220 ;
        RECT 1778.660 2790.900 1778.980 2791.220 ;
        RECT 1587.300 2789.540 1587.620 2789.860 ;
        RECT 1602.940 2789.540 1603.260 2789.860 ;
        RECT 1689.420 2789.540 1689.740 2789.860 ;
        RECT 1001.260 2788.860 1001.580 2789.180 ;
        RECT 993.900 2788.180 994.220 2788.500 ;
        RECT 1035.300 2788.180 1035.620 2788.500 ;
        RECT 1051.860 2788.180 1052.180 2788.500 ;
        RECT 1086.820 2788.180 1087.140 2788.500 ;
        RECT 1128.220 2788.180 1128.540 2788.500 ;
        RECT 1163.180 2788.180 1163.500 2788.500 ;
        RECT 1724.380 2788.180 1724.700 2788.500 ;
        RECT 1765.780 2790.220 1766.100 2790.540 ;
        RECT 1772.220 2789.540 1772.540 2789.860 ;
        RECT 1783.260 2788.180 1783.580 2788.500 ;
        RECT 1034.380 2787.500 1034.700 2787.820 ;
        RECT 1039.900 2787.500 1040.220 2787.820 ;
        RECT 1046.340 2787.500 1046.660 2787.820 ;
        RECT 1061.980 2787.500 1062.300 2787.820 ;
        RECT 1067.500 2787.500 1067.820 2787.820 ;
        RECT 1073.940 2787.500 1074.260 2787.820 ;
        RECT 1081.300 2787.500 1081.620 2787.820 ;
        RECT 1089.580 2787.500 1089.900 2787.820 ;
        RECT 1096.020 2787.500 1096.340 2787.820 ;
        RECT 1103.380 2787.500 1103.700 2787.820 ;
        RECT 1109.820 2787.500 1110.140 2787.820 ;
        RECT 1116.260 2787.500 1116.580 2787.820 ;
        RECT 1121.780 2787.500 1122.100 2787.820 ;
        RECT 1130.980 2787.500 1131.300 2787.820 ;
        RECT 1137.420 2787.500 1137.740 2787.820 ;
        RECT 1143.860 2787.500 1144.180 2787.820 ;
        RECT 1151.220 2787.500 1151.540 2787.820 ;
        RECT 1153.980 2787.500 1154.300 2787.820 ;
        RECT 1165.020 2787.500 1165.340 2787.820 ;
        RECT 1172.380 2787.500 1172.700 2787.820 ;
        RECT 1178.820 2787.500 1179.140 2787.820 ;
        RECT 1186.180 2787.500 1186.500 2787.820 ;
        RECT 1191.700 2787.500 1192.020 2787.820 ;
        RECT 1198.140 2787.500 1198.460 2787.820 ;
        RECT 1581.780 2787.500 1582.100 2787.820 ;
        RECT 1594.660 2787.500 1594.980 2787.820 ;
        RECT 1604.780 2787.500 1605.100 2787.820 ;
        RECT 1708.740 2787.500 1709.060 2787.820 ;
        RECT 1713.340 2787.500 1713.660 2787.820 ;
        RECT 1719.780 2787.500 1720.100 2787.820 ;
        RECT 1730.820 2787.500 1731.140 2787.820 ;
        RECT 1737.260 2787.500 1737.580 2787.820 ;
        RECT 1743.700 2787.500 1744.020 2787.820 ;
        RECT 1748.300 2787.500 1748.620 2787.820 ;
        RECT 1754.740 2787.500 1755.060 2787.820 ;
        RECT 1644.340 2785.460 1644.660 2785.780 ;
        RECT 1838.460 2069.420 1838.780 2069.740 ;
        RECT 1844.900 2069.420 1845.220 2069.740 ;
        RECT 1851.340 2069.420 1851.660 2069.740 ;
        RECT 1857.780 2069.420 1858.100 2069.740 ;
        RECT 1863.300 2069.420 1863.620 2069.740 ;
        RECT 1869.740 2069.420 1870.060 2069.740 ;
        RECT 1879.860 2069.420 1880.180 2069.740 ;
        RECT 1886.300 2069.420 1886.620 2069.740 ;
        RECT 1891.820 2069.420 1892.140 2069.740 ;
        RECT 1898.260 2069.420 1898.580 2069.740 ;
        RECT 1904.700 2069.420 1905.020 2069.740 ;
        RECT 1911.140 2069.420 1911.460 2069.740 ;
        RECT 1925.860 2069.420 1926.180 2069.740 ;
        RECT 1873.420 2068.740 1873.740 2069.060 ;
        RECT 1914.820 2068.740 1915.140 2069.060 ;
        RECT 1920.340 2068.740 1920.660 2069.060 ;
        RECT 1981.980 2068.060 1982.300 2068.380 ;
        RECT 1987.500 2068.060 1987.820 2068.380 ;
        RECT 2028.900 2067.380 2029.220 2067.700 ;
        RECT 1841.220 2066.700 1841.540 2067.020 ;
        RECT 1848.580 2066.700 1848.900 2067.020 ;
        RECT 1889.980 2066.700 1890.300 2067.020 ;
        RECT 1941.500 2066.700 1941.820 2067.020 ;
        RECT 2023.380 2066.700 2023.700 2067.020 ;
        RECT 1855.020 2066.020 1855.340 2066.340 ;
        RECT 1901.020 2066.020 1901.340 2066.340 ;
        RECT 1934.140 2066.020 1934.460 2066.340 ;
        RECT 2011.420 2066.020 2011.740 2066.340 ;
        RECT 2016.940 2066.020 2017.260 2066.340 ;
        RECT 2037.180 2066.020 2037.500 2066.340 ;
        RECT 1859.620 2065.340 1859.940 2065.660 ;
        RECT 1865.140 2065.340 1865.460 2065.660 ;
        RECT 1894.580 2065.340 1894.900 2065.660 ;
        RECT 1907.460 2065.340 1907.780 2065.660 ;
        RECT 1912.060 2065.340 1912.380 2065.660 ;
        RECT 1935.980 2065.340 1936.300 2065.660 ;
        RECT 1999.460 2065.340 1999.780 2065.660 ;
        RECT 2043.620 2065.340 2043.940 2065.660 ;
        RECT 1871.580 2064.660 1871.900 2064.980 ;
        RECT 1917.580 2064.660 1917.900 2064.980 ;
        RECT 1924.020 2064.660 1924.340 2064.980 ;
        RECT 1929.540 2064.660 1929.860 2064.980 ;
        RECT 2005.900 2064.660 2006.220 2064.980 ;
        RECT 1877.100 2063.980 1877.420 2064.300 ;
        RECT 1882.620 2063.980 1882.940 2064.300 ;
        RECT 1967.260 2063.980 1967.580 2064.300 ;
        RECT 1993.020 2063.980 1993.340 2064.300 ;
        RECT 1947.940 2063.300 1948.260 2063.620 ;
        RECT 1954.380 2063.300 1954.700 2063.620 ;
        RECT 1958.980 2063.300 1959.300 2063.620 ;
        RECT 1965.420 2063.300 1965.740 2063.620 ;
        RECT 1970.020 2063.300 1970.340 2063.620 ;
        RECT 1973.700 2063.300 1974.020 2063.620 ;
        RECT 1976.460 2063.300 1976.780 2063.620 ;
        RECT 1980.140 2063.300 1980.460 2063.620 ;
        RECT 2031.660 2063.300 2031.980 2063.620 ;
        RECT 1940.580 2058.540 1940.900 2058.860 ;
        RECT 1955.300 2057.860 1955.620 2058.180 ;
        RECT 1987.300 2057.860 1987.620 2058.180 ;
        RECT 1995.780 2057.860 1996.100 2058.180 ;
        RECT 1946.420 2057.180 1946.740 2057.500 ;
        RECT 1990.260 2057.180 1990.580 2057.500 ;
        RECT 2004.820 2057.180 2005.140 2057.500 ;
        RECT 2016.500 2057.180 2016.820 2057.500 ;
        RECT 2008.660 2056.500 2008.980 2056.820 ;
        RECT 2021.540 2056.500 2021.860 2056.820 ;
        RECT 1948.860 2055.140 1949.180 2055.460 ;
        RECT 1961.510 2051.740 1961.830 2052.060 ;
        RECT 2050.060 2051.740 2050.380 2052.060 ;
        RECT 1418.020 1985.780 1418.340 1986.100 ;
        RECT 1418.940 1980.340 1419.260 1980.660 ;
        RECT 1417.100 1975.580 1417.420 1975.900 ;
        RECT 1411.580 1955.180 1411.900 1955.500 ;
        RECT 1719.780 1593.420 1720.100 1593.740 ;
        RECT 1740.020 1592.060 1740.340 1592.380 ;
      LAYER met4 ;
        RECT 646.135 3264.175 646.465 3264.505 ;
        RECT 668.215 3264.175 668.545 3264.505 ;
        RECT 1292.895 3264.175 1293.225 3264.505 ;
        RECT 1890.895 3264.175 1891.225 3264.505 ;
        RECT 1917.575 3264.175 1917.905 3264.505 ;
        RECT 394.025 3251.635 394.325 3256.235 ;
        RECT 400.265 3251.635 400.565 3256.235 ;
        RECT 406.505 3251.635 406.805 3256.235 ;
        RECT 412.745 3251.635 413.045 3256.235 ;
        RECT 418.985 3251.635 419.285 3256.235 ;
        RECT 425.225 3251.635 425.525 3256.235 ;
        RECT 431.465 3251.635 431.765 3256.235 ;
        RECT 437.705 3251.635 438.005 3256.235 ;
        RECT 443.945 3251.635 444.245 3256.235 ;
        RECT 450.185 3251.635 450.485 3256.235 ;
        RECT 456.425 3251.635 456.725 3256.235 ;
        RECT 462.665 3251.635 462.965 3256.235 ;
        RECT 468.905 3251.635 469.205 3256.235 ;
        RECT 475.145 3251.635 475.445 3256.235 ;
        RECT 481.385 3251.635 481.685 3256.235 ;
        RECT 487.625 3251.635 487.925 3256.235 ;
        RECT 493.865 3251.635 494.165 3256.235 ;
        RECT 500.105 3251.635 500.405 3256.235 ;
        RECT 506.345 3251.635 506.645 3256.235 ;
        RECT 512.585 3251.635 512.885 3256.235 ;
        RECT 518.825 3251.635 519.125 3256.235 ;
        RECT 525.065 3251.635 525.365 3256.235 ;
        RECT 531.305 3251.635 531.605 3256.235 ;
        RECT 537.545 3251.635 537.845 3256.235 ;
        RECT 543.785 3251.635 544.085 3256.235 ;
        RECT 550.025 3251.635 550.325 3256.235 ;
        RECT 556.265 3251.635 556.565 3256.235 ;
        RECT 562.505 3251.635 562.805 3256.235 ;
        RECT 568.745 3251.635 569.045 3256.235 ;
        RECT 574.985 3251.635 575.285 3256.235 ;
        RECT 581.225 3251.635 581.525 3256.235 ;
        RECT 587.465 3251.635 587.765 3256.235 ;
        RECT 642.890 3255.650 643.190 3256.235 ;
        RECT 646.150 3255.650 646.450 3264.175 ;
        RECT 668.230 3259.050 668.530 3264.175 ;
        RECT 642.890 3255.350 646.450 3255.650 ;
        RECT 667.865 3258.750 668.530 3259.050 ;
        RECT 642.890 3251.635 643.190 3255.350 ;
        RECT 667.865 3251.635 668.165 3258.750 ;
        RECT 1292.910 3256.235 1293.210 3264.175 ;
        RECT 1317.850 3258.055 1318.180 3258.385 ;
        RECT 1044.025 3251.635 1044.325 3256.235 ;
        RECT 1050.265 3251.635 1050.565 3256.235 ;
        RECT 1056.505 3251.635 1056.805 3256.235 ;
        RECT 1062.745 3251.635 1063.045 3256.235 ;
        RECT 1068.985 3251.635 1069.285 3256.235 ;
        RECT 1075.225 3251.635 1075.525 3256.235 ;
        RECT 1081.465 3251.635 1081.765 3256.235 ;
        RECT 1087.705 3251.635 1088.005 3256.235 ;
        RECT 1093.945 3251.635 1094.245 3256.235 ;
        RECT 1100.185 3251.635 1100.485 3256.235 ;
        RECT 1106.425 3251.635 1106.725 3256.235 ;
        RECT 1112.665 3251.635 1112.965 3256.235 ;
        RECT 1118.905 3251.635 1119.205 3256.235 ;
        RECT 1125.145 3251.635 1125.445 3256.235 ;
        RECT 1131.385 3251.635 1131.685 3256.235 ;
        RECT 1137.625 3251.635 1137.925 3256.235 ;
        RECT 1143.865 3251.635 1144.165 3256.235 ;
        RECT 1150.105 3251.635 1150.405 3256.235 ;
        RECT 1156.345 3251.635 1156.645 3256.235 ;
        RECT 1162.585 3251.635 1162.885 3256.235 ;
        RECT 1168.825 3251.635 1169.125 3256.235 ;
        RECT 1175.065 3251.635 1175.365 3256.235 ;
        RECT 1181.305 3251.635 1181.605 3256.235 ;
        RECT 1187.545 3251.635 1187.845 3256.235 ;
        RECT 1193.785 3251.635 1194.085 3256.235 ;
        RECT 1200.025 3251.635 1200.325 3256.235 ;
        RECT 1206.265 3251.635 1206.565 3256.235 ;
        RECT 1212.505 3251.635 1212.805 3256.235 ;
        RECT 1218.745 3251.635 1219.045 3256.235 ;
        RECT 1224.985 3251.635 1225.285 3256.235 ;
        RECT 1231.225 3251.635 1231.525 3256.235 ;
        RECT 1237.465 3251.635 1237.765 3256.235 ;
        RECT 1292.890 3255.350 1293.210 3256.235 ;
        RECT 1292.890 3251.635 1293.190 3255.350 ;
        RECT 1317.865 3251.635 1318.165 3258.055 ;
        RECT 1644.025 3251.635 1644.325 3256.235 ;
        RECT 1650.265 3251.635 1650.565 3256.235 ;
        RECT 1656.505 3251.635 1656.805 3256.235 ;
        RECT 1662.745 3251.635 1663.045 3256.235 ;
        RECT 1668.985 3251.635 1669.285 3256.235 ;
        RECT 1675.225 3251.635 1675.525 3256.235 ;
        RECT 1681.465 3251.635 1681.765 3256.235 ;
        RECT 1687.705 3251.635 1688.005 3256.235 ;
        RECT 1693.945 3251.635 1694.245 3256.235 ;
        RECT 1700.185 3251.635 1700.485 3256.235 ;
        RECT 1706.425 3251.635 1706.725 3256.235 ;
        RECT 1712.665 3251.635 1712.965 3256.235 ;
        RECT 1718.905 3251.635 1719.205 3256.235 ;
        RECT 1725.145 3251.635 1725.445 3256.235 ;
        RECT 1731.385 3251.635 1731.685 3256.235 ;
        RECT 1737.625 3251.635 1737.925 3256.235 ;
        RECT 1743.865 3251.635 1744.165 3256.235 ;
        RECT 1750.105 3251.635 1750.405 3256.235 ;
        RECT 1756.345 3251.635 1756.645 3256.235 ;
        RECT 1762.585 3251.635 1762.885 3256.235 ;
        RECT 1768.825 3251.635 1769.125 3256.235 ;
        RECT 1775.065 3251.635 1775.365 3256.235 ;
        RECT 1781.305 3251.635 1781.605 3256.235 ;
        RECT 1787.545 3251.635 1787.845 3256.235 ;
        RECT 1793.785 3251.635 1794.085 3256.235 ;
        RECT 1800.025 3251.635 1800.325 3256.235 ;
        RECT 1806.265 3251.635 1806.565 3256.235 ;
        RECT 1812.505 3251.635 1812.805 3256.235 ;
        RECT 1818.745 3251.635 1819.045 3256.235 ;
        RECT 1824.985 3251.635 1825.285 3256.235 ;
        RECT 1831.225 3251.635 1831.525 3256.235 ;
        RECT 1837.465 3251.635 1837.765 3256.235 ;
        RECT 1890.910 3255.650 1891.210 3264.175 ;
        RECT 1917.590 3256.235 1917.890 3264.175 ;
        RECT 1892.890 3255.650 1893.190 3256.235 ;
        RECT 1890.910 3255.350 1893.190 3255.650 ;
        RECT 1917.590 3255.350 1918.165 3256.235 ;
        RECT 1892.890 3251.635 1893.190 3255.350 ;
        RECT 1917.865 3251.635 1918.165 3255.350 ;
      LAYER met4 ;
        RECT 305.000 2805.000 681.480 3251.235 ;
        RECT 955.000 2805.000 1331.480 3251.235 ;
        RECT 1555.000 2805.000 1931.480 3251.235 ;
      LAYER met4 ;
        RECT 334.010 2801.750 334.310 2804.600 ;
        RECT 339.850 2801.750 340.150 2804.600 ;
        RECT 345.690 2801.750 345.990 2804.600 ;
        RECT 351.530 2801.750 351.830 2804.600 ;
        RECT 334.010 2801.450 337.330 2801.750 ;
        RECT 334.010 2800.000 334.310 2801.450 ;
        RECT 337.030 2794.625 337.330 2801.450 ;
        RECT 339.850 2801.450 342.850 2801.750 ;
        RECT 339.850 2800.000 340.150 2801.450 ;
        RECT 342.550 2794.625 342.850 2801.450 ;
        RECT 345.690 2801.450 349.290 2801.750 ;
        RECT 345.690 2800.000 345.990 2801.450 ;
        RECT 337.015 2794.295 337.345 2794.625 ;
        RECT 342.535 2794.295 342.865 2794.625 ;
        RECT 348.990 2793.265 349.290 2801.450 ;
        RECT 350.830 2801.450 351.830 2801.750 ;
        RECT 350.830 2794.625 351.130 2801.450 ;
        RECT 351.530 2800.000 351.830 2801.450 ;
        RECT 357.370 2801.750 357.670 2804.600 ;
        RECT 363.210 2802.450 363.510 2804.600 ;
        RECT 361.870 2802.150 363.510 2802.450 ;
        RECT 357.370 2801.450 358.490 2801.750 ;
        RECT 357.370 2800.000 357.670 2801.450 ;
        RECT 358.190 2794.625 358.490 2801.450 ;
        RECT 361.870 2794.625 362.170 2802.150 ;
        RECT 363.210 2800.000 363.510 2802.150 ;
        RECT 363.830 2801.750 364.130 2804.600 ;
        RECT 369.050 2801.750 369.350 2804.600 ;
        RECT 363.830 2801.450 364.930 2801.750 ;
        RECT 363.830 2800.000 364.130 2801.450 ;
        RECT 364.630 2794.625 364.930 2801.450 ;
        RECT 368.310 2801.450 369.350 2801.750 ;
        RECT 368.310 2794.625 368.610 2801.450 ;
        RECT 369.050 2800.000 369.350 2801.450 ;
        RECT 369.670 2801.750 369.970 2804.600 ;
        RECT 374.890 2801.750 375.190 2804.600 ;
        RECT 369.670 2801.450 371.370 2801.750 ;
        RECT 369.670 2800.000 369.970 2801.450 ;
        RECT 371.070 2794.625 371.370 2801.450 ;
        RECT 374.750 2800.000 375.190 2801.750 ;
        RECT 375.510 2801.750 375.810 2804.600 ;
        RECT 380.730 2801.750 381.030 2804.600 ;
        RECT 375.510 2801.450 378.730 2801.750 ;
        RECT 375.510 2800.000 375.810 2801.450 ;
        RECT 374.750 2794.625 375.050 2800.000 ;
        RECT 350.815 2794.295 351.145 2794.625 ;
        RECT 358.175 2794.295 358.505 2794.625 ;
        RECT 361.855 2794.295 362.185 2794.625 ;
        RECT 364.615 2794.295 364.945 2794.625 ;
        RECT 368.295 2794.295 368.625 2794.625 ;
        RECT 371.055 2794.295 371.385 2794.625 ;
        RECT 374.735 2794.295 375.065 2794.625 ;
        RECT 348.975 2792.935 349.305 2793.265 ;
        RECT 378.430 2791.225 378.730 2801.450 ;
        RECT 379.350 2801.450 381.030 2801.750 ;
        RECT 379.350 2794.625 379.650 2801.450 ;
        RECT 380.730 2800.000 381.030 2801.450 ;
        RECT 381.350 2801.750 381.650 2804.600 ;
        RECT 381.350 2801.450 384.250 2801.750 ;
        RECT 381.350 2800.000 381.650 2801.450 ;
        RECT 383.950 2794.625 384.250 2801.450 ;
        RECT 386.570 2796.650 386.870 2804.600 ;
        RECT 387.190 2801.750 387.490 2804.600 ;
        RECT 392.410 2801.750 392.710 2804.600 ;
        RECT 387.190 2801.450 390.690 2801.750 ;
        RECT 387.190 2800.000 387.490 2801.450 ;
        RECT 386.570 2796.350 387.010 2796.650 ;
        RECT 386.710 2794.625 387.010 2796.350 ;
        RECT 379.335 2794.295 379.665 2794.625 ;
        RECT 383.935 2794.295 384.265 2794.625 ;
        RECT 386.695 2794.295 387.025 2794.625 ;
        RECT 390.390 2791.905 390.690 2801.450 ;
        RECT 392.230 2800.000 392.710 2801.750 ;
        RECT 393.030 2801.750 393.330 2804.600 ;
        RECT 398.250 2802.450 398.550 2804.600 ;
        RECT 396.830 2802.150 398.550 2802.450 ;
        RECT 393.030 2801.450 396.210 2801.750 ;
        RECT 393.030 2800.000 393.330 2801.450 ;
        RECT 392.230 2794.625 392.530 2800.000 ;
        RECT 395.910 2794.625 396.210 2801.450 ;
        RECT 392.215 2794.295 392.545 2794.625 ;
        RECT 395.895 2794.295 396.225 2794.625 ;
        RECT 396.830 2793.265 397.130 2802.150 ;
        RECT 398.250 2800.000 398.550 2802.150 ;
        RECT 398.870 2801.750 399.170 2804.600 ;
        RECT 404.090 2801.750 404.390 2804.600 ;
        RECT 398.870 2801.450 399.890 2801.750 ;
        RECT 398.870 2800.000 399.170 2801.450 ;
        RECT 399.590 2794.625 399.890 2801.450 ;
        RECT 403.270 2801.450 404.390 2801.750 ;
        RECT 403.270 2794.625 403.570 2801.450 ;
        RECT 404.090 2800.000 404.390 2801.450 ;
        RECT 404.710 2801.750 405.010 2804.600 ;
        RECT 409.930 2801.750 410.230 2804.600 ;
        RECT 404.710 2801.450 406.330 2801.750 ;
        RECT 404.710 2800.000 405.010 2801.450 ;
        RECT 406.030 2794.625 406.330 2801.450 ;
        RECT 409.710 2800.000 410.230 2801.750 ;
        RECT 410.550 2801.750 410.850 2804.600 ;
        RECT 415.770 2801.750 416.070 2804.600 ;
        RECT 410.550 2801.450 413.690 2801.750 ;
        RECT 410.550 2800.000 410.850 2801.450 ;
        RECT 409.710 2794.625 410.010 2800.000 ;
        RECT 413.390 2794.625 413.690 2801.450 ;
        RECT 414.310 2801.450 416.070 2801.750 ;
        RECT 399.575 2794.295 399.905 2794.625 ;
        RECT 403.255 2794.295 403.585 2794.625 ;
        RECT 406.015 2794.295 406.345 2794.625 ;
        RECT 409.695 2794.295 410.025 2794.625 ;
        RECT 413.375 2794.295 413.705 2794.625 ;
        RECT 414.310 2793.265 414.610 2801.450 ;
        RECT 415.770 2800.000 416.070 2801.450 ;
        RECT 416.390 2801.750 416.690 2804.600 ;
        RECT 421.610 2801.750 421.910 2804.600 ;
        RECT 416.390 2801.450 419.210 2801.750 ;
        RECT 416.390 2800.000 416.690 2801.450 ;
        RECT 418.910 2794.625 419.210 2801.450 ;
        RECT 420.750 2801.450 421.910 2801.750 ;
        RECT 420.750 2794.625 421.050 2801.450 ;
        RECT 421.610 2800.000 421.910 2801.450 ;
        RECT 422.230 2801.750 422.530 2804.600 ;
        RECT 427.450 2801.750 427.750 2804.600 ;
        RECT 422.230 2801.450 425.650 2801.750 ;
        RECT 422.230 2800.000 422.530 2801.450 ;
        RECT 425.350 2794.625 425.650 2801.450 ;
        RECT 427.190 2800.000 427.750 2801.750 ;
        RECT 428.070 2801.750 428.370 2804.600 ;
        RECT 433.290 2802.450 433.590 2804.600 ;
        RECT 431.790 2802.150 433.590 2802.450 ;
        RECT 428.070 2801.450 431.170 2801.750 ;
        RECT 428.070 2800.000 428.370 2801.450 ;
        RECT 418.895 2794.295 419.225 2794.625 ;
        RECT 420.735 2794.295 421.065 2794.625 ;
        RECT 425.335 2794.295 425.665 2794.625 ;
        RECT 427.190 2793.265 427.490 2800.000 ;
        RECT 430.870 2793.265 431.170 2801.450 ;
        RECT 431.790 2794.625 432.090 2802.150 ;
        RECT 433.290 2800.000 433.590 2802.150 ;
        RECT 433.910 2796.650 434.210 2804.600 ;
        RECT 439.130 2800.050 439.430 2804.600 ;
        RECT 439.750 2801.750 440.050 2804.600 ;
        RECT 444.970 2801.750 445.270 2804.600 ;
        RECT 439.750 2801.450 441.290 2801.750 ;
        RECT 439.130 2799.750 439.450 2800.050 ;
        RECT 439.750 2800.000 440.050 2801.450 ;
        RECT 433.630 2796.350 434.210 2796.650 ;
        RECT 433.630 2794.625 433.930 2796.350 ;
        RECT 439.150 2794.625 439.450 2799.750 ;
        RECT 440.990 2794.625 441.290 2801.450 ;
        RECT 444.670 2800.000 445.270 2801.750 ;
        RECT 444.670 2794.625 444.970 2800.000 ;
        RECT 445.590 2794.625 445.890 2804.600 ;
        RECT 450.810 2801.750 451.110 2804.600 ;
        RECT 449.270 2801.450 451.110 2801.750 ;
        RECT 449.270 2794.625 449.570 2801.450 ;
        RECT 450.810 2800.000 451.110 2801.450 ;
        RECT 451.430 2801.750 451.730 2804.600 ;
        RECT 456.650 2801.750 456.950 2804.600 ;
        RECT 451.430 2801.450 455.090 2801.750 ;
        RECT 451.430 2800.000 451.730 2801.450 ;
        RECT 454.790 2794.625 455.090 2801.450 ;
        RECT 455.710 2801.450 456.950 2801.750 ;
        RECT 431.775 2794.295 432.105 2794.625 ;
        RECT 433.615 2794.295 433.945 2794.625 ;
        RECT 439.135 2794.295 439.465 2794.625 ;
        RECT 440.975 2794.295 441.305 2794.625 ;
        RECT 444.655 2794.295 444.985 2794.625 ;
        RECT 445.575 2794.295 445.905 2794.625 ;
        RECT 449.255 2794.295 449.585 2794.625 ;
        RECT 454.775 2794.295 455.105 2794.625 ;
        RECT 455.710 2793.265 456.010 2801.450 ;
        RECT 456.650 2800.000 456.950 2801.450 ;
        RECT 457.270 2801.750 457.570 2804.600 ;
        RECT 457.270 2801.450 460.610 2801.750 ;
        RECT 457.270 2800.000 457.570 2801.450 ;
        RECT 396.815 2792.935 397.145 2793.265 ;
        RECT 414.295 2792.935 414.625 2793.265 ;
        RECT 427.175 2792.935 427.505 2793.265 ;
        RECT 430.855 2792.935 431.185 2793.265 ;
        RECT 455.695 2792.935 456.025 2793.265 ;
        RECT 460.310 2791.905 460.610 2801.450 ;
        RECT 462.490 2800.050 462.790 2804.600 ;
        RECT 462.150 2799.750 462.790 2800.050 ;
        RECT 463.110 2801.750 463.410 2804.600 ;
        RECT 468.330 2801.750 468.630 2804.600 ;
        RECT 463.110 2801.450 466.130 2801.750 ;
        RECT 463.110 2800.000 463.410 2801.450 ;
        RECT 462.150 2794.625 462.450 2799.750 ;
        RECT 465.830 2794.625 466.130 2801.450 ;
        RECT 466.750 2801.450 468.630 2801.750 ;
        RECT 462.135 2794.295 462.465 2794.625 ;
        RECT 465.815 2794.295 466.145 2794.625 ;
        RECT 466.750 2793.265 467.050 2801.450 ;
        RECT 468.330 2800.000 468.630 2801.450 ;
        RECT 468.950 2796.650 469.250 2804.600 ;
        RECT 474.170 2801.750 474.470 2804.600 ;
        RECT 468.590 2796.350 469.250 2796.650 ;
        RECT 474.110 2800.000 474.470 2801.750 ;
        RECT 474.790 2801.750 475.090 2804.600 ;
        RECT 480.010 2802.450 480.310 2804.600 ;
        RECT 478.710 2802.150 480.310 2802.450 ;
        RECT 474.790 2800.000 475.330 2801.750 ;
        RECT 468.590 2793.265 468.890 2796.350 ;
        RECT 474.110 2794.625 474.410 2800.000 ;
        RECT 475.030 2794.625 475.330 2800.000 ;
        RECT 478.710 2794.625 479.010 2802.150 ;
        RECT 480.010 2800.000 480.310 2802.150 ;
        RECT 480.630 2801.750 480.930 2804.600 ;
        RECT 485.850 2801.750 486.150 2804.600 ;
        RECT 480.630 2801.450 482.690 2801.750 ;
        RECT 480.630 2800.000 480.930 2801.450 ;
        RECT 482.390 2794.625 482.690 2801.450 ;
        RECT 485.150 2801.450 486.150 2801.750 ;
        RECT 485.150 2794.625 485.450 2801.450 ;
        RECT 485.850 2800.000 486.150 2801.450 ;
        RECT 486.470 2801.750 486.770 2804.600 ;
        RECT 491.690 2801.750 491.990 2804.600 ;
        RECT 486.470 2801.450 489.130 2801.750 ;
        RECT 486.470 2800.000 486.770 2801.450 ;
        RECT 488.830 2794.625 489.130 2801.450 ;
        RECT 490.670 2801.450 491.990 2801.750 ;
        RECT 490.670 2794.625 490.970 2801.450 ;
        RECT 491.690 2800.000 491.990 2801.450 ;
        RECT 492.310 2801.750 492.610 2804.600 ;
        RECT 492.310 2801.450 495.570 2801.750 ;
        RECT 492.310 2800.000 492.610 2801.450 ;
        RECT 495.270 2794.625 495.570 2801.450 ;
        RECT 497.530 2796.650 497.830 2804.600 ;
        RECT 498.150 2801.750 498.450 2804.600 ;
        RECT 503.370 2801.750 503.670 2804.600 ;
        RECT 498.150 2801.450 501.090 2801.750 ;
        RECT 498.150 2800.000 498.450 2801.450 ;
        RECT 497.530 2796.350 498.330 2796.650 ;
        RECT 498.030 2794.625 498.330 2796.350 ;
        RECT 500.790 2794.625 501.090 2801.450 ;
        RECT 501.710 2801.450 503.670 2801.750 ;
        RECT 474.095 2794.295 474.425 2794.625 ;
        RECT 475.015 2794.295 475.345 2794.625 ;
        RECT 478.695 2794.295 479.025 2794.625 ;
        RECT 482.375 2794.295 482.705 2794.625 ;
        RECT 485.135 2794.295 485.465 2794.625 ;
        RECT 488.815 2794.295 489.145 2794.625 ;
        RECT 490.655 2794.295 490.985 2794.625 ;
        RECT 495.255 2794.295 495.585 2794.625 ;
        RECT 498.015 2794.295 498.345 2794.625 ;
        RECT 500.775 2794.295 501.105 2794.625 ;
        RECT 501.710 2793.265 502.010 2801.450 ;
        RECT 503.370 2800.000 503.670 2801.450 ;
        RECT 503.990 2801.750 504.290 2804.600 ;
        RECT 509.210 2801.750 509.510 2804.600 ;
        RECT 503.990 2801.450 507.530 2801.750 ;
        RECT 503.990 2800.000 504.290 2801.450 ;
        RECT 507.230 2794.625 507.530 2801.450 ;
        RECT 508.150 2801.450 509.510 2801.750 ;
        RECT 507.215 2794.295 507.545 2794.625 ;
        RECT 466.735 2792.935 467.065 2793.265 ;
        RECT 468.575 2792.935 468.905 2793.265 ;
        RECT 501.695 2792.935 502.025 2793.265 ;
        RECT 508.150 2791.905 508.450 2801.450 ;
        RECT 509.210 2800.000 509.510 2801.450 ;
        RECT 509.830 2801.750 510.130 2804.600 ;
        RECT 515.050 2802.450 515.350 2804.600 ;
        RECT 513.670 2802.150 515.350 2802.450 ;
        RECT 509.830 2800.000 510.290 2801.750 ;
        RECT 509.990 2793.265 510.290 2800.000 ;
        RECT 513.670 2793.265 513.970 2802.150 ;
        RECT 515.050 2800.000 515.350 2802.150 ;
        RECT 515.670 2801.750 515.970 2804.600 ;
        RECT 520.890 2801.750 521.190 2804.600 ;
        RECT 515.670 2801.450 516.730 2801.750 ;
        RECT 515.670 2800.000 515.970 2801.450 ;
        RECT 516.430 2794.625 516.730 2801.450 ;
        RECT 520.110 2801.450 521.190 2801.750 ;
        RECT 516.415 2794.295 516.745 2794.625 ;
        RECT 520.110 2793.265 520.410 2801.450 ;
        RECT 520.890 2800.000 521.190 2801.450 ;
        RECT 521.510 2801.750 521.810 2804.600 ;
        RECT 526.730 2801.750 527.030 2804.600 ;
        RECT 521.510 2801.450 524.090 2801.750 ;
        RECT 521.510 2800.000 521.810 2801.450 ;
        RECT 523.790 2794.625 524.090 2801.450 ;
        RECT 526.550 2800.000 527.030 2801.750 ;
        RECT 527.350 2801.750 527.650 2804.600 ;
        RECT 532.570 2802.450 532.870 2804.600 ;
        RECT 531.150 2802.150 532.870 2802.450 ;
        RECT 527.350 2801.450 530.530 2801.750 ;
        RECT 527.350 2800.000 527.650 2801.450 ;
        RECT 526.550 2794.625 526.850 2800.000 ;
        RECT 530.230 2794.625 530.530 2801.450 ;
        RECT 523.775 2794.295 524.105 2794.625 ;
        RECT 526.535 2794.295 526.865 2794.625 ;
        RECT 530.215 2794.295 530.545 2794.625 ;
        RECT 531.150 2793.265 531.450 2802.150 ;
        RECT 532.570 2800.000 532.870 2802.150 ;
        RECT 533.190 2801.750 533.490 2804.600 ;
        RECT 533.190 2801.450 536.050 2801.750 ;
        RECT 533.190 2800.000 533.490 2801.450 ;
        RECT 535.750 2794.625 536.050 2801.450 ;
        RECT 538.410 2796.650 538.710 2804.600 ;
        RECT 539.030 2801.750 539.330 2804.600 ;
        RECT 544.250 2801.750 544.550 2804.600 ;
        RECT 539.030 2801.450 542.490 2801.750 ;
        RECT 539.030 2800.000 539.330 2801.450 ;
        RECT 538.410 2796.350 538.810 2796.650 ;
        RECT 535.735 2794.295 536.065 2794.625 ;
        RECT 538.510 2793.265 538.810 2796.350 ;
        RECT 542.190 2794.625 542.490 2801.450 ;
        RECT 543.110 2801.450 544.550 2801.750 ;
        RECT 542.175 2794.295 542.505 2794.625 ;
        RECT 543.110 2793.265 543.410 2801.450 ;
        RECT 544.250 2800.000 544.550 2801.450 ;
        RECT 544.870 2801.750 545.170 2804.600 ;
        RECT 984.010 2801.750 984.310 2804.600 ;
        RECT 989.850 2801.750 990.150 2804.600 ;
        RECT 995.690 2801.750 995.990 2804.600 ;
        RECT 1001.530 2801.750 1001.830 2804.600 ;
        RECT 544.870 2801.450 548.010 2801.750 ;
        RECT 544.870 2800.000 545.170 2801.450 ;
        RECT 547.710 2794.625 548.010 2801.450 ;
        RECT 981.030 2801.450 984.310 2801.750 ;
        RECT 981.030 2794.625 981.330 2801.450 ;
        RECT 984.010 2800.000 984.310 2801.450 ;
        RECT 987.470 2801.450 990.150 2801.750 ;
        RECT 987.470 2794.625 987.770 2801.450 ;
        RECT 989.850 2800.000 990.150 2801.450 ;
        RECT 993.910 2801.450 995.990 2801.750 ;
        RECT 547.695 2794.295 548.025 2794.625 ;
        RECT 981.015 2794.295 981.345 2794.625 ;
        RECT 987.455 2794.295 987.785 2794.625 ;
        RECT 509.975 2792.935 510.305 2793.265 ;
        RECT 513.655 2792.935 513.985 2793.265 ;
        RECT 520.095 2792.935 520.425 2793.265 ;
        RECT 531.135 2792.935 531.465 2793.265 ;
        RECT 538.495 2792.935 538.825 2793.265 ;
        RECT 543.095 2792.935 543.425 2793.265 ;
        RECT 390.375 2791.575 390.705 2791.905 ;
        RECT 460.295 2791.575 460.625 2791.905 ;
        RECT 508.135 2791.575 508.465 2791.905 ;
        RECT 378.415 2790.895 378.745 2791.225 ;
        RECT 993.910 2788.505 994.210 2801.450 ;
        RECT 995.690 2800.000 995.990 2801.450 ;
        RECT 1001.270 2800.000 1001.830 2801.750 ;
        RECT 1007.370 2802.450 1007.670 2804.600 ;
        RECT 1007.370 2802.150 1008.930 2802.450 ;
        RECT 1007.370 2800.000 1007.670 2802.150 ;
        RECT 1001.270 2789.185 1001.570 2800.000 ;
        RECT 1008.630 2794.625 1008.930 2802.150 ;
        RECT 1013.210 2801.750 1013.510 2804.600 ;
        RECT 1012.310 2801.450 1013.510 2801.750 ;
        RECT 1008.615 2794.295 1008.945 2794.625 ;
        RECT 1012.310 2793.265 1012.610 2801.450 ;
        RECT 1013.210 2800.000 1013.510 2801.450 ;
        RECT 1013.830 2796.650 1014.130 2804.600 ;
        RECT 1019.050 2801.750 1019.350 2804.600 ;
        RECT 1013.230 2796.350 1014.130 2796.650 ;
        RECT 1018.750 2800.000 1019.350 2801.750 ;
        RECT 1013.230 2794.625 1013.530 2796.350 ;
        RECT 1013.215 2794.295 1013.545 2794.625 ;
        RECT 1018.750 2793.945 1019.050 2800.000 ;
        RECT 1019.670 2794.625 1019.970 2804.600 ;
        RECT 1024.890 2801.750 1025.190 2804.600 ;
        RECT 1024.270 2801.450 1025.190 2801.750 ;
        RECT 1019.655 2794.295 1019.985 2794.625 ;
        RECT 1018.735 2793.615 1019.065 2793.945 ;
        RECT 1024.270 2793.265 1024.570 2801.450 ;
        RECT 1024.890 2800.000 1025.190 2801.450 ;
        RECT 1025.510 2801.750 1025.810 2804.600 ;
        RECT 1030.730 2801.750 1031.030 2804.600 ;
        RECT 1025.510 2801.450 1027.330 2801.750 ;
        RECT 1025.510 2800.000 1025.810 2801.450 ;
        RECT 1027.030 2794.625 1027.330 2801.450 ;
        RECT 1030.710 2800.000 1031.030 2801.750 ;
        RECT 1031.350 2801.750 1031.650 2804.600 ;
        RECT 1036.570 2802.450 1036.870 2804.600 ;
        RECT 1035.310 2802.150 1036.870 2802.450 ;
        RECT 1031.350 2801.450 1034.690 2801.750 ;
        RECT 1031.350 2800.000 1031.650 2801.450 ;
        RECT 1030.710 2794.625 1031.010 2800.000 ;
        RECT 1027.015 2794.295 1027.345 2794.625 ;
        RECT 1030.695 2794.295 1031.025 2794.625 ;
        RECT 1012.295 2792.935 1012.625 2793.265 ;
        RECT 1024.255 2792.935 1024.585 2793.265 ;
        RECT 1001.255 2788.855 1001.585 2789.185 ;
        RECT 993.895 2788.175 994.225 2788.505 ;
        RECT 1034.390 2787.825 1034.690 2801.450 ;
        RECT 1035.310 2788.505 1035.610 2802.150 ;
        RECT 1036.570 2800.000 1036.870 2802.150 ;
        RECT 1037.190 2801.750 1037.490 2804.600 ;
        RECT 1042.410 2801.750 1042.710 2804.600 ;
        RECT 1037.190 2801.450 1040.210 2801.750 ;
        RECT 1037.190 2800.000 1037.490 2801.450 ;
        RECT 1035.295 2788.175 1035.625 2788.505 ;
        RECT 1039.910 2787.825 1040.210 2801.450 ;
        RECT 1041.750 2801.450 1042.710 2801.750 ;
        RECT 1041.750 2794.625 1042.050 2801.450 ;
        RECT 1042.410 2800.000 1042.710 2801.450 ;
        RECT 1043.030 2801.750 1043.330 2804.600 ;
        RECT 1048.250 2801.750 1048.550 2804.600 ;
        RECT 1043.030 2801.450 1046.650 2801.750 ;
        RECT 1043.030 2800.000 1043.330 2801.450 ;
        RECT 1041.735 2794.295 1042.065 2794.625 ;
        RECT 1046.350 2787.825 1046.650 2801.450 ;
        RECT 1048.190 2800.000 1048.550 2801.750 ;
        RECT 1048.870 2801.750 1049.170 2804.600 ;
        RECT 1054.090 2801.750 1054.390 2804.600 ;
        RECT 1048.870 2801.450 1052.170 2801.750 ;
        RECT 1048.870 2800.000 1049.170 2801.450 ;
        RECT 1048.190 2793.265 1048.490 2800.000 ;
        RECT 1048.175 2792.935 1048.505 2793.265 ;
        RECT 1051.870 2788.505 1052.170 2801.450 ;
        RECT 1052.790 2801.450 1054.390 2801.750 ;
        RECT 1052.790 2794.625 1053.090 2801.450 ;
        RECT 1054.090 2800.000 1054.390 2801.450 ;
        RECT 1054.710 2800.050 1055.010 2804.600 ;
        RECT 1059.930 2801.750 1060.230 2804.600 ;
        RECT 1059.230 2801.450 1060.230 2801.750 ;
        RECT 1055.535 2800.050 1055.865 2800.065 ;
        RECT 1054.710 2799.750 1055.865 2800.050 ;
        RECT 1055.535 2799.735 1055.865 2799.750 ;
        RECT 1059.230 2794.625 1059.530 2801.450 ;
        RECT 1059.930 2800.000 1060.230 2801.450 ;
        RECT 1060.550 2801.750 1060.850 2804.600 ;
        RECT 1065.770 2801.750 1066.070 2804.600 ;
        RECT 1060.550 2801.450 1062.290 2801.750 ;
        RECT 1060.550 2800.000 1060.850 2801.450 ;
        RECT 1052.775 2794.295 1053.105 2794.625 ;
        RECT 1059.215 2794.295 1059.545 2794.625 ;
        RECT 1051.855 2788.175 1052.185 2788.505 ;
        RECT 1061.990 2787.825 1062.290 2801.450 ;
        RECT 1065.670 2800.000 1066.070 2801.750 ;
        RECT 1066.390 2801.750 1066.690 2804.600 ;
        RECT 1071.610 2801.750 1071.910 2804.600 ;
        RECT 1066.390 2801.450 1067.810 2801.750 ;
        RECT 1066.390 2800.000 1066.690 2801.450 ;
        RECT 1065.670 2794.625 1065.970 2800.000 ;
        RECT 1065.655 2794.295 1065.985 2794.625 ;
        RECT 1067.510 2787.825 1067.810 2801.450 ;
        RECT 1070.270 2801.450 1071.910 2801.750 ;
        RECT 1070.270 2794.625 1070.570 2801.450 ;
        RECT 1071.610 2800.000 1071.910 2801.450 ;
        RECT 1072.230 2801.750 1072.530 2804.600 ;
        RECT 1077.450 2801.750 1077.750 2804.600 ;
        RECT 1072.230 2801.450 1074.250 2801.750 ;
        RECT 1072.230 2800.000 1072.530 2801.450 ;
        RECT 1070.255 2794.295 1070.585 2794.625 ;
        RECT 1073.950 2787.825 1074.250 2801.450 ;
        RECT 1076.710 2801.450 1077.750 2801.750 ;
        RECT 1076.710 2794.625 1077.010 2801.450 ;
        RECT 1077.450 2800.000 1077.750 2801.450 ;
        RECT 1078.070 2801.750 1078.370 2804.600 ;
        RECT 1083.290 2801.750 1083.590 2804.600 ;
        RECT 1078.070 2801.450 1081.610 2801.750 ;
        RECT 1078.070 2800.000 1078.370 2801.450 ;
        RECT 1076.695 2794.295 1077.025 2794.625 ;
        RECT 1081.310 2787.825 1081.610 2801.450 ;
        RECT 1083.150 2800.000 1083.590 2801.750 ;
        RECT 1083.910 2801.750 1084.210 2804.600 ;
        RECT 1089.130 2802.450 1089.430 2804.600 ;
        RECT 1087.750 2802.150 1089.430 2802.450 ;
        RECT 1083.910 2801.450 1087.130 2801.750 ;
        RECT 1083.910 2800.000 1084.210 2801.450 ;
        RECT 1083.150 2793.945 1083.450 2800.000 ;
        RECT 1083.135 2793.615 1083.465 2793.945 ;
        RECT 1086.830 2788.505 1087.130 2801.450 ;
        RECT 1087.750 2794.625 1088.050 2802.150 ;
        RECT 1089.130 2800.000 1089.430 2802.150 ;
        RECT 1089.750 2796.650 1090.050 2804.600 ;
        RECT 1094.970 2801.750 1095.270 2804.600 ;
        RECT 1089.590 2796.350 1090.050 2796.650 ;
        RECT 1094.190 2801.450 1095.270 2801.750 ;
        RECT 1087.735 2794.295 1088.065 2794.625 ;
        RECT 1086.815 2788.175 1087.145 2788.505 ;
        RECT 1089.590 2787.825 1089.890 2796.350 ;
        RECT 1094.190 2794.625 1094.490 2801.450 ;
        RECT 1094.970 2800.000 1095.270 2801.450 ;
        RECT 1095.590 2800.050 1095.890 2804.600 ;
        RECT 1100.810 2801.750 1101.110 2804.600 ;
        RECT 1095.590 2799.750 1096.330 2800.050 ;
        RECT 1094.175 2794.295 1094.505 2794.625 ;
        RECT 1096.030 2787.825 1096.330 2799.750 ;
        RECT 1100.630 2800.000 1101.110 2801.750 ;
        RECT 1101.430 2801.750 1101.730 2804.600 ;
        RECT 1106.650 2802.450 1106.950 2804.600 ;
        RECT 1105.230 2802.150 1106.950 2802.450 ;
        RECT 1101.430 2801.450 1103.690 2801.750 ;
        RECT 1101.430 2800.000 1101.730 2801.450 ;
        RECT 1100.630 2795.305 1100.930 2800.000 ;
        RECT 1100.615 2794.975 1100.945 2795.305 ;
        RECT 1103.390 2787.825 1103.690 2801.450 ;
        RECT 1105.230 2791.905 1105.530 2802.150 ;
        RECT 1106.650 2800.000 1106.950 2802.150 ;
        RECT 1107.270 2801.750 1107.570 2804.600 ;
        RECT 1112.490 2801.750 1112.790 2804.600 ;
        RECT 1107.270 2801.450 1110.130 2801.750 ;
        RECT 1107.270 2800.000 1107.570 2801.450 ;
        RECT 1105.215 2791.575 1105.545 2791.905 ;
        RECT 1109.830 2787.825 1110.130 2801.450 ;
        RECT 1111.670 2801.450 1112.790 2801.750 ;
        RECT 1111.670 2794.625 1111.970 2801.450 ;
        RECT 1112.490 2800.000 1112.790 2801.450 ;
        RECT 1113.110 2801.750 1113.410 2804.600 ;
        RECT 1118.330 2801.750 1118.630 2804.600 ;
        RECT 1113.110 2801.450 1116.570 2801.750 ;
        RECT 1113.110 2800.000 1113.410 2801.450 ;
        RECT 1111.655 2794.295 1111.985 2794.625 ;
        RECT 1116.270 2787.825 1116.570 2801.450 ;
        RECT 1118.110 2800.000 1118.630 2801.750 ;
        RECT 1118.950 2801.750 1119.250 2804.600 ;
        RECT 1124.170 2801.750 1124.470 2804.600 ;
        RECT 1118.950 2801.450 1122.090 2801.750 ;
        RECT 1118.950 2800.000 1119.250 2801.450 ;
        RECT 1118.110 2794.625 1118.410 2800.000 ;
        RECT 1118.095 2794.295 1118.425 2794.625 ;
        RECT 1121.790 2787.825 1122.090 2801.450 ;
        RECT 1122.710 2801.450 1124.470 2801.750 ;
        RECT 1122.710 2794.625 1123.010 2801.450 ;
        RECT 1124.170 2800.000 1124.470 2801.450 ;
        RECT 1124.790 2801.750 1125.090 2804.600 ;
        RECT 1130.010 2801.750 1130.310 2804.600 ;
        RECT 1124.790 2801.450 1128.530 2801.750 ;
        RECT 1124.790 2800.000 1125.090 2801.450 ;
        RECT 1122.695 2794.295 1123.025 2794.625 ;
        RECT 1128.230 2788.505 1128.530 2801.450 ;
        RECT 1129.150 2801.450 1130.310 2801.750 ;
        RECT 1129.150 2794.625 1129.450 2801.450 ;
        RECT 1130.010 2800.000 1130.310 2801.450 ;
        RECT 1130.630 2800.050 1130.930 2804.600 ;
        RECT 1135.850 2801.750 1136.150 2804.600 ;
        RECT 1130.630 2799.750 1131.290 2800.050 ;
        RECT 1129.135 2794.295 1129.465 2794.625 ;
        RECT 1128.215 2788.175 1128.545 2788.505 ;
        RECT 1130.990 2787.825 1131.290 2799.750 ;
        RECT 1135.590 2800.000 1136.150 2801.750 ;
        RECT 1136.470 2801.750 1136.770 2804.600 ;
        RECT 1136.470 2801.450 1137.730 2801.750 ;
        RECT 1136.470 2800.000 1136.770 2801.450 ;
        RECT 1135.590 2794.625 1135.890 2800.000 ;
        RECT 1135.575 2794.295 1135.905 2794.625 ;
        RECT 1137.430 2787.825 1137.730 2801.450 ;
        RECT 1141.690 2796.650 1141.990 2804.600 ;
        RECT 1142.310 2801.750 1142.610 2804.600 ;
        RECT 1142.310 2801.450 1144.170 2801.750 ;
        RECT 1142.310 2800.000 1142.610 2801.450 ;
        RECT 1141.110 2796.350 1141.990 2796.650 ;
        RECT 1141.110 2794.625 1141.410 2796.350 ;
        RECT 1141.095 2794.295 1141.425 2794.625 ;
        RECT 1143.870 2787.825 1144.170 2801.450 ;
        RECT 1147.530 2800.050 1147.830 2804.600 ;
        RECT 1148.150 2801.750 1148.450 2804.600 ;
        RECT 1153.370 2801.750 1153.670 2804.600 ;
        RECT 1148.150 2801.450 1151.530 2801.750 ;
        RECT 1147.530 2799.750 1147.850 2800.050 ;
        RECT 1148.150 2800.000 1148.450 2801.450 ;
        RECT 1147.550 2794.625 1147.850 2799.750 ;
        RECT 1147.535 2794.295 1147.865 2794.625 ;
        RECT 1151.230 2787.825 1151.530 2801.450 ;
        RECT 1153.070 2800.000 1153.670 2801.750 ;
        RECT 1153.070 2791.905 1153.370 2800.000 ;
        RECT 1153.055 2791.575 1153.385 2791.905 ;
        RECT 1153.990 2787.825 1154.290 2804.600 ;
        RECT 1159.210 2796.650 1159.510 2804.600 ;
        RECT 1159.830 2801.750 1160.130 2804.600 ;
        RECT 1165.050 2801.750 1165.350 2804.600 ;
        RECT 1159.830 2801.450 1163.490 2801.750 ;
        RECT 1159.830 2800.000 1160.130 2801.450 ;
        RECT 1159.210 2796.350 1159.810 2796.650 ;
        RECT 1159.510 2791.905 1159.810 2796.350 ;
        RECT 1159.495 2791.575 1159.825 2791.905 ;
        RECT 1163.190 2788.505 1163.490 2801.450 ;
        RECT 1164.110 2801.450 1165.350 2801.750 ;
        RECT 1164.110 2793.945 1164.410 2801.450 ;
        RECT 1165.050 2800.000 1165.350 2801.450 ;
        RECT 1165.670 2796.650 1165.970 2804.600 ;
        RECT 1170.890 2801.750 1171.190 2804.600 ;
        RECT 1165.030 2796.350 1165.970 2796.650 ;
        RECT 1167.790 2801.450 1171.190 2801.750 ;
        RECT 1164.095 2793.615 1164.425 2793.945 ;
        RECT 1163.175 2788.175 1163.505 2788.505 ;
        RECT 1165.030 2787.825 1165.330 2796.350 ;
        RECT 1167.790 2793.945 1168.090 2801.450 ;
        RECT 1170.890 2800.000 1171.190 2801.450 ;
        RECT 1171.510 2801.750 1171.810 2804.600 ;
        RECT 1176.730 2801.750 1177.030 2804.600 ;
        RECT 1171.510 2801.450 1172.690 2801.750 ;
        RECT 1171.510 2800.000 1171.810 2801.450 ;
        RECT 1167.775 2793.615 1168.105 2793.945 ;
        RECT 1172.390 2787.825 1172.690 2801.450 ;
        RECT 1175.150 2801.450 1177.030 2801.750 ;
        RECT 1175.150 2793.265 1175.450 2801.450 ;
        RECT 1176.730 2800.000 1177.030 2801.450 ;
        RECT 1177.350 2801.750 1177.650 2804.600 ;
        RECT 1182.570 2801.750 1182.870 2804.600 ;
        RECT 1177.350 2801.450 1179.130 2801.750 ;
        RECT 1177.350 2800.000 1177.650 2801.450 ;
        RECT 1175.135 2792.935 1175.465 2793.265 ;
        RECT 1178.830 2787.825 1179.130 2801.450 ;
        RECT 1180.670 2801.450 1182.870 2801.750 ;
        RECT 1180.670 2792.585 1180.970 2801.450 ;
        RECT 1182.570 2800.000 1182.870 2801.450 ;
        RECT 1183.190 2801.750 1183.490 2804.600 ;
        RECT 1188.410 2801.750 1188.710 2804.600 ;
        RECT 1183.190 2801.450 1186.490 2801.750 ;
        RECT 1183.190 2800.000 1183.490 2801.450 ;
        RECT 1180.655 2792.255 1180.985 2792.585 ;
        RECT 1186.190 2787.825 1186.490 2801.450 ;
        RECT 1187.110 2801.450 1188.710 2801.750 ;
        RECT 1187.110 2793.265 1187.410 2801.450 ;
        RECT 1188.410 2800.000 1188.710 2801.450 ;
        RECT 1189.030 2801.750 1189.330 2804.600 ;
        RECT 1194.250 2801.750 1194.550 2804.600 ;
        RECT 1189.030 2801.450 1192.010 2801.750 ;
        RECT 1189.030 2800.000 1189.330 2801.450 ;
        RECT 1187.095 2792.935 1187.425 2793.265 ;
        RECT 1191.710 2787.825 1192.010 2801.450 ;
        RECT 1193.550 2801.450 1194.550 2801.750 ;
        RECT 1193.550 2792.585 1193.850 2801.450 ;
        RECT 1194.250 2800.000 1194.550 2801.450 ;
        RECT 1194.870 2801.750 1195.170 2804.600 ;
        RECT 1584.010 2801.750 1584.310 2804.600 ;
        RECT 1589.850 2801.750 1590.150 2804.600 ;
        RECT 1595.690 2801.750 1595.990 2804.600 ;
        RECT 1194.870 2801.450 1198.450 2801.750 ;
        RECT 1194.870 2800.000 1195.170 2801.450 ;
        RECT 1193.535 2792.255 1193.865 2792.585 ;
        RECT 1198.150 2787.825 1198.450 2801.450 ;
        RECT 1581.790 2801.450 1584.310 2801.750 ;
        RECT 1411.575 2792.935 1411.905 2793.265 ;
        RECT 1034.375 2787.495 1034.705 2787.825 ;
        RECT 1039.895 2787.495 1040.225 2787.825 ;
        RECT 1046.335 2787.495 1046.665 2787.825 ;
        RECT 1061.975 2787.495 1062.305 2787.825 ;
        RECT 1067.495 2787.495 1067.825 2787.825 ;
        RECT 1073.935 2787.495 1074.265 2787.825 ;
        RECT 1081.295 2787.495 1081.625 2787.825 ;
        RECT 1089.575 2787.495 1089.905 2787.825 ;
        RECT 1096.015 2787.495 1096.345 2787.825 ;
        RECT 1103.375 2787.495 1103.705 2787.825 ;
        RECT 1109.815 2787.495 1110.145 2787.825 ;
        RECT 1116.255 2787.495 1116.585 2787.825 ;
        RECT 1121.775 2787.495 1122.105 2787.825 ;
        RECT 1130.975 2787.495 1131.305 2787.825 ;
        RECT 1137.415 2787.495 1137.745 2787.825 ;
        RECT 1143.855 2787.495 1144.185 2787.825 ;
        RECT 1151.215 2787.495 1151.545 2787.825 ;
        RECT 1153.975 2787.495 1154.305 2787.825 ;
        RECT 1165.015 2787.495 1165.345 2787.825 ;
        RECT 1172.375 2787.495 1172.705 2787.825 ;
        RECT 1178.815 2787.495 1179.145 2787.825 ;
        RECT 1186.175 2787.495 1186.505 2787.825 ;
        RECT 1191.695 2787.495 1192.025 2787.825 ;
        RECT 1198.135 2787.495 1198.465 2787.825 ;
        RECT 292.020 2715.000 295.020 2785.000 ;
        RECT 310.020 2715.000 313.020 2785.000 ;
        RECT 328.020 2715.000 331.020 2785.000 ;
        RECT 364.020 2715.000 367.020 2785.000 ;
        RECT 454.020 2715.000 457.020 2785.000 ;
        RECT 472.020 2715.000 475.020 2785.000 ;
        RECT 490.020 2715.000 493.020 2785.000 ;
        RECT 508.020 2715.000 511.020 2785.000 ;
        RECT 544.020 2715.000 547.020 2785.000 ;
        RECT 634.020 2715.000 637.020 2785.000 ;
        RECT 652.020 2715.000 655.020 2785.000 ;
        RECT 670.020 2715.000 673.020 2785.000 ;
        RECT 688.020 2715.000 691.020 2785.000 ;
        RECT 994.020 2715.000 997.020 2785.000 ;
        RECT 1012.020 2715.000 1015.020 2785.000 ;
        RECT 1030.020 2715.000 1033.020 2785.000 ;
        RECT 1048.020 2715.000 1051.020 2785.000 ;
        RECT 1084.020 2715.000 1087.020 2785.000 ;
        RECT 1174.020 2715.000 1177.020 2785.000 ;
        RECT 1192.020 2715.000 1195.020 2785.000 ;
        RECT 1210.020 2715.000 1213.020 2785.000 ;
        RECT 1228.020 2715.000 1231.020 2785.000 ;
        RECT 1264.020 2715.000 1267.020 2785.000 ;
      LAYER met4 ;
        RECT 323.295 2688.640 1389.905 2697.345 ;
        RECT 323.295 1610.240 397.440 2688.640 ;
        RECT 399.840 1610.240 1389.905 2688.640 ;
      LAYER met4 ;
        RECT 1411.590 1955.505 1411.890 2792.935 ;
        RECT 1417.095 2792.255 1417.425 2792.585 ;
        RECT 1417.110 1975.905 1417.410 2792.255 ;
        RECT 1418.935 2791.575 1419.265 2791.905 ;
        RECT 1418.015 2790.895 1418.345 2791.225 ;
        RECT 1418.030 1986.105 1418.330 2790.895 ;
        RECT 1418.015 1985.775 1418.345 1986.105 ;
        RECT 1418.950 1980.665 1419.250 2791.575 ;
        RECT 1581.790 2787.825 1582.090 2801.450 ;
        RECT 1584.010 2800.000 1584.310 2801.450 ;
        RECT 1587.310 2801.450 1590.150 2801.750 ;
        RECT 1587.310 2789.865 1587.610 2801.450 ;
        RECT 1589.850 2800.000 1590.150 2801.450 ;
        RECT 1594.670 2801.450 1595.990 2801.750 ;
        RECT 1587.295 2789.535 1587.625 2789.865 ;
        RECT 1594.670 2787.825 1594.970 2801.450 ;
        RECT 1595.690 2800.000 1595.990 2801.450 ;
        RECT 1601.530 2802.450 1601.830 2804.600 ;
        RECT 1601.530 2802.150 1603.250 2802.450 ;
        RECT 1601.530 2800.000 1601.830 2802.150 ;
        RECT 1602.950 2789.865 1603.250 2802.150 ;
        RECT 1607.370 2801.750 1607.670 2804.600 ;
        RECT 1613.210 2801.750 1613.510 2804.600 ;
        RECT 1604.790 2801.450 1607.670 2801.750 ;
        RECT 1602.935 2789.535 1603.265 2789.865 ;
        RECT 1604.790 2787.825 1605.090 2801.450 ;
        RECT 1607.370 2800.000 1607.670 2801.450 ;
        RECT 1611.230 2801.450 1613.510 2801.750 ;
        RECT 1611.230 2793.945 1611.530 2801.450 ;
        RECT 1613.210 2800.000 1613.510 2801.450 ;
        RECT 1613.830 2801.750 1614.130 2804.600 ;
        RECT 1619.050 2802.450 1619.350 2804.600 ;
        RECT 1617.670 2802.150 1619.350 2802.450 ;
        RECT 1613.830 2800.000 1614.290 2801.750 ;
        RECT 1613.990 2794.625 1614.290 2800.000 ;
        RECT 1613.975 2794.295 1614.305 2794.625 ;
        RECT 1617.670 2793.945 1617.970 2802.150 ;
        RECT 1619.050 2800.000 1619.350 2802.150 ;
        RECT 1619.670 2801.750 1619.970 2804.600 ;
        RECT 1624.890 2801.750 1625.190 2804.600 ;
        RECT 1619.670 2801.450 1620.730 2801.750 ;
        RECT 1619.670 2800.000 1619.970 2801.450 ;
        RECT 1620.430 2794.625 1620.730 2801.450 ;
        RECT 1624.110 2801.450 1625.190 2801.750 ;
        RECT 1620.415 2794.295 1620.745 2794.625 ;
        RECT 1624.110 2793.945 1624.410 2801.450 ;
        RECT 1624.890 2800.000 1625.190 2801.450 ;
        RECT 1625.510 2800.050 1625.810 2804.600 ;
        RECT 1630.730 2801.750 1631.030 2804.600 ;
        RECT 1625.510 2799.750 1626.250 2800.050 ;
        RECT 1625.950 2794.625 1626.250 2799.750 ;
        RECT 1630.550 2800.000 1631.030 2801.750 ;
        RECT 1631.350 2801.750 1631.650 2804.600 ;
        RECT 1636.570 2802.450 1636.870 2804.600 ;
        RECT 1635.150 2802.150 1636.870 2802.450 ;
        RECT 1631.350 2800.000 1631.770 2801.750 ;
        RECT 1625.935 2794.295 1626.265 2794.625 ;
        RECT 1630.550 2793.945 1630.850 2800.000 ;
        RECT 1631.470 2794.625 1631.770 2800.000 ;
        RECT 1631.455 2794.295 1631.785 2794.625 ;
        RECT 1635.150 2793.945 1635.450 2802.150 ;
        RECT 1636.570 2800.000 1636.870 2802.150 ;
        RECT 1637.190 2801.750 1637.490 2804.600 ;
        RECT 1637.190 2801.450 1638.210 2801.750 ;
        RECT 1637.190 2800.000 1637.490 2801.450 ;
        RECT 1637.910 2794.625 1638.210 2801.450 ;
        RECT 1642.410 2799.385 1642.710 2804.600 ;
        RECT 1643.030 2802.450 1643.330 2804.600 ;
        RECT 1643.030 2802.150 1644.650 2802.450 ;
        RECT 1643.030 2800.000 1643.330 2802.150 ;
        RECT 1642.395 2799.055 1642.725 2799.385 ;
        RECT 1637.895 2794.295 1638.225 2794.625 ;
        RECT 1611.215 2793.615 1611.545 2793.945 ;
        RECT 1617.655 2793.615 1617.985 2793.945 ;
        RECT 1624.095 2793.615 1624.425 2793.945 ;
        RECT 1630.535 2793.615 1630.865 2793.945 ;
        RECT 1635.135 2793.615 1635.465 2793.945 ;
        RECT 1581.775 2787.495 1582.105 2787.825 ;
        RECT 1594.655 2787.495 1594.985 2787.825 ;
        RECT 1604.775 2787.495 1605.105 2787.825 ;
        RECT 1644.350 2785.785 1644.650 2802.150 ;
        RECT 1648.250 2801.750 1648.550 2804.600 ;
        RECT 1648.030 2800.000 1648.550 2801.750 ;
        RECT 1648.870 2801.750 1649.170 2804.600 ;
        RECT 1654.090 2802.450 1654.390 2804.600 ;
        RECT 1652.630 2802.150 1654.390 2802.450 ;
        RECT 1648.870 2800.000 1649.250 2801.750 ;
        RECT 1648.030 2794.625 1648.330 2800.000 ;
        RECT 1648.950 2794.625 1649.250 2800.000 ;
        RECT 1652.630 2794.625 1652.930 2802.150 ;
        RECT 1654.090 2800.000 1654.390 2802.150 ;
        RECT 1654.710 2801.750 1655.010 2804.600 ;
        RECT 1659.930 2801.750 1660.230 2804.600 ;
        RECT 1654.710 2801.450 1655.690 2801.750 ;
        RECT 1654.710 2800.000 1655.010 2801.450 ;
        RECT 1648.015 2794.295 1648.345 2794.625 ;
        RECT 1648.935 2794.295 1649.265 2794.625 ;
        RECT 1652.615 2794.295 1652.945 2794.625 ;
        RECT 1655.390 2793.945 1655.690 2801.450 ;
        RECT 1659.070 2801.450 1660.230 2801.750 ;
        RECT 1659.070 2793.945 1659.370 2801.450 ;
        RECT 1659.930 2800.000 1660.230 2801.450 ;
        RECT 1660.550 2802.450 1660.850 2804.600 ;
        RECT 1660.550 2802.150 1662.130 2802.450 ;
        RECT 1660.550 2800.000 1660.850 2802.150 ;
        RECT 1661.830 2794.625 1662.130 2802.150 ;
        RECT 1665.770 2801.750 1666.070 2804.600 ;
        RECT 1663.670 2801.450 1666.070 2801.750 ;
        RECT 1661.815 2794.295 1662.145 2794.625 ;
        RECT 1663.670 2793.945 1663.970 2801.450 ;
        RECT 1665.770 2800.000 1666.070 2801.450 ;
        RECT 1666.390 2801.750 1666.690 2804.600 ;
        RECT 1671.610 2802.450 1671.910 2804.600 ;
        RECT 1670.110 2802.150 1671.910 2802.450 ;
        RECT 1666.390 2800.000 1666.730 2801.750 ;
        RECT 1666.430 2794.625 1666.730 2800.000 ;
        RECT 1666.415 2794.295 1666.745 2794.625 ;
        RECT 1670.110 2793.945 1670.410 2802.150 ;
        RECT 1671.610 2800.000 1671.910 2802.150 ;
        RECT 1672.230 2801.750 1672.530 2804.600 ;
        RECT 1672.230 2801.450 1673.170 2801.750 ;
        RECT 1672.230 2800.000 1672.530 2801.450 ;
        RECT 1672.870 2794.625 1673.170 2801.450 ;
        RECT 1677.450 2800.050 1677.750 2804.600 ;
        RECT 1678.070 2802.450 1678.370 2804.600 ;
        RECT 1678.070 2802.150 1679.610 2802.450 ;
        RECT 1677.450 2799.750 1677.770 2800.050 ;
        RECT 1678.070 2800.000 1678.370 2802.150 ;
        RECT 1672.855 2794.295 1673.185 2794.625 ;
        RECT 1677.470 2793.945 1677.770 2799.750 ;
        RECT 1679.310 2794.625 1679.610 2802.150 ;
        RECT 1683.290 2801.750 1683.590 2804.600 ;
        RECT 1682.990 2800.000 1683.590 2801.750 ;
        RECT 1679.295 2794.295 1679.625 2794.625 ;
        RECT 1682.990 2793.945 1683.290 2800.000 ;
        RECT 1683.910 2794.625 1684.210 2804.600 ;
        RECT 1689.130 2801.750 1689.430 2804.600 ;
        RECT 1688.510 2801.450 1689.430 2801.750 ;
        RECT 1688.510 2799.385 1688.810 2801.450 ;
        RECT 1689.130 2800.000 1689.430 2801.450 ;
        RECT 1688.495 2799.055 1688.825 2799.385 ;
        RECT 1689.750 2796.650 1690.050 2804.600 ;
        RECT 1694.970 2801.750 1695.270 2804.600 ;
        RECT 1689.430 2796.350 1690.050 2796.650 ;
        RECT 1694.950 2800.000 1695.270 2801.750 ;
        RECT 1695.590 2801.750 1695.890 2804.600 ;
        RECT 1700.810 2802.450 1701.110 2804.600 ;
        RECT 1699.550 2802.150 1701.110 2802.450 ;
        RECT 1695.590 2800.000 1696.170 2801.750 ;
        RECT 1683.895 2794.295 1684.225 2794.625 ;
        RECT 1655.375 2793.615 1655.705 2793.945 ;
        RECT 1659.055 2793.615 1659.385 2793.945 ;
        RECT 1663.655 2793.615 1663.985 2793.945 ;
        RECT 1670.095 2793.615 1670.425 2793.945 ;
        RECT 1677.455 2793.615 1677.785 2793.945 ;
        RECT 1682.975 2793.615 1683.305 2793.945 ;
        RECT 1689.430 2789.865 1689.730 2796.350 ;
        RECT 1694.950 2793.945 1695.250 2800.000 ;
        RECT 1695.870 2794.625 1696.170 2800.000 ;
        RECT 1695.855 2794.295 1696.185 2794.625 ;
        RECT 1699.550 2793.945 1699.850 2802.150 ;
        RECT 1700.810 2800.000 1701.110 2802.150 ;
        RECT 1701.430 2801.750 1701.730 2804.600 ;
        RECT 1706.650 2801.750 1706.950 2804.600 ;
        RECT 1701.430 2801.450 1702.610 2801.750 ;
        RECT 1701.430 2800.000 1701.730 2801.450 ;
        RECT 1702.310 2794.625 1702.610 2801.450 ;
        RECT 1705.990 2801.450 1706.950 2801.750 ;
        RECT 1705.990 2794.625 1706.290 2801.450 ;
        RECT 1706.650 2800.000 1706.950 2801.450 ;
        RECT 1707.270 2802.450 1707.570 2804.600 ;
        RECT 1707.270 2802.150 1709.050 2802.450 ;
        RECT 1707.270 2800.000 1707.570 2802.150 ;
        RECT 1702.295 2794.295 1702.625 2794.625 ;
        RECT 1705.975 2794.295 1706.305 2794.625 ;
        RECT 1694.935 2793.615 1695.265 2793.945 ;
        RECT 1699.535 2793.615 1699.865 2793.945 ;
        RECT 1689.415 2789.535 1689.745 2789.865 ;
        RECT 1708.750 2787.825 1709.050 2802.150 ;
        RECT 1712.490 2801.750 1712.790 2804.600 ;
        RECT 1712.430 2800.000 1712.790 2801.750 ;
        RECT 1713.110 2801.750 1713.410 2804.600 ;
        RECT 1713.110 2800.000 1713.650 2801.750 ;
        RECT 1718.330 2800.050 1718.630 2804.600 ;
        RECT 1712.430 2794.625 1712.730 2800.000 ;
        RECT 1712.415 2794.295 1712.745 2794.625 ;
        RECT 1713.350 2787.825 1713.650 2800.000 ;
        RECT 1717.950 2799.750 1718.630 2800.050 ;
        RECT 1718.950 2801.750 1719.250 2804.600 ;
        RECT 1724.170 2801.750 1724.470 2804.600 ;
        RECT 1718.950 2801.450 1720.090 2801.750 ;
        RECT 1718.950 2800.000 1719.250 2801.450 ;
        RECT 1717.950 2794.625 1718.250 2799.750 ;
        RECT 1717.935 2794.295 1718.265 2794.625 ;
        RECT 1719.790 2787.825 1720.090 2801.450 ;
        RECT 1723.470 2801.450 1724.470 2801.750 ;
        RECT 1723.470 2794.625 1723.770 2801.450 ;
        RECT 1724.170 2800.000 1724.470 2801.450 ;
        RECT 1724.790 2796.650 1725.090 2804.600 ;
        RECT 1730.010 2801.750 1730.310 2804.600 ;
        RECT 1724.390 2796.350 1725.090 2796.650 ;
        RECT 1728.990 2801.450 1730.310 2801.750 ;
        RECT 1723.455 2794.295 1723.785 2794.625 ;
        RECT 1724.390 2788.505 1724.690 2796.350 ;
        RECT 1728.990 2794.625 1729.290 2801.450 ;
        RECT 1730.010 2800.000 1730.310 2801.450 ;
        RECT 1730.630 2801.750 1730.930 2804.600 ;
        RECT 1735.850 2802.450 1736.150 2804.600 ;
        RECT 1734.510 2802.150 1736.150 2802.450 ;
        RECT 1730.630 2800.000 1731.130 2801.750 ;
        RECT 1728.975 2794.295 1729.305 2794.625 ;
        RECT 1724.375 2788.175 1724.705 2788.505 ;
        RECT 1730.830 2787.825 1731.130 2800.000 ;
        RECT 1734.510 2794.625 1734.810 2802.150 ;
        RECT 1735.850 2800.000 1736.150 2802.150 ;
        RECT 1736.470 2801.750 1736.770 2804.600 ;
        RECT 1741.690 2801.750 1741.990 2804.600 ;
        RECT 1736.470 2801.450 1737.570 2801.750 ;
        RECT 1736.470 2800.000 1736.770 2801.450 ;
        RECT 1734.495 2794.295 1734.825 2794.625 ;
        RECT 1737.270 2787.825 1737.570 2801.450 ;
        RECT 1740.950 2801.450 1741.990 2801.750 ;
        RECT 1740.950 2794.625 1741.250 2801.450 ;
        RECT 1741.690 2800.000 1741.990 2801.450 ;
        RECT 1742.310 2802.450 1742.610 2804.600 ;
        RECT 1742.310 2802.150 1744.010 2802.450 ;
        RECT 1742.310 2800.000 1742.610 2802.150 ;
        RECT 1740.935 2794.295 1741.265 2794.625 ;
        RECT 1743.710 2787.825 1744.010 2802.150 ;
        RECT 1747.530 2801.750 1747.830 2804.600 ;
        RECT 1747.390 2800.000 1747.830 2801.750 ;
        RECT 1748.150 2801.750 1748.450 2804.600 ;
        RECT 1748.150 2800.000 1748.610 2801.750 ;
        RECT 1753.370 2800.050 1753.670 2804.600 ;
        RECT 1747.390 2794.625 1747.690 2800.000 ;
        RECT 1747.375 2794.295 1747.705 2794.625 ;
        RECT 1748.310 2787.825 1748.610 2800.000 ;
        RECT 1752.910 2799.750 1753.670 2800.050 ;
        RECT 1753.990 2801.750 1754.290 2804.600 ;
        RECT 1753.990 2801.450 1755.050 2801.750 ;
        RECT 1753.990 2800.000 1754.290 2801.450 ;
        RECT 1752.910 2792.585 1753.210 2799.750 ;
        RECT 1752.895 2792.255 1753.225 2792.585 ;
        RECT 1754.750 2787.825 1755.050 2801.450 ;
        RECT 1759.210 2796.665 1759.510 2804.600 ;
        RECT 1759.830 2802.450 1760.130 2804.600 ;
        RECT 1759.830 2802.150 1761.490 2802.450 ;
        RECT 1759.830 2800.000 1760.130 2802.150 ;
        RECT 1759.210 2796.350 1759.665 2796.665 ;
        RECT 1759.335 2796.335 1759.665 2796.350 ;
        RECT 1761.190 2795.985 1761.490 2802.150 ;
        RECT 1765.050 2801.750 1765.350 2804.600 ;
        RECT 1762.110 2801.450 1765.350 2801.750 ;
        RECT 1761.175 2795.655 1761.505 2795.985 ;
        RECT 1762.110 2791.225 1762.410 2801.450 ;
        RECT 1765.050 2800.000 1765.350 2801.450 ;
        RECT 1765.670 2801.750 1765.970 2804.600 ;
        RECT 1770.890 2801.750 1771.190 2804.600 ;
        RECT 1765.670 2800.000 1766.090 2801.750 ;
        RECT 1762.095 2790.895 1762.425 2791.225 ;
        RECT 1765.790 2790.545 1766.090 2800.000 ;
        RECT 1767.630 2801.450 1771.190 2801.750 ;
        RECT 1767.630 2793.945 1767.930 2801.450 ;
        RECT 1770.890 2800.000 1771.190 2801.450 ;
        RECT 1771.510 2801.750 1771.810 2804.600 ;
        RECT 1776.730 2801.750 1777.030 2804.600 ;
        RECT 1771.510 2801.450 1772.530 2801.750 ;
        RECT 1771.510 2800.000 1771.810 2801.450 ;
        RECT 1767.615 2793.615 1767.945 2793.945 ;
        RECT 1765.775 2790.215 1766.105 2790.545 ;
        RECT 1772.230 2789.865 1772.530 2801.450 ;
        RECT 1774.070 2801.450 1777.030 2801.750 ;
        RECT 1774.070 2793.945 1774.370 2801.450 ;
        RECT 1776.730 2800.000 1777.030 2801.450 ;
        RECT 1777.350 2802.450 1777.650 2804.600 ;
        RECT 1777.350 2802.150 1778.970 2802.450 ;
        RECT 1777.350 2800.000 1777.650 2802.150 ;
        RECT 1774.055 2793.615 1774.385 2793.945 ;
        RECT 1778.670 2791.225 1778.970 2802.150 ;
        RECT 1782.570 2801.750 1782.870 2804.600 ;
        RECT 1780.510 2801.450 1782.870 2801.750 ;
        RECT 1780.510 2793.945 1780.810 2801.450 ;
        RECT 1782.570 2800.000 1782.870 2801.450 ;
        RECT 1783.190 2801.750 1783.490 2804.600 ;
        RECT 1783.190 2800.000 1783.570 2801.750 ;
        RECT 1788.410 2800.050 1788.710 2804.600 ;
        RECT 1780.495 2793.615 1780.825 2793.945 ;
        RECT 1778.655 2790.895 1778.985 2791.225 ;
        RECT 1772.215 2789.535 1772.545 2789.865 ;
        RECT 1783.270 2788.505 1783.570 2800.000 ;
        RECT 1787.870 2799.750 1788.710 2800.050 ;
        RECT 1789.030 2801.750 1789.330 2804.600 ;
        RECT 1789.030 2801.450 1790.010 2801.750 ;
        RECT 1789.030 2800.000 1789.330 2801.450 ;
        RECT 1787.870 2792.585 1788.170 2799.750 ;
        RECT 1789.710 2793.265 1790.010 2801.450 ;
        RECT 1794.250 2799.385 1794.550 2804.600 ;
        RECT 1794.870 2803.450 1795.170 2804.600 ;
        RECT 1794.870 2803.150 1797.370 2803.450 ;
        RECT 1794.870 2800.000 1795.170 2803.150 ;
        RECT 1794.235 2799.055 1794.565 2799.385 ;
        RECT 1797.070 2798.705 1797.370 2803.150 ;
        RECT 1794.295 2798.375 1794.625 2798.705 ;
        RECT 1797.055 2798.375 1797.385 2798.705 ;
        RECT 1794.310 2794.625 1794.610 2798.375 ;
        RECT 1794.295 2794.295 1794.625 2794.625 ;
        RECT 1789.695 2792.935 1790.025 2793.265 ;
        RECT 1787.855 2792.255 1788.185 2792.585 ;
        RECT 1783.255 2788.175 1783.585 2788.505 ;
        RECT 1708.735 2787.495 1709.065 2787.825 ;
        RECT 1713.335 2787.495 1713.665 2787.825 ;
        RECT 1719.775 2787.495 1720.105 2787.825 ;
        RECT 1730.815 2787.495 1731.145 2787.825 ;
        RECT 1737.255 2787.495 1737.585 2787.825 ;
        RECT 1743.695 2787.495 1744.025 2787.825 ;
        RECT 1748.295 2787.495 1748.625 2787.825 ;
        RECT 1754.735 2787.495 1755.065 2787.825 ;
        RECT 1644.335 2785.455 1644.665 2785.785 ;
        RECT 1838.455 2069.415 1838.785 2069.745 ;
        RECT 1844.895 2069.415 1845.225 2069.745 ;
        RECT 1851.335 2069.415 1851.665 2069.745 ;
        RECT 1857.775 2069.415 1858.105 2069.745 ;
        RECT 1863.295 2069.415 1863.625 2069.745 ;
        RECT 1869.735 2069.415 1870.065 2069.745 ;
        RECT 1879.855 2069.415 1880.185 2069.745 ;
        RECT 1886.295 2069.415 1886.625 2069.745 ;
        RECT 1891.815 2069.415 1892.145 2069.745 ;
        RECT 1898.255 2069.415 1898.585 2069.745 ;
        RECT 1904.695 2069.415 1905.025 2069.745 ;
        RECT 1911.135 2069.415 1911.465 2069.745 ;
        RECT 1925.855 2069.415 1926.185 2069.745 ;
        RECT 1838.470 2055.450 1838.770 2069.415 ;
        RECT 1841.215 2066.695 1841.545 2067.025 ;
        RECT 1841.230 2058.850 1841.530 2066.695 ;
        RECT 1841.230 2058.550 1842.230 2058.850 ;
        RECT 1841.310 2055.450 1841.610 2056.235 ;
        RECT 1838.470 2055.150 1841.610 2055.450 ;
        RECT 1841.310 2051.635 1841.610 2055.150 ;
        RECT 1841.930 2051.635 1842.230 2058.550 ;
        RECT 1844.910 2055.450 1845.210 2069.415 ;
        RECT 1848.575 2066.695 1848.905 2067.025 ;
        RECT 1847.150 2055.450 1847.450 2056.235 ;
        RECT 1844.910 2055.150 1847.450 2055.450 ;
        RECT 1847.150 2051.635 1847.450 2055.150 ;
        RECT 1847.770 2055.450 1848.070 2056.235 ;
        RECT 1848.590 2055.450 1848.890 2066.695 ;
        RECT 1847.770 2055.150 1848.890 2055.450 ;
        RECT 1851.350 2055.450 1851.650 2069.415 ;
        RECT 1855.015 2066.015 1855.345 2066.345 ;
        RECT 1852.990 2055.450 1853.290 2056.235 ;
        RECT 1851.350 2055.150 1853.290 2055.450 ;
        RECT 1847.770 2051.635 1848.070 2055.150 ;
        RECT 1852.990 2051.635 1853.290 2055.150 ;
        RECT 1853.610 2055.450 1853.910 2056.235 ;
        RECT 1855.030 2055.450 1855.330 2066.015 ;
        RECT 1853.610 2055.150 1855.330 2055.450 ;
        RECT 1857.790 2055.450 1858.090 2069.415 ;
        RECT 1859.615 2065.335 1859.945 2065.665 ;
        RECT 1859.630 2056.235 1859.930 2065.335 ;
        RECT 1858.830 2055.450 1859.130 2056.235 ;
        RECT 1857.790 2055.150 1859.130 2055.450 ;
        RECT 1853.610 2051.635 1853.910 2055.150 ;
        RECT 1858.830 2051.635 1859.130 2055.150 ;
        RECT 1859.450 2055.150 1859.930 2056.235 ;
        RECT 1859.450 2051.635 1859.750 2055.150 ;
        RECT 1863.310 2053.750 1863.610 2069.415 ;
        RECT 1865.135 2065.335 1865.465 2065.665 ;
        RECT 1865.150 2058.850 1865.450 2065.335 ;
        RECT 1865.150 2058.550 1865.590 2058.850 ;
        RECT 1864.670 2053.750 1864.970 2056.235 ;
        RECT 1863.310 2053.450 1864.970 2053.750 ;
        RECT 1864.670 2051.635 1864.970 2053.450 ;
        RECT 1865.290 2051.635 1865.590 2058.550 ;
        RECT 1869.750 2055.450 1870.050 2069.415 ;
        RECT 1873.415 2068.735 1873.745 2069.065 ;
        RECT 1871.575 2064.655 1871.905 2064.985 ;
        RECT 1871.590 2058.850 1871.890 2064.655 ;
        RECT 1871.130 2058.550 1871.890 2058.850 ;
        RECT 1870.510 2055.450 1870.810 2056.235 ;
        RECT 1869.750 2055.150 1870.810 2055.450 ;
        RECT 1870.510 2051.635 1870.810 2055.150 ;
        RECT 1871.130 2051.635 1871.430 2058.550 ;
        RECT 1873.430 2055.450 1873.730 2068.735 ;
        RECT 1877.095 2063.975 1877.425 2064.305 ;
        RECT 1877.110 2056.235 1877.410 2063.975 ;
        RECT 1876.350 2055.450 1876.650 2056.235 ;
        RECT 1873.430 2055.150 1876.650 2055.450 ;
        RECT 1876.350 2051.635 1876.650 2055.150 ;
        RECT 1876.970 2055.150 1877.410 2056.235 ;
        RECT 1879.870 2055.450 1880.170 2069.415 ;
        RECT 1882.615 2063.975 1882.945 2064.305 ;
        RECT 1882.630 2058.850 1882.930 2063.975 ;
        RECT 1882.630 2058.550 1883.110 2058.850 ;
        RECT 1882.190 2055.450 1882.490 2056.235 ;
        RECT 1879.870 2055.150 1882.490 2055.450 ;
        RECT 1876.970 2051.635 1877.270 2055.150 ;
        RECT 1882.190 2051.635 1882.490 2055.150 ;
        RECT 1882.810 2051.635 1883.110 2058.550 ;
        RECT 1886.310 2055.450 1886.610 2069.415 ;
        RECT 1889.975 2066.695 1890.305 2067.025 ;
        RECT 1888.030 2055.450 1888.330 2056.235 ;
        RECT 1886.310 2055.150 1888.330 2055.450 ;
        RECT 1888.030 2051.635 1888.330 2055.150 ;
        RECT 1888.650 2055.450 1888.950 2056.235 ;
        RECT 1889.990 2055.450 1890.290 2066.695 ;
        RECT 1888.650 2055.150 1890.290 2055.450 ;
        RECT 1891.830 2055.450 1892.130 2069.415 ;
        RECT 1894.575 2065.335 1894.905 2065.665 ;
        RECT 1894.590 2056.235 1894.890 2065.335 ;
        RECT 1893.870 2055.450 1894.170 2056.235 ;
        RECT 1891.830 2055.150 1894.170 2055.450 ;
        RECT 1888.650 2051.635 1888.950 2055.150 ;
        RECT 1893.870 2051.635 1894.170 2055.150 ;
        RECT 1894.490 2055.150 1894.890 2056.235 ;
        RECT 1898.270 2055.450 1898.570 2069.415 ;
        RECT 1901.015 2066.015 1901.345 2066.345 ;
        RECT 1899.710 2055.450 1900.010 2056.235 ;
        RECT 1898.270 2055.150 1900.010 2055.450 ;
        RECT 1894.490 2051.635 1894.790 2055.150 ;
        RECT 1899.710 2051.635 1900.010 2055.150 ;
        RECT 1900.330 2055.450 1900.630 2056.235 ;
        RECT 1901.030 2055.450 1901.330 2066.015 ;
        RECT 1900.330 2055.150 1901.330 2055.450 ;
        RECT 1904.710 2055.450 1905.010 2069.415 ;
        RECT 1907.455 2065.335 1907.785 2065.665 ;
        RECT 1905.550 2055.450 1905.850 2056.235 ;
        RECT 1904.710 2055.150 1905.850 2055.450 ;
        RECT 1900.330 2051.635 1900.630 2055.150 ;
        RECT 1905.550 2051.635 1905.850 2055.150 ;
        RECT 1906.170 2055.450 1906.470 2056.235 ;
        RECT 1907.470 2055.450 1907.770 2065.335 ;
        RECT 1906.170 2055.150 1907.770 2055.450 ;
        RECT 1911.150 2056.235 1911.450 2069.415 ;
        RECT 1914.815 2068.735 1915.145 2069.065 ;
        RECT 1920.335 2068.735 1920.665 2069.065 ;
        RECT 1912.055 2065.335 1912.385 2065.665 ;
        RECT 1912.070 2056.235 1912.370 2065.335 ;
        RECT 1911.150 2055.150 1911.690 2056.235 ;
        RECT 1906.170 2051.635 1906.470 2055.150 ;
        RECT 1911.390 2051.635 1911.690 2055.150 ;
        RECT 1912.010 2055.150 1912.370 2056.235 ;
        RECT 1914.830 2055.450 1915.130 2068.735 ;
        RECT 1917.575 2064.655 1917.905 2064.985 ;
        RECT 1917.590 2058.850 1917.890 2064.655 ;
        RECT 1917.590 2058.550 1918.150 2058.850 ;
        RECT 1917.230 2055.450 1917.530 2056.235 ;
        RECT 1914.830 2055.150 1917.530 2055.450 ;
        RECT 1912.010 2051.635 1912.310 2055.150 ;
        RECT 1917.230 2051.635 1917.530 2055.150 ;
        RECT 1917.850 2051.635 1918.150 2058.550 ;
        RECT 1920.350 2055.450 1920.650 2068.735 ;
        RECT 1924.015 2064.655 1924.345 2064.985 ;
        RECT 1924.030 2058.850 1924.330 2064.655 ;
        RECT 1923.690 2058.550 1924.330 2058.850 ;
        RECT 1923.070 2055.450 1923.370 2056.235 ;
        RECT 1920.350 2055.150 1923.370 2055.450 ;
        RECT 1923.070 2051.635 1923.370 2055.150 ;
        RECT 1923.690 2051.635 1923.990 2058.550 ;
        RECT 1925.870 2055.450 1926.170 2069.415 ;
        RECT 1981.975 2068.055 1982.305 2068.385 ;
        RECT 1987.495 2068.055 1987.825 2068.385 ;
        RECT 1941.495 2066.695 1941.825 2067.025 ;
        RECT 1934.135 2066.015 1934.465 2066.345 ;
        RECT 1929.535 2064.655 1929.865 2064.985 ;
        RECT 1929.550 2056.235 1929.850 2064.655 ;
        RECT 1928.910 2055.450 1929.210 2056.235 ;
        RECT 1925.870 2055.150 1929.210 2055.450 ;
        RECT 1928.910 2051.635 1929.210 2055.150 ;
        RECT 1929.530 2055.150 1929.850 2056.235 ;
        RECT 1934.150 2055.450 1934.450 2066.015 ;
        RECT 1935.975 2065.335 1936.305 2065.665 ;
        RECT 1934.750 2055.450 1935.050 2056.235 ;
        RECT 1934.150 2055.150 1935.050 2055.450 ;
        RECT 1929.530 2051.635 1929.830 2055.150 ;
        RECT 1934.750 2051.635 1935.050 2055.150 ;
        RECT 1935.370 2055.450 1935.670 2056.235 ;
        RECT 1935.990 2055.450 1936.290 2065.335 ;
        RECT 1940.575 2058.535 1940.905 2058.865 ;
        RECT 1935.370 2055.150 1936.290 2055.450 ;
        RECT 1935.370 2051.635 1935.670 2055.150 ;
        RECT 1940.590 2051.635 1940.890 2058.535 ;
        RECT 1941.510 2056.235 1941.810 2066.695 ;
        RECT 1967.255 2063.975 1967.585 2064.305 ;
        RECT 1947.935 2063.295 1948.265 2063.625 ;
        RECT 1954.375 2063.295 1954.705 2063.625 ;
        RECT 1958.975 2063.295 1959.305 2063.625 ;
        RECT 1965.415 2063.295 1965.745 2063.625 ;
        RECT 1946.415 2057.175 1946.745 2057.505 ;
        RECT 1941.210 2055.150 1941.810 2056.235 ;
        RECT 1941.210 2051.635 1941.510 2055.150 ;
        RECT 1946.430 2051.635 1946.730 2057.175 ;
        RECT 1947.050 2055.450 1947.350 2056.235 ;
        RECT 1947.950 2055.450 1948.250 2063.295 ;
        RECT 1947.050 2055.150 1948.250 2055.450 ;
        RECT 1948.855 2055.450 1949.185 2055.465 ;
        RECT 1952.270 2055.450 1952.570 2056.235 ;
        RECT 1948.855 2055.150 1952.570 2055.450 ;
        RECT 1947.050 2051.635 1947.350 2055.150 ;
        RECT 1948.855 2055.135 1949.185 2055.150 ;
        RECT 1952.270 2051.635 1952.570 2055.150 ;
        RECT 1952.890 2053.750 1953.190 2056.235 ;
        RECT 1954.390 2053.750 1954.690 2063.295 ;
        RECT 1955.295 2057.855 1955.625 2058.185 ;
        RECT 1955.310 2055.450 1955.610 2057.855 ;
        RECT 1958.990 2056.235 1959.290 2063.295 ;
        RECT 1958.110 2055.450 1958.410 2056.235 ;
        RECT 1955.310 2055.150 1958.410 2055.450 ;
        RECT 1952.890 2053.450 1954.690 2053.750 ;
        RECT 1952.890 2051.635 1953.190 2053.450 ;
        RECT 1958.110 2051.635 1958.410 2055.150 ;
        RECT 1958.730 2055.150 1959.290 2056.235 ;
        RECT 1958.730 2051.635 1959.030 2055.150 ;
        RECT 1961.505 2052.050 1961.835 2052.065 ;
        RECT 1963.950 2052.050 1964.250 2056.235 ;
        RECT 1961.505 2051.750 1964.250 2052.050 ;
        RECT 1961.505 2051.735 1961.835 2051.750 ;
        RECT 1963.950 2051.635 1964.250 2051.750 ;
        RECT 1964.570 2055.450 1964.870 2056.235 ;
        RECT 1965.430 2055.450 1965.730 2063.295 ;
        RECT 1964.570 2055.150 1965.730 2055.450 ;
        RECT 1967.270 2055.450 1967.570 2063.975 ;
        RECT 1970.015 2063.295 1970.345 2063.625 ;
        RECT 1973.695 2063.295 1974.025 2063.625 ;
        RECT 1976.455 2063.295 1976.785 2063.625 ;
        RECT 1980.135 2063.295 1980.465 2063.625 ;
        RECT 1970.030 2058.170 1970.330 2063.295 ;
        RECT 1970.030 2057.870 1970.710 2058.170 ;
        RECT 1969.790 2055.450 1970.090 2056.235 ;
        RECT 1967.270 2055.150 1970.090 2055.450 ;
        RECT 1964.570 2051.635 1964.870 2055.150 ;
        RECT 1969.790 2051.635 1970.090 2055.150 ;
        RECT 1970.410 2051.635 1970.710 2057.870 ;
        RECT 1973.710 2055.450 1974.010 2063.295 ;
        RECT 1976.470 2056.235 1976.770 2063.295 ;
        RECT 1975.630 2055.450 1975.930 2056.235 ;
        RECT 1973.710 2055.150 1975.930 2055.450 ;
        RECT 1975.630 2051.635 1975.930 2055.150 ;
        RECT 1976.250 2055.150 1976.770 2056.235 ;
        RECT 1976.250 2051.635 1976.550 2055.150 ;
        RECT 1980.150 2053.750 1980.450 2063.295 ;
        RECT 1981.990 2058.170 1982.290 2068.055 ;
        RECT 1987.510 2058.850 1987.810 2068.055 ;
        RECT 2028.895 2067.375 2029.225 2067.705 ;
        RECT 2023.375 2066.695 2023.705 2067.025 ;
        RECT 2011.415 2066.015 2011.745 2066.345 ;
        RECT 2016.935 2066.015 2017.265 2066.345 ;
        RECT 1999.455 2065.335 1999.785 2065.665 ;
        RECT 1993.015 2063.975 1993.345 2064.305 ;
        RECT 1987.510 2058.550 1988.230 2058.850 ;
        RECT 1981.990 2057.870 1982.390 2058.170 ;
        RECT 1981.470 2053.750 1981.770 2056.235 ;
        RECT 1980.150 2053.450 1981.770 2053.750 ;
        RECT 1981.470 2051.635 1981.770 2053.450 ;
        RECT 1982.090 2051.635 1982.390 2057.870 ;
        RECT 1987.295 2057.855 1987.625 2058.185 ;
        RECT 1987.310 2051.635 1987.610 2057.855 ;
        RECT 1987.930 2051.635 1988.230 2058.550 ;
        RECT 1993.030 2058.170 1993.330 2063.975 ;
        RECT 1993.030 2057.870 1994.070 2058.170 ;
        RECT 1990.255 2057.175 1990.585 2057.505 ;
        RECT 1990.270 2055.450 1990.570 2057.175 ;
        RECT 1993.150 2055.450 1993.450 2056.235 ;
        RECT 1990.270 2055.150 1993.450 2055.450 ;
        RECT 1993.150 2051.635 1993.450 2055.150 ;
        RECT 1993.770 2051.635 1994.070 2057.870 ;
        RECT 1995.775 2057.855 1996.105 2058.185 ;
        RECT 1995.790 2055.450 1996.090 2057.855 ;
        RECT 1999.470 2057.490 1999.770 2065.335 ;
        RECT 2005.895 2064.655 2006.225 2064.985 ;
        RECT 1999.470 2057.190 1999.910 2057.490 ;
        RECT 1998.990 2055.450 1999.290 2056.235 ;
        RECT 1995.790 2055.150 1999.290 2055.450 ;
        RECT 1998.990 2051.635 1999.290 2055.150 ;
        RECT 1999.610 2051.635 1999.910 2057.190 ;
        RECT 2004.815 2057.175 2005.145 2057.505 ;
        RECT 2005.910 2057.490 2006.210 2064.655 ;
        RECT 2005.450 2057.190 2006.210 2057.490 ;
        RECT 2004.830 2051.635 2005.130 2057.175 ;
        RECT 2005.450 2051.635 2005.750 2057.190 ;
        RECT 2008.655 2056.495 2008.985 2056.825 ;
        RECT 2008.670 2055.450 2008.970 2056.495 ;
        RECT 2011.430 2056.235 2011.730 2066.015 ;
        RECT 2016.950 2058.850 2017.250 2066.015 ;
        RECT 2023.390 2058.850 2023.690 2066.695 ;
        RECT 2016.950 2058.550 2017.430 2058.850 ;
        RECT 2016.495 2057.175 2016.825 2057.505 ;
        RECT 2010.670 2055.450 2010.970 2056.235 ;
        RECT 2008.670 2055.150 2010.970 2055.450 ;
        RECT 2010.670 2051.635 2010.970 2055.150 ;
        RECT 2011.290 2055.150 2011.730 2056.235 ;
        RECT 2011.290 2051.635 2011.590 2055.150 ;
        RECT 2016.510 2051.635 2016.810 2057.175 ;
        RECT 2017.130 2051.635 2017.430 2058.550 ;
        RECT 2022.970 2058.550 2023.690 2058.850 ;
        RECT 2021.535 2056.495 2021.865 2056.825 ;
        RECT 2021.550 2055.450 2021.850 2056.495 ;
        RECT 2022.350 2055.450 2022.650 2056.235 ;
        RECT 2021.550 2055.150 2022.650 2055.450 ;
        RECT 2022.350 2051.635 2022.650 2055.150 ;
        RECT 2022.970 2051.635 2023.270 2058.550 ;
        RECT 2028.910 2056.235 2029.210 2067.375 ;
        RECT 2037.175 2066.015 2037.505 2066.345 ;
        RECT 2031.655 2063.295 2031.985 2063.625 ;
        RECT 2028.810 2055.150 2029.210 2056.235 ;
        RECT 2031.670 2055.450 2031.970 2063.295 ;
        RECT 2034.650 2055.450 2034.950 2056.235 ;
        RECT 2031.670 2055.150 2034.950 2055.450 ;
        RECT 2037.190 2055.450 2037.490 2066.015 ;
        RECT 2043.615 2065.335 2043.945 2065.665 ;
        RECT 2040.490 2055.450 2040.790 2056.235 ;
        RECT 2037.190 2055.150 2040.790 2055.450 ;
        RECT 2043.630 2055.450 2043.930 2065.335 ;
        RECT 2046.330 2055.450 2046.630 2056.235 ;
        RECT 2043.630 2055.150 2046.630 2055.450 ;
        RECT 2028.810 2051.635 2029.110 2055.150 ;
        RECT 2034.650 2051.635 2034.950 2055.150 ;
        RECT 2040.490 2051.635 2040.790 2055.150 ;
        RECT 2046.330 2051.635 2046.630 2055.150 ;
        RECT 2050.055 2052.050 2050.385 2052.065 ;
        RECT 2052.170 2052.050 2052.470 2056.235 ;
        RECT 2050.055 2051.750 2052.470 2052.050 ;
        RECT 2050.055 2051.735 2050.385 2051.750 ;
        RECT 2052.170 2051.635 2052.470 2051.750 ;
        RECT 1418.935 1980.335 1419.265 1980.665 ;
        RECT 1417.095 1975.575 1417.425 1975.905 ;
        RECT 1411.575 1955.175 1411.905 1955.505 ;
      LAYER met4 ;
        RECT 323.295 1606.975 1389.905 1610.240 ;
        RECT 1705.000 1605.000 2081.480 2051.235 ;
      LAYER met4 ;
        RECT 1718.315 1602.450 1718.615 1604.600 ;
        RECT 1718.315 1602.150 1720.090 1602.450 ;
        RECT 1718.315 1600.000 1718.615 1602.150 ;
        RECT 1719.790 1593.745 1720.090 1602.150 ;
        RECT 1743.290 1601.550 1743.590 1604.600 ;
        RECT 1740.030 1601.250 1743.590 1601.550 ;
        RECT 1719.775 1593.415 1720.105 1593.745 ;
        RECT 1740.030 1592.385 1740.330 1601.250 ;
        RECT 1743.290 1600.000 1743.590 1601.250 ;
        RECT 1798.715 1600.000 1799.015 1604.600 ;
        RECT 1804.955 1600.000 1805.255 1604.600 ;
        RECT 1811.195 1600.000 1811.495 1604.600 ;
        RECT 1817.435 1600.000 1817.735 1604.600 ;
        RECT 1823.675 1600.000 1823.975 1604.600 ;
        RECT 1829.915 1600.000 1830.215 1604.600 ;
        RECT 1836.155 1600.000 1836.455 1604.600 ;
        RECT 1842.395 1600.000 1842.695 1604.600 ;
        RECT 1848.635 1600.000 1848.935 1604.600 ;
        RECT 1854.875 1600.000 1855.175 1604.600 ;
        RECT 1861.115 1600.000 1861.415 1604.600 ;
        RECT 1867.355 1600.000 1867.655 1604.600 ;
        RECT 1873.595 1600.000 1873.895 1604.600 ;
        RECT 1879.835 1600.000 1880.135 1604.600 ;
        RECT 1886.075 1600.000 1886.375 1604.600 ;
        RECT 1892.315 1600.000 1892.615 1604.600 ;
        RECT 1898.555 1600.000 1898.855 1604.600 ;
        RECT 1904.795 1600.000 1905.095 1604.600 ;
        RECT 1911.035 1600.000 1911.335 1604.600 ;
        RECT 1917.275 1600.000 1917.575 1604.600 ;
        RECT 1923.515 1600.000 1923.815 1604.600 ;
        RECT 1929.755 1600.000 1930.055 1604.600 ;
        RECT 1935.995 1600.000 1936.295 1604.600 ;
        RECT 1942.235 1600.000 1942.535 1604.600 ;
        RECT 1948.475 1600.000 1948.775 1604.600 ;
        RECT 1954.715 1600.000 1955.015 1604.600 ;
        RECT 1960.955 1600.000 1961.255 1604.600 ;
        RECT 1967.195 1600.000 1967.495 1604.600 ;
        RECT 1973.435 1600.000 1973.735 1604.600 ;
        RECT 1979.675 1600.000 1979.975 1604.600 ;
        RECT 1985.915 1600.000 1986.215 1604.600 ;
        RECT 1992.155 1600.000 1992.455 1604.600 ;
        RECT 1740.015 1592.055 1740.345 1592.385 ;
  END
END user_project_wrapper
END LIBRARY

