VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO hs32_core1
  CLASS BLOCK ;
  FOREIGN hs32_core1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1200.000 BY 1200.000 ;
  PIN cpu_addr_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 489.640 1200.000 490.240 ;
    END
  END cpu_addr_e[0]
  PIN cpu_addr_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 599.800 1200.000 600.400 ;
    END
  END cpu_addr_e[10]
  PIN cpu_addr_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 610.680 1200.000 611.280 ;
    END
  END cpu_addr_e[11]
  PIN cpu_addr_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 621.560 1200.000 622.160 ;
    END
  END cpu_addr_e[12]
  PIN cpu_addr_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 632.440 1200.000 633.040 ;
    END
  END cpu_addr_e[13]
  PIN cpu_addr_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 644.000 1200.000 644.600 ;
    END
  END cpu_addr_e[14]
  PIN cpu_addr_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 654.880 1200.000 655.480 ;
    END
  END cpu_addr_e[15]
  PIN cpu_addr_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 500.520 1200.000 501.120 ;
    END
  END cpu_addr_e[1]
  PIN cpu_addr_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 511.400 1200.000 512.000 ;
    END
  END cpu_addr_e[2]
  PIN cpu_addr_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 522.960 1200.000 523.560 ;
    END
  END cpu_addr_e[3]
  PIN cpu_addr_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 533.840 1200.000 534.440 ;
    END
  END cpu_addr_e[4]
  PIN cpu_addr_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 544.720 1200.000 545.320 ;
    END
  END cpu_addr_e[5]
  PIN cpu_addr_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 555.600 1200.000 556.200 ;
    END
  END cpu_addr_e[6]
  PIN cpu_addr_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 566.480 1200.000 567.080 ;
    END
  END cpu_addr_e[7]
  PIN cpu_addr_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 578.040 1200.000 578.640 ;
    END
  END cpu_addr_e[8]
  PIN cpu_addr_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 588.920 1200.000 589.520 ;
    END
  END cpu_addr_e[9]
  PIN cpu_addr_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 367.630 1196.000 367.910 1200.000 ;
    END
  END cpu_addr_n[0]
  PIN cpu_addr_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 480.790 1196.000 481.070 1200.000 ;
    END
  END cpu_addr_n[10]
  PIN cpu_addr_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.290 1196.000 492.570 1200.000 ;
    END
  END cpu_addr_n[11]
  PIN cpu_addr_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 1196.000 503.610 1200.000 ;
    END
  END cpu_addr_n[12]
  PIN cpu_addr_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.830 1196.000 515.110 1200.000 ;
    END
  END cpu_addr_n[13]
  PIN cpu_addr_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.330 1196.000 526.610 1200.000 ;
    END
  END cpu_addr_n[14]
  PIN cpu_addr_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.370 1196.000 537.650 1200.000 ;
    END
  END cpu_addr_n[15]
  PIN cpu_addr_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.130 1196.000 379.410 1200.000 ;
    END
  END cpu_addr_n[1]
  PIN cpu_addr_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 390.170 1196.000 390.450 1200.000 ;
    END
  END cpu_addr_n[2]
  PIN cpu_addr_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.670 1196.000 401.950 1200.000 ;
    END
  END cpu_addr_n[3]
  PIN cpu_addr_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 413.170 1196.000 413.450 1200.000 ;
    END
  END cpu_addr_n[4]
  PIN cpu_addr_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.210 1196.000 424.490 1200.000 ;
    END
  END cpu_addr_n[5]
  PIN cpu_addr_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.710 1196.000 435.990 1200.000 ;
    END
  END cpu_addr_n[6]
  PIN cpu_addr_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.750 1196.000 447.030 1200.000 ;
    END
  END cpu_addr_n[7]
  PIN cpu_addr_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 458.250 1196.000 458.530 1200.000 ;
    END
  END cpu_addr_n[8]
  PIN cpu_addr_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 469.750 1196.000 470.030 1200.000 ;
    END
  END cpu_addr_n[9]
  PIN cpu_dtr_e0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 27.240 1200.000 27.840 ;
    END
  END cpu_dtr_e0[0]
  PIN cpu_dtr_e0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 137.400 1200.000 138.000 ;
    END
  END cpu_dtr_e0[10]
  PIN cpu_dtr_e0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 148.280 1200.000 148.880 ;
    END
  END cpu_dtr_e0[11]
  PIN cpu_dtr_e0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 159.160 1200.000 159.760 ;
    END
  END cpu_dtr_e0[12]
  PIN cpu_dtr_e0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 170.040 1200.000 170.640 ;
    END
  END cpu_dtr_e0[13]
  PIN cpu_dtr_e0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 181.600 1200.000 182.200 ;
    END
  END cpu_dtr_e0[14]
  PIN cpu_dtr_e0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 192.480 1200.000 193.080 ;
    END
  END cpu_dtr_e0[15]
  PIN cpu_dtr_e0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 203.360 1200.000 203.960 ;
    END
  END cpu_dtr_e0[16]
  PIN cpu_dtr_e0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 214.240 1200.000 214.840 ;
    END
  END cpu_dtr_e0[17]
  PIN cpu_dtr_e0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 225.120 1200.000 225.720 ;
    END
  END cpu_dtr_e0[18]
  PIN cpu_dtr_e0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 236.680 1200.000 237.280 ;
    END
  END cpu_dtr_e0[19]
  PIN cpu_dtr_e0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 38.120 1200.000 38.720 ;
    END
  END cpu_dtr_e0[1]
  PIN cpu_dtr_e0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 247.560 1200.000 248.160 ;
    END
  END cpu_dtr_e0[20]
  PIN cpu_dtr_e0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 258.440 1200.000 259.040 ;
    END
  END cpu_dtr_e0[21]
  PIN cpu_dtr_e0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 269.320 1200.000 269.920 ;
    END
  END cpu_dtr_e0[22]
  PIN cpu_dtr_e0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 280.200 1200.000 280.800 ;
    END
  END cpu_dtr_e0[23]
  PIN cpu_dtr_e0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 291.760 1200.000 292.360 ;
    END
  END cpu_dtr_e0[24]
  PIN cpu_dtr_e0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 302.640 1200.000 303.240 ;
    END
  END cpu_dtr_e0[25]
  PIN cpu_dtr_e0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 313.520 1200.000 314.120 ;
    END
  END cpu_dtr_e0[26]
  PIN cpu_dtr_e0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 324.400 1200.000 325.000 ;
    END
  END cpu_dtr_e0[27]
  PIN cpu_dtr_e0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 335.280 1200.000 335.880 ;
    END
  END cpu_dtr_e0[28]
  PIN cpu_dtr_e0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 346.160 1200.000 346.760 ;
    END
  END cpu_dtr_e0[29]
  PIN cpu_dtr_e0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 49.000 1200.000 49.600 ;
    END
  END cpu_dtr_e0[2]
  PIN cpu_dtr_e0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 357.720 1200.000 358.320 ;
    END
  END cpu_dtr_e0[30]
  PIN cpu_dtr_e0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 368.600 1200.000 369.200 ;
    END
  END cpu_dtr_e0[31]
  PIN cpu_dtr_e0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 59.880 1200.000 60.480 ;
    END
  END cpu_dtr_e0[3]
  PIN cpu_dtr_e0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 71.440 1200.000 72.040 ;
    END
  END cpu_dtr_e0[4]
  PIN cpu_dtr_e0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 82.320 1200.000 82.920 ;
    END
  END cpu_dtr_e0[5]
  PIN cpu_dtr_e0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 93.200 1200.000 93.800 ;
    END
  END cpu_dtr_e0[6]
  PIN cpu_dtr_e0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 104.080 1200.000 104.680 ;
    END
  END cpu_dtr_e0[7]
  PIN cpu_dtr_e0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 114.960 1200.000 115.560 ;
    END
  END cpu_dtr_e0[8]
  PIN cpu_dtr_e0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 126.520 1200.000 127.120 ;
    END
  END cpu_dtr_e0[9]
  PIN cpu_dtr_e1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 841.880 1200.000 842.480 ;
    END
  END cpu_dtr_e1[0]
  PIN cpu_dtr_e1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 952.040 1200.000 952.640 ;
    END
  END cpu_dtr_e1[10]
  PIN cpu_dtr_e1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 962.920 1200.000 963.520 ;
    END
  END cpu_dtr_e1[11]
  PIN cpu_dtr_e1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 973.800 1200.000 974.400 ;
    END
  END cpu_dtr_e1[12]
  PIN cpu_dtr_e1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 985.360 1200.000 985.960 ;
    END
  END cpu_dtr_e1[13]
  PIN cpu_dtr_e1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 996.240 1200.000 996.840 ;
    END
  END cpu_dtr_e1[14]
  PIN cpu_dtr_e1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1007.120 1200.000 1007.720 ;
    END
  END cpu_dtr_e1[15]
  PIN cpu_dtr_e1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1018.000 1200.000 1018.600 ;
    END
  END cpu_dtr_e1[16]
  PIN cpu_dtr_e1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1028.880 1200.000 1029.480 ;
    END
  END cpu_dtr_e1[17]
  PIN cpu_dtr_e1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1040.440 1200.000 1041.040 ;
    END
  END cpu_dtr_e1[18]
  PIN cpu_dtr_e1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1051.320 1200.000 1051.920 ;
    END
  END cpu_dtr_e1[19]
  PIN cpu_dtr_e1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 852.760 1200.000 853.360 ;
    END
  END cpu_dtr_e1[1]
  PIN cpu_dtr_e1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1062.200 1200.000 1062.800 ;
    END
  END cpu_dtr_e1[20]
  PIN cpu_dtr_e1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1073.080 1200.000 1073.680 ;
    END
  END cpu_dtr_e1[21]
  PIN cpu_dtr_e1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1083.960 1200.000 1084.560 ;
    END
  END cpu_dtr_e1[22]
  PIN cpu_dtr_e1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1095.520 1200.000 1096.120 ;
    END
  END cpu_dtr_e1[23]
  PIN cpu_dtr_e1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1106.400 1200.000 1107.000 ;
    END
  END cpu_dtr_e1[24]
  PIN cpu_dtr_e1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1117.280 1200.000 1117.880 ;
    END
  END cpu_dtr_e1[25]
  PIN cpu_dtr_e1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1128.160 1200.000 1128.760 ;
    END
  END cpu_dtr_e1[26]
  PIN cpu_dtr_e1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1139.040 1200.000 1139.640 ;
    END
  END cpu_dtr_e1[27]
  PIN cpu_dtr_e1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1150.600 1200.000 1151.200 ;
    END
  END cpu_dtr_e1[28]
  PIN cpu_dtr_e1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1161.480 1200.000 1162.080 ;
    END
  END cpu_dtr_e1[29]
  PIN cpu_dtr_e1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 864.320 1200.000 864.920 ;
    END
  END cpu_dtr_e1[2]
  PIN cpu_dtr_e1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1172.360 1200.000 1172.960 ;
    END
  END cpu_dtr_e1[30]
  PIN cpu_dtr_e1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1183.240 1200.000 1183.840 ;
    END
  END cpu_dtr_e1[31]
  PIN cpu_dtr_e1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 875.200 1200.000 875.800 ;
    END
  END cpu_dtr_e1[3]
  PIN cpu_dtr_e1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 886.080 1200.000 886.680 ;
    END
  END cpu_dtr_e1[4]
  PIN cpu_dtr_e1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 896.960 1200.000 897.560 ;
    END
  END cpu_dtr_e1[5]
  PIN cpu_dtr_e1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 907.840 1200.000 908.440 ;
    END
  END cpu_dtr_e1[6]
  PIN cpu_dtr_e1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 918.720 1200.000 919.320 ;
    END
  END cpu_dtr_e1[7]
  PIN cpu_dtr_e1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 930.280 1200.000 930.880 ;
    END
  END cpu_dtr_e1[8]
  PIN cpu_dtr_e1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1196.000 941.160 1200.000 941.760 ;
    END
  END cpu_dtr_e1[9]
  PIN cpu_dtr_n0[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.610 1196.000 5.890 1200.000 ;
    END
  END cpu_dtr_n0[0]
  PIN cpu_dtr_n0[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.770 1196.000 119.050 1200.000 ;
    END
  END cpu_dtr_n0[10]
  PIN cpu_dtr_n0[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.810 1196.000 130.090 1200.000 ;
    END
  END cpu_dtr_n0[11]
  PIN cpu_dtr_n0[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.310 1196.000 141.590 1200.000 ;
    END
  END cpu_dtr_n0[12]
  PIN cpu_dtr_n0[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.350 1196.000 152.630 1200.000 ;
    END
  END cpu_dtr_n0[13]
  PIN cpu_dtr_n0[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.850 1196.000 164.130 1200.000 ;
    END
  END cpu_dtr_n0[14]
  PIN cpu_dtr_n0[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.350 1196.000 175.630 1200.000 ;
    END
  END cpu_dtr_n0[15]
  PIN cpu_dtr_n0[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.390 1196.000 186.670 1200.000 ;
    END
  END cpu_dtr_n0[16]
  PIN cpu_dtr_n0[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.890 1196.000 198.170 1200.000 ;
    END
  END cpu_dtr_n0[17]
  PIN cpu_dtr_n0[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.390 1196.000 209.670 1200.000 ;
    END
  END cpu_dtr_n0[18]
  PIN cpu_dtr_n0[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 1196.000 220.710 1200.000 ;
    END
  END cpu_dtr_n0[19]
  PIN cpu_dtr_n0[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 1196.000 16.930 1200.000 ;
    END
  END cpu_dtr_n0[1]
  PIN cpu_dtr_n0[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 231.930 1196.000 232.210 1200.000 ;
    END
  END cpu_dtr_n0[20]
  PIN cpu_dtr_n0[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 1196.000 243.250 1200.000 ;
    END
  END cpu_dtr_n0[21]
  PIN cpu_dtr_n0[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.470 1196.000 254.750 1200.000 ;
    END
  END cpu_dtr_n0[22]
  PIN cpu_dtr_n0[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 265.970 1196.000 266.250 1200.000 ;
    END
  END cpu_dtr_n0[23]
  PIN cpu_dtr_n0[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 1196.000 277.290 1200.000 ;
    END
  END cpu_dtr_n0[24]
  PIN cpu_dtr_n0[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.510 1196.000 288.790 1200.000 ;
    END
  END cpu_dtr_n0[25]
  PIN cpu_dtr_n0[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.550 1196.000 299.830 1200.000 ;
    END
  END cpu_dtr_n0[26]
  PIN cpu_dtr_n0[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.050 1196.000 311.330 1200.000 ;
    END
  END cpu_dtr_n0[27]
  PIN cpu_dtr_n0[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.550 1196.000 322.830 1200.000 ;
    END
  END cpu_dtr_n0[28]
  PIN cpu_dtr_n0[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.590 1196.000 333.870 1200.000 ;
    END
  END cpu_dtr_n0[29]
  PIN cpu_dtr_n0[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.150 1196.000 28.430 1200.000 ;
    END
  END cpu_dtr_n0[2]
  PIN cpu_dtr_n0[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.090 1196.000 345.370 1200.000 ;
    END
  END cpu_dtr_n0[30]
  PIN cpu_dtr_n0[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.590 1196.000 356.870 1200.000 ;
    END
  END cpu_dtr_n0[31]
  PIN cpu_dtr_n0[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.190 1196.000 39.470 1200.000 ;
    END
  END cpu_dtr_n0[3]
  PIN cpu_dtr_n0[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 1196.000 50.970 1200.000 ;
    END
  END cpu_dtr_n0[4]
  PIN cpu_dtr_n0[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 1196.000 62.470 1200.000 ;
    END
  END cpu_dtr_n0[5]
  PIN cpu_dtr_n0[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.230 1196.000 73.510 1200.000 ;
    END
  END cpu_dtr_n0[6]
  PIN cpu_dtr_n0[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 84.730 1196.000 85.010 1200.000 ;
    END
  END cpu_dtr_n0[7]
  PIN cpu_dtr_n0[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 95.770 1196.000 96.050 1200.000 ;
    END
  END cpu_dtr_n0[8]
  PIN cpu_dtr_n0[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.270 1196.000 107.550 1200.000 ;
    END
  END cpu_dtr_n0[9]
  PIN cpu_dtr_n1[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 843.270 1196.000 843.550 1200.000 ;
    END
  END cpu_dtr_n1[0]
  PIN cpu_dtr_n1[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.430 1196.000 956.710 1200.000 ;
    END
  END cpu_dtr_n1[10]
  PIN cpu_dtr_n1[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.930 1196.000 968.210 1200.000 ;
    END
  END cpu_dtr_n1[11]
  PIN cpu_dtr_n1[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.970 1196.000 979.250 1200.000 ;
    END
  END cpu_dtr_n1[12]
  PIN cpu_dtr_n1[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.470 1196.000 990.750 1200.000 ;
    END
  END cpu_dtr_n1[13]
  PIN cpu_dtr_n1[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.510 1196.000 1001.790 1200.000 ;
    END
  END cpu_dtr_n1[14]
  PIN cpu_dtr_n1[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.010 1196.000 1013.290 1200.000 ;
    END
  END cpu_dtr_n1[15]
  PIN cpu_dtr_n1[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1024.510 1196.000 1024.790 1200.000 ;
    END
  END cpu_dtr_n1[16]
  PIN cpu_dtr_n1[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.550 1196.000 1035.830 1200.000 ;
    END
  END cpu_dtr_n1[17]
  PIN cpu_dtr_n1[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1047.050 1196.000 1047.330 1200.000 ;
    END
  END cpu_dtr_n1[18]
  PIN cpu_dtr_n1[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.550 1196.000 1058.830 1200.000 ;
    END
  END cpu_dtr_n1[19]
  PIN cpu_dtr_n1[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.310 1196.000 854.590 1200.000 ;
    END
  END cpu_dtr_n1[1]
  PIN cpu_dtr_n1[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.590 1196.000 1069.870 1200.000 ;
    END
  END cpu_dtr_n1[20]
  PIN cpu_dtr_n1[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.090 1196.000 1081.370 1200.000 ;
    END
  END cpu_dtr_n1[21]
  PIN cpu_dtr_n1[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.130 1196.000 1092.410 1200.000 ;
    END
  END cpu_dtr_n1[22]
  PIN cpu_dtr_n1[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1103.630 1196.000 1103.910 1200.000 ;
    END
  END cpu_dtr_n1[23]
  PIN cpu_dtr_n1[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1115.130 1196.000 1115.410 1200.000 ;
    END
  END cpu_dtr_n1[24]
  PIN cpu_dtr_n1[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.170 1196.000 1126.450 1200.000 ;
    END
  END cpu_dtr_n1[25]
  PIN cpu_dtr_n1[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1137.670 1196.000 1137.950 1200.000 ;
    END
  END cpu_dtr_n1[26]
  PIN cpu_dtr_n1[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1148.710 1196.000 1148.990 1200.000 ;
    END
  END cpu_dtr_n1[27]
  PIN cpu_dtr_n1[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.210 1196.000 1160.490 1200.000 ;
    END
  END cpu_dtr_n1[28]
  PIN cpu_dtr_n1[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1171.710 1196.000 1171.990 1200.000 ;
    END
  END cpu_dtr_n1[29]
  PIN cpu_dtr_n1[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 865.810 1196.000 866.090 1200.000 ;
    END
  END cpu_dtr_n1[2]
  PIN cpu_dtr_n1[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1182.750 1196.000 1183.030 1200.000 ;
    END
  END cpu_dtr_n1[30]
  PIN cpu_dtr_n1[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.250 1196.000 1194.530 1200.000 ;
    END
  END cpu_dtr_n1[31]
  PIN cpu_dtr_n1[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 877.310 1196.000 877.590 1200.000 ;
    END
  END cpu_dtr_n1[3]
  PIN cpu_dtr_n1[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.350 1196.000 888.630 1200.000 ;
    END
  END cpu_dtr_n1[4]
  PIN cpu_dtr_n1[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 899.850 1196.000 900.130 1200.000 ;
    END
  END cpu_dtr_n1[5]
  PIN cpu_dtr_n1[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.350 1196.000 911.630 1200.000 ;
    END
  END cpu_dtr_n1[6]
  PIN cpu_dtr_n1[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.390 1196.000 922.670 1200.000 ;
    END
  END cpu_dtr_n1[7]
  PIN cpu_dtr_n1[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 933.890 1196.000 934.170 1200.000 ;
    END
  END cpu_dtr_n1[8]
  PIN cpu_dtr_n1[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.930 1196.000 945.210 1200.000 ;
    END
  END cpu_dtr_n1[9]
  PIN cpu_dtw_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 665.760 1200.000 666.360 ;
    END
  END cpu_dtw_e[0]
  PIN cpu_dtw_e[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 775.920 1200.000 776.520 ;
    END
  END cpu_dtw_e[10]
  PIN cpu_dtw_e[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 786.800 1200.000 787.400 ;
    END
  END cpu_dtw_e[11]
  PIN cpu_dtw_e[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 797.680 1200.000 798.280 ;
    END
  END cpu_dtw_e[12]
  PIN cpu_dtw_e[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 809.240 1200.000 809.840 ;
    END
  END cpu_dtw_e[13]
  PIN cpu_dtw_e[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 820.120 1200.000 820.720 ;
    END
  END cpu_dtw_e[14]
  PIN cpu_dtw_e[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 831.000 1200.000 831.600 ;
    END
  END cpu_dtw_e[15]
  PIN cpu_dtw_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 676.640 1200.000 677.240 ;
    END
  END cpu_dtw_e[1]
  PIN cpu_dtw_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 687.520 1200.000 688.120 ;
    END
  END cpu_dtw_e[2]
  PIN cpu_dtw_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 699.080 1200.000 699.680 ;
    END
  END cpu_dtw_e[3]
  PIN cpu_dtw_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 709.960 1200.000 710.560 ;
    END
  END cpu_dtw_e[4]
  PIN cpu_dtw_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 720.840 1200.000 721.440 ;
    END
  END cpu_dtw_e[5]
  PIN cpu_dtw_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 731.720 1200.000 732.320 ;
    END
  END cpu_dtw_e[6]
  PIN cpu_dtw_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 742.600 1200.000 743.200 ;
    END
  END cpu_dtw_e[7]
  PIN cpu_dtw_e[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 754.160 1200.000 754.760 ;
    END
  END cpu_dtw_e[8]
  PIN cpu_dtw_e[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 765.040 1200.000 765.640 ;
    END
  END cpu_dtw_e[9]
  PIN cpu_dtw_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 662.030 1196.000 662.310 1200.000 ;
    END
  END cpu_dtw_n[0]
  PIN cpu_dtw_n[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.190 1196.000 775.470 1200.000 ;
    END
  END cpu_dtw_n[10]
  PIN cpu_dtw_n[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.690 1196.000 786.970 1200.000 ;
    END
  END cpu_dtw_n[11]
  PIN cpu_dtw_n[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.730 1196.000 798.010 1200.000 ;
    END
  END cpu_dtw_n[12]
  PIN cpu_dtw_n[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 809.230 1196.000 809.510 1200.000 ;
    END
  END cpu_dtw_n[13]
  PIN cpu_dtw_n[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 820.730 1196.000 821.010 1200.000 ;
    END
  END cpu_dtw_n[14]
  PIN cpu_dtw_n[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 831.770 1196.000 832.050 1200.000 ;
    END
  END cpu_dtw_n[15]
  PIN cpu_dtw_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.530 1196.000 673.810 1200.000 ;
    END
  END cpu_dtw_n[1]
  PIN cpu_dtw_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 684.570 1196.000 684.850 1200.000 ;
    END
  END cpu_dtw_n[2]
  PIN cpu_dtw_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.070 1196.000 696.350 1200.000 ;
    END
  END cpu_dtw_n[3]
  PIN cpu_dtw_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.570 1196.000 707.850 1200.000 ;
    END
  END cpu_dtw_n[4]
  PIN cpu_dtw_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.610 1196.000 718.890 1200.000 ;
    END
  END cpu_dtw_n[5]
  PIN cpu_dtw_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 730.110 1196.000 730.390 1200.000 ;
    END
  END cpu_dtw_n[6]
  PIN cpu_dtw_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.150 1196.000 741.430 1200.000 ;
    END
  END cpu_dtw_n[7]
  PIN cpu_dtw_n[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 752.650 1196.000 752.930 1200.000 ;
    END
  END cpu_dtw_n[8]
  PIN cpu_dtw_n[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 764.150 1196.000 764.430 1200.000 ;
    END
  END cpu_dtw_n[9]
  PIN cpu_mask_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 379.480 1200.000 380.080 ;
    END
  END cpu_mask_e[0]
  PIN cpu_mask_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 390.360 1200.000 390.960 ;
    END
  END cpu_mask_e[1]
  PIN cpu_mask_e[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 401.240 1200.000 401.840 ;
    END
  END cpu_mask_e[2]
  PIN cpu_mask_e[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 412.800 1200.000 413.400 ;
    END
  END cpu_mask_e[3]
  PIN cpu_mask_e[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 423.680 1200.000 424.280 ;
    END
  END cpu_mask_e[4]
  PIN cpu_mask_e[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 434.560 1200.000 435.160 ;
    END
  END cpu_mask_e[5]
  PIN cpu_mask_e[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 445.440 1200.000 446.040 ;
    END
  END cpu_mask_e[6]
  PIN cpu_mask_e[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 456.320 1200.000 456.920 ;
    END
  END cpu_mask_e[7]
  PIN cpu_mask_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 548.870 1196.000 549.150 1200.000 ;
    END
  END cpu_mask_n[0]
  PIN cpu_mask_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 560.370 1196.000 560.650 1200.000 ;
    END
  END cpu_mask_n[1]
  PIN cpu_mask_n[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.410 1196.000 571.690 1200.000 ;
    END
  END cpu_mask_n[2]
  PIN cpu_mask_n[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.910 1196.000 583.190 1200.000 ;
    END
  END cpu_mask_n[3]
  PIN cpu_mask_n[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.950 1196.000 594.230 1200.000 ;
    END
  END cpu_mask_n[4]
  PIN cpu_mask_n[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 605.450 1196.000 605.730 1200.000 ;
    END
  END cpu_mask_n[5]
  PIN cpu_mask_n[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.950 1196.000 617.230 1200.000 ;
    END
  END cpu_mask_n[6]
  PIN cpu_mask_n[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 627.990 1196.000 628.270 1200.000 ;
    END
  END cpu_mask_n[7]
  PIN cpu_wen_e[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 467.880 1200.000 468.480 ;
    END
  END cpu_wen_e[0]
  PIN cpu_wen_e[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 478.760 1200.000 479.360 ;
    END
  END cpu_wen_e[1]
  PIN cpu_wen_n[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 639.490 1196.000 639.770 1200.000 ;
    END
  END cpu_wen_n[0]
  PIN cpu_wen_n[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.530 1196.000 650.810 1200.000 ;
    END
  END cpu_wen_n[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 351.600 4.000 352.200 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 383.560 4.000 384.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.280 4.000 573.880 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 762.320 4.000 762.920 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 857.520 4.000 858.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 888.800 4.000 889.400 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 920.080 4.000 920.680 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.360 4.000 67.960 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 952.040 4.000 952.640 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 983.320 4.000 983.920 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1015.280 4.000 1015.880 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1046.560 4.000 1047.160 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1078.520 4.000 1079.120 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.800 4.000 1110.400 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1141.760 4.000 1142.360 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1173.040 4.000 1173.640 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 99.320 4.000 99.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 130.600 4.000 131.200 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.000 4.000 15.600 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.520 4.000 331.120 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 362.480 4.000 363.080 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.720 4.000 426.320 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.760 4.000 615.360 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.720 4.000 647.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 709.960 4.000 710.560 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 804.480 4.000 805.080 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 867.720 4.000 868.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 899.680 4.000 900.280 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 930.960 4.000 931.560 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 962.240 4.000 962.840 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 994.200 4.000 994.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1025.480 4.000 1026.080 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1057.440 4.000 1058.040 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1088.720 4.000 1089.320 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1120.680 4.000 1121.280 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.960 4.000 1152.560 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1183.920 4.000 1184.520 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 109.520 4.000 110.120 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.000 4.000 236.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.960 4.000 268.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 4.000 499.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.120 4.000 531.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 594.360 4.000 594.960 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 625.640 4.000 626.240 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.920 4.000 657.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.880 4.000 689.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.160 4.000 720.760 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 752.120 4.000 752.720 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 815.360 4.000 815.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 4.000 847.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 878.600 4.000 879.200 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 909.880 4.000 910.480 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 973.120 4.000 973.720 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1004.400 4.000 1005.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1036.360 4.000 1036.960 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1067.640 4.000 1068.240 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1099.600 4.000 1100.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1130.880 4.000 1131.480 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1162.840 4.000 1163.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.120 4.000 1194.720 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.160 4.000 278.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1141.350 0.000 1141.630 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.090 0.000 1173.370 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1194.250 0.000 1194.530 4.000 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1151.930 0.000 1152.210 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1183.670 0.000 1183.950 4.000 ;
    END
  END la_oen[1]
  PIN one
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 16.360 1200.000 16.960 ;
    END
  END one
  PIN ram_ce
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 1194.120 1200.000 1194.720 ;
    END
  END ram_ce
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.730 0.000 16.010 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 493.670 0.000 493.950 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.930 0.000 876.210 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.350 0.000 1003.630 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.090 0.000 1035.370 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 153.730 0.000 154.010 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1066.830 0.000 1067.110 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1099.030 0.000 1099.310 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.310 0.000 440.590 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.250 0.000 504.530 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.990 0.000 536.270 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.350 0.000 727.630 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 790.830 0.000 791.110 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.770 0.000 855.050 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.510 0.000 886.790 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.250 0.000 918.530 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.990 0.000 950.270 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 982.190 0.000 982.470 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.930 0.000 1014.210 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.670 0.000 1045.950 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.410 0.000 1077.690 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.630 0.000 206.910 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 546.570 0.000 546.850 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 642.250 0.000 642.530 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 833.150 0.000 833.430 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 897.090 0.000 897.370 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 928.830 0.000 929.110 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.570 0.000 960.850 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.770 0.000 993.050 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.510 0.000 1024.790 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1056.250 0.000 1056.530 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.450 0.000 1088.730 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.190 0.000 1120.470 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 387.410 0.000 387.690 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.470 0.000 47.750 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END wbs_we_i
  PIN zero
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1196.000 5.480 1200.000 6.080 ;
    END
  END zero
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1188.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1188.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1194.160 1188.725 ;
      LAYER met1 ;
        RECT 5.130 4.460 1194.550 1189.280 ;
      LAYER met2 ;
        RECT 5.160 1195.720 5.330 1196.000 ;
        RECT 6.170 1195.720 16.370 1196.000 ;
        RECT 17.210 1195.720 27.870 1196.000 ;
        RECT 28.710 1195.720 38.910 1196.000 ;
        RECT 39.750 1195.720 50.410 1196.000 ;
        RECT 51.250 1195.720 61.910 1196.000 ;
        RECT 62.750 1195.720 72.950 1196.000 ;
        RECT 73.790 1195.720 84.450 1196.000 ;
        RECT 85.290 1195.720 95.490 1196.000 ;
        RECT 96.330 1195.720 106.990 1196.000 ;
        RECT 107.830 1195.720 118.490 1196.000 ;
        RECT 119.330 1195.720 129.530 1196.000 ;
        RECT 130.370 1195.720 141.030 1196.000 ;
        RECT 141.870 1195.720 152.070 1196.000 ;
        RECT 152.910 1195.720 163.570 1196.000 ;
        RECT 164.410 1195.720 175.070 1196.000 ;
        RECT 175.910 1195.720 186.110 1196.000 ;
        RECT 186.950 1195.720 197.610 1196.000 ;
        RECT 198.450 1195.720 209.110 1196.000 ;
        RECT 209.950 1195.720 220.150 1196.000 ;
        RECT 220.990 1195.720 231.650 1196.000 ;
        RECT 232.490 1195.720 242.690 1196.000 ;
        RECT 243.530 1195.720 254.190 1196.000 ;
        RECT 255.030 1195.720 265.690 1196.000 ;
        RECT 266.530 1195.720 276.730 1196.000 ;
        RECT 277.570 1195.720 288.230 1196.000 ;
        RECT 289.070 1195.720 299.270 1196.000 ;
        RECT 300.110 1195.720 310.770 1196.000 ;
        RECT 311.610 1195.720 322.270 1196.000 ;
        RECT 323.110 1195.720 333.310 1196.000 ;
        RECT 334.150 1195.720 344.810 1196.000 ;
        RECT 345.650 1195.720 356.310 1196.000 ;
        RECT 357.150 1195.720 367.350 1196.000 ;
        RECT 368.190 1195.720 378.850 1196.000 ;
        RECT 379.690 1195.720 389.890 1196.000 ;
        RECT 390.730 1195.720 401.390 1196.000 ;
        RECT 402.230 1195.720 412.890 1196.000 ;
        RECT 413.730 1195.720 423.930 1196.000 ;
        RECT 424.770 1195.720 435.430 1196.000 ;
        RECT 436.270 1195.720 446.470 1196.000 ;
        RECT 447.310 1195.720 457.970 1196.000 ;
        RECT 458.810 1195.720 469.470 1196.000 ;
        RECT 470.310 1195.720 480.510 1196.000 ;
        RECT 481.350 1195.720 492.010 1196.000 ;
        RECT 492.850 1195.720 503.050 1196.000 ;
        RECT 503.890 1195.720 514.550 1196.000 ;
        RECT 515.390 1195.720 526.050 1196.000 ;
        RECT 526.890 1195.720 537.090 1196.000 ;
        RECT 537.930 1195.720 548.590 1196.000 ;
        RECT 549.430 1195.720 560.090 1196.000 ;
        RECT 560.930 1195.720 571.130 1196.000 ;
        RECT 571.970 1195.720 582.630 1196.000 ;
        RECT 583.470 1195.720 593.670 1196.000 ;
        RECT 594.510 1195.720 605.170 1196.000 ;
        RECT 606.010 1195.720 616.670 1196.000 ;
        RECT 617.510 1195.720 627.710 1196.000 ;
        RECT 628.550 1195.720 639.210 1196.000 ;
        RECT 640.050 1195.720 650.250 1196.000 ;
        RECT 651.090 1195.720 661.750 1196.000 ;
        RECT 662.590 1195.720 673.250 1196.000 ;
        RECT 674.090 1195.720 684.290 1196.000 ;
        RECT 685.130 1195.720 695.790 1196.000 ;
        RECT 696.630 1195.720 707.290 1196.000 ;
        RECT 708.130 1195.720 718.330 1196.000 ;
        RECT 719.170 1195.720 729.830 1196.000 ;
        RECT 730.670 1195.720 740.870 1196.000 ;
        RECT 741.710 1195.720 752.370 1196.000 ;
        RECT 753.210 1195.720 763.870 1196.000 ;
        RECT 764.710 1195.720 774.910 1196.000 ;
        RECT 775.750 1195.720 786.410 1196.000 ;
        RECT 787.250 1195.720 797.450 1196.000 ;
        RECT 798.290 1195.720 808.950 1196.000 ;
        RECT 809.790 1195.720 820.450 1196.000 ;
        RECT 821.290 1195.720 831.490 1196.000 ;
        RECT 832.330 1195.720 842.990 1196.000 ;
        RECT 843.830 1195.720 854.030 1196.000 ;
        RECT 854.870 1195.720 865.530 1196.000 ;
        RECT 866.370 1195.720 877.030 1196.000 ;
        RECT 877.870 1195.720 888.070 1196.000 ;
        RECT 888.910 1195.720 899.570 1196.000 ;
        RECT 900.410 1195.720 911.070 1196.000 ;
        RECT 911.910 1195.720 922.110 1196.000 ;
        RECT 922.950 1195.720 933.610 1196.000 ;
        RECT 934.450 1195.720 944.650 1196.000 ;
        RECT 945.490 1195.720 956.150 1196.000 ;
        RECT 956.990 1195.720 967.650 1196.000 ;
        RECT 968.490 1195.720 978.690 1196.000 ;
        RECT 979.530 1195.720 990.190 1196.000 ;
        RECT 991.030 1195.720 1001.230 1196.000 ;
        RECT 1002.070 1195.720 1012.730 1196.000 ;
        RECT 1013.570 1195.720 1024.230 1196.000 ;
        RECT 1025.070 1195.720 1035.270 1196.000 ;
        RECT 1036.110 1195.720 1046.770 1196.000 ;
        RECT 1047.610 1195.720 1058.270 1196.000 ;
        RECT 1059.110 1195.720 1069.310 1196.000 ;
        RECT 1070.150 1195.720 1080.810 1196.000 ;
        RECT 1081.650 1195.720 1091.850 1196.000 ;
        RECT 1092.690 1195.720 1103.350 1196.000 ;
        RECT 1104.190 1195.720 1114.850 1196.000 ;
        RECT 1115.690 1195.720 1125.890 1196.000 ;
        RECT 1126.730 1195.720 1137.390 1196.000 ;
        RECT 1138.230 1195.720 1148.430 1196.000 ;
        RECT 1149.270 1195.720 1159.930 1196.000 ;
        RECT 1160.770 1195.720 1171.430 1196.000 ;
        RECT 1172.270 1195.720 1182.470 1196.000 ;
        RECT 1183.310 1195.720 1193.970 1196.000 ;
        RECT 5.160 4.280 1194.520 1195.720 ;
        RECT 5.710 4.000 15.450 4.280 ;
        RECT 16.290 4.000 26.030 4.280 ;
        RECT 26.870 4.000 36.610 4.280 ;
        RECT 37.450 4.000 47.190 4.280 ;
        RECT 48.030 4.000 57.770 4.280 ;
        RECT 58.610 4.000 68.350 4.280 ;
        RECT 69.190 4.000 78.930 4.280 ;
        RECT 79.770 4.000 89.510 4.280 ;
        RECT 90.350 4.000 100.090 4.280 ;
        RECT 100.930 4.000 110.670 4.280 ;
        RECT 111.510 4.000 121.250 4.280 ;
        RECT 122.090 4.000 132.290 4.280 ;
        RECT 133.130 4.000 142.870 4.280 ;
        RECT 143.710 4.000 153.450 4.280 ;
        RECT 154.290 4.000 164.030 4.280 ;
        RECT 164.870 4.000 174.610 4.280 ;
        RECT 175.450 4.000 185.190 4.280 ;
        RECT 186.030 4.000 195.770 4.280 ;
        RECT 196.610 4.000 206.350 4.280 ;
        RECT 207.190 4.000 216.930 4.280 ;
        RECT 217.770 4.000 227.510 4.280 ;
        RECT 228.350 4.000 238.090 4.280 ;
        RECT 238.930 4.000 249.130 4.280 ;
        RECT 249.970 4.000 259.710 4.280 ;
        RECT 260.550 4.000 270.290 4.280 ;
        RECT 271.130 4.000 280.870 4.280 ;
        RECT 281.710 4.000 291.450 4.280 ;
        RECT 292.290 4.000 302.030 4.280 ;
        RECT 302.870 4.000 312.610 4.280 ;
        RECT 313.450 4.000 323.190 4.280 ;
        RECT 324.030 4.000 333.770 4.280 ;
        RECT 334.610 4.000 344.350 4.280 ;
        RECT 345.190 4.000 354.930 4.280 ;
        RECT 355.770 4.000 365.970 4.280 ;
        RECT 366.810 4.000 376.550 4.280 ;
        RECT 377.390 4.000 387.130 4.280 ;
        RECT 387.970 4.000 397.710 4.280 ;
        RECT 398.550 4.000 408.290 4.280 ;
        RECT 409.130 4.000 418.870 4.280 ;
        RECT 419.710 4.000 429.450 4.280 ;
        RECT 430.290 4.000 440.030 4.280 ;
        RECT 440.870 4.000 450.610 4.280 ;
        RECT 451.450 4.000 461.190 4.280 ;
        RECT 462.030 4.000 471.770 4.280 ;
        RECT 472.610 4.000 482.350 4.280 ;
        RECT 483.190 4.000 493.390 4.280 ;
        RECT 494.230 4.000 503.970 4.280 ;
        RECT 504.810 4.000 514.550 4.280 ;
        RECT 515.390 4.000 525.130 4.280 ;
        RECT 525.970 4.000 535.710 4.280 ;
        RECT 536.550 4.000 546.290 4.280 ;
        RECT 547.130 4.000 556.870 4.280 ;
        RECT 557.710 4.000 567.450 4.280 ;
        RECT 568.290 4.000 578.030 4.280 ;
        RECT 578.870 4.000 588.610 4.280 ;
        RECT 589.450 4.000 599.190 4.280 ;
        RECT 600.030 4.000 610.230 4.280 ;
        RECT 611.070 4.000 620.810 4.280 ;
        RECT 621.650 4.000 631.390 4.280 ;
        RECT 632.230 4.000 641.970 4.280 ;
        RECT 642.810 4.000 652.550 4.280 ;
        RECT 653.390 4.000 663.130 4.280 ;
        RECT 663.970 4.000 673.710 4.280 ;
        RECT 674.550 4.000 684.290 4.280 ;
        RECT 685.130 4.000 694.870 4.280 ;
        RECT 695.710 4.000 705.450 4.280 ;
        RECT 706.290 4.000 716.030 4.280 ;
        RECT 716.870 4.000 727.070 4.280 ;
        RECT 727.910 4.000 737.650 4.280 ;
        RECT 738.490 4.000 748.230 4.280 ;
        RECT 749.070 4.000 758.810 4.280 ;
        RECT 759.650 4.000 769.390 4.280 ;
        RECT 770.230 4.000 779.970 4.280 ;
        RECT 780.810 4.000 790.550 4.280 ;
        RECT 791.390 4.000 801.130 4.280 ;
        RECT 801.970 4.000 811.710 4.280 ;
        RECT 812.550 4.000 822.290 4.280 ;
        RECT 823.130 4.000 832.870 4.280 ;
        RECT 833.710 4.000 843.450 4.280 ;
        RECT 844.290 4.000 854.490 4.280 ;
        RECT 855.330 4.000 865.070 4.280 ;
        RECT 865.910 4.000 875.650 4.280 ;
        RECT 876.490 4.000 886.230 4.280 ;
        RECT 887.070 4.000 896.810 4.280 ;
        RECT 897.650 4.000 907.390 4.280 ;
        RECT 908.230 4.000 917.970 4.280 ;
        RECT 918.810 4.000 928.550 4.280 ;
        RECT 929.390 4.000 939.130 4.280 ;
        RECT 939.970 4.000 949.710 4.280 ;
        RECT 950.550 4.000 960.290 4.280 ;
        RECT 961.130 4.000 971.330 4.280 ;
        RECT 972.170 4.000 981.910 4.280 ;
        RECT 982.750 4.000 992.490 4.280 ;
        RECT 993.330 4.000 1003.070 4.280 ;
        RECT 1003.910 4.000 1013.650 4.280 ;
        RECT 1014.490 4.000 1024.230 4.280 ;
        RECT 1025.070 4.000 1034.810 4.280 ;
        RECT 1035.650 4.000 1045.390 4.280 ;
        RECT 1046.230 4.000 1055.970 4.280 ;
        RECT 1056.810 4.000 1066.550 4.280 ;
        RECT 1067.390 4.000 1077.130 4.280 ;
        RECT 1077.970 4.000 1088.170 4.280 ;
        RECT 1089.010 4.000 1098.750 4.280 ;
        RECT 1099.590 4.000 1109.330 4.280 ;
        RECT 1110.170 4.000 1119.910 4.280 ;
        RECT 1120.750 4.000 1130.490 4.280 ;
        RECT 1131.330 4.000 1141.070 4.280 ;
        RECT 1141.910 4.000 1151.650 4.280 ;
        RECT 1152.490 4.000 1162.230 4.280 ;
        RECT 1163.070 4.000 1172.810 4.280 ;
        RECT 1173.650 4.000 1183.390 4.280 ;
        RECT 1184.230 4.000 1193.970 4.280 ;
      LAYER met3 ;
        RECT 4.400 1193.720 1195.600 1194.585 ;
        RECT 4.000 1184.920 1196.000 1193.720 ;
        RECT 4.400 1184.240 1196.000 1184.920 ;
        RECT 4.400 1183.520 1195.600 1184.240 ;
        RECT 4.000 1182.840 1195.600 1183.520 ;
        RECT 4.000 1174.040 1196.000 1182.840 ;
        RECT 4.400 1173.360 1196.000 1174.040 ;
        RECT 4.400 1172.640 1195.600 1173.360 ;
        RECT 4.000 1171.960 1195.600 1172.640 ;
        RECT 4.000 1163.840 1196.000 1171.960 ;
        RECT 4.400 1162.480 1196.000 1163.840 ;
        RECT 4.400 1162.440 1195.600 1162.480 ;
        RECT 4.000 1161.080 1195.600 1162.440 ;
        RECT 4.000 1152.960 1196.000 1161.080 ;
        RECT 4.400 1151.600 1196.000 1152.960 ;
        RECT 4.400 1151.560 1195.600 1151.600 ;
        RECT 4.000 1150.200 1195.600 1151.560 ;
        RECT 4.000 1142.760 1196.000 1150.200 ;
        RECT 4.400 1141.360 1196.000 1142.760 ;
        RECT 4.000 1140.040 1196.000 1141.360 ;
        RECT 4.000 1138.640 1195.600 1140.040 ;
        RECT 4.000 1131.880 1196.000 1138.640 ;
        RECT 4.400 1130.480 1196.000 1131.880 ;
        RECT 4.000 1129.160 1196.000 1130.480 ;
        RECT 4.000 1127.760 1195.600 1129.160 ;
        RECT 4.000 1121.680 1196.000 1127.760 ;
        RECT 4.400 1120.280 1196.000 1121.680 ;
        RECT 4.000 1118.280 1196.000 1120.280 ;
        RECT 4.000 1116.880 1195.600 1118.280 ;
        RECT 4.000 1110.800 1196.000 1116.880 ;
        RECT 4.400 1109.400 1196.000 1110.800 ;
        RECT 4.000 1107.400 1196.000 1109.400 ;
        RECT 4.000 1106.000 1195.600 1107.400 ;
        RECT 4.000 1100.600 1196.000 1106.000 ;
        RECT 4.400 1099.200 1196.000 1100.600 ;
        RECT 4.000 1096.520 1196.000 1099.200 ;
        RECT 4.000 1095.120 1195.600 1096.520 ;
        RECT 4.000 1089.720 1196.000 1095.120 ;
        RECT 4.400 1088.320 1196.000 1089.720 ;
        RECT 4.000 1084.960 1196.000 1088.320 ;
        RECT 4.000 1083.560 1195.600 1084.960 ;
        RECT 4.000 1079.520 1196.000 1083.560 ;
        RECT 4.400 1078.120 1196.000 1079.520 ;
        RECT 4.000 1074.080 1196.000 1078.120 ;
        RECT 4.000 1072.680 1195.600 1074.080 ;
        RECT 4.000 1068.640 1196.000 1072.680 ;
        RECT 4.400 1067.240 1196.000 1068.640 ;
        RECT 4.000 1063.200 1196.000 1067.240 ;
        RECT 4.000 1061.800 1195.600 1063.200 ;
        RECT 4.000 1058.440 1196.000 1061.800 ;
        RECT 4.400 1057.040 1196.000 1058.440 ;
        RECT 4.000 1052.320 1196.000 1057.040 ;
        RECT 4.000 1050.920 1195.600 1052.320 ;
        RECT 4.000 1047.560 1196.000 1050.920 ;
        RECT 4.400 1046.160 1196.000 1047.560 ;
        RECT 4.000 1041.440 1196.000 1046.160 ;
        RECT 4.000 1040.040 1195.600 1041.440 ;
        RECT 4.000 1037.360 1196.000 1040.040 ;
        RECT 4.400 1035.960 1196.000 1037.360 ;
        RECT 4.000 1029.880 1196.000 1035.960 ;
        RECT 4.000 1028.480 1195.600 1029.880 ;
        RECT 4.000 1026.480 1196.000 1028.480 ;
        RECT 4.400 1025.080 1196.000 1026.480 ;
        RECT 4.000 1019.000 1196.000 1025.080 ;
        RECT 4.000 1017.600 1195.600 1019.000 ;
        RECT 4.000 1016.280 1196.000 1017.600 ;
        RECT 4.400 1014.880 1196.000 1016.280 ;
        RECT 4.000 1008.120 1196.000 1014.880 ;
        RECT 4.000 1006.720 1195.600 1008.120 ;
        RECT 4.000 1005.400 1196.000 1006.720 ;
        RECT 4.400 1004.000 1196.000 1005.400 ;
        RECT 4.000 997.240 1196.000 1004.000 ;
        RECT 4.000 995.840 1195.600 997.240 ;
        RECT 4.000 995.200 1196.000 995.840 ;
        RECT 4.400 993.800 1196.000 995.200 ;
        RECT 4.000 986.360 1196.000 993.800 ;
        RECT 4.000 984.960 1195.600 986.360 ;
        RECT 4.000 984.320 1196.000 984.960 ;
        RECT 4.400 982.920 1196.000 984.320 ;
        RECT 4.000 974.800 1196.000 982.920 ;
        RECT 4.000 974.120 1195.600 974.800 ;
        RECT 4.400 973.400 1195.600 974.120 ;
        RECT 4.400 972.720 1196.000 973.400 ;
        RECT 4.000 963.920 1196.000 972.720 ;
        RECT 4.000 963.240 1195.600 963.920 ;
        RECT 4.400 962.520 1195.600 963.240 ;
        RECT 4.400 961.840 1196.000 962.520 ;
        RECT 4.000 953.040 1196.000 961.840 ;
        RECT 4.400 951.640 1195.600 953.040 ;
        RECT 4.000 942.160 1196.000 951.640 ;
        RECT 4.400 940.760 1195.600 942.160 ;
        RECT 4.000 931.960 1196.000 940.760 ;
        RECT 4.400 931.280 1196.000 931.960 ;
        RECT 4.400 930.560 1195.600 931.280 ;
        RECT 4.000 929.880 1195.600 930.560 ;
        RECT 4.000 921.080 1196.000 929.880 ;
        RECT 4.400 919.720 1196.000 921.080 ;
        RECT 4.400 919.680 1195.600 919.720 ;
        RECT 4.000 918.320 1195.600 919.680 ;
        RECT 4.000 910.880 1196.000 918.320 ;
        RECT 4.400 909.480 1196.000 910.880 ;
        RECT 4.000 908.840 1196.000 909.480 ;
        RECT 4.000 907.440 1195.600 908.840 ;
        RECT 4.000 900.680 1196.000 907.440 ;
        RECT 4.400 899.280 1196.000 900.680 ;
        RECT 4.000 897.960 1196.000 899.280 ;
        RECT 4.000 896.560 1195.600 897.960 ;
        RECT 4.000 889.800 1196.000 896.560 ;
        RECT 4.400 888.400 1196.000 889.800 ;
        RECT 4.000 887.080 1196.000 888.400 ;
        RECT 4.000 885.680 1195.600 887.080 ;
        RECT 4.000 879.600 1196.000 885.680 ;
        RECT 4.400 878.200 1196.000 879.600 ;
        RECT 4.000 876.200 1196.000 878.200 ;
        RECT 4.000 874.800 1195.600 876.200 ;
        RECT 4.000 868.720 1196.000 874.800 ;
        RECT 4.400 867.320 1196.000 868.720 ;
        RECT 4.000 865.320 1196.000 867.320 ;
        RECT 4.000 863.920 1195.600 865.320 ;
        RECT 4.000 858.520 1196.000 863.920 ;
        RECT 4.400 857.120 1196.000 858.520 ;
        RECT 4.000 853.760 1196.000 857.120 ;
        RECT 4.000 852.360 1195.600 853.760 ;
        RECT 4.000 847.640 1196.000 852.360 ;
        RECT 4.400 846.240 1196.000 847.640 ;
        RECT 4.000 842.880 1196.000 846.240 ;
        RECT 4.000 841.480 1195.600 842.880 ;
        RECT 4.000 837.440 1196.000 841.480 ;
        RECT 4.400 836.040 1196.000 837.440 ;
        RECT 4.000 832.000 1196.000 836.040 ;
        RECT 4.000 830.600 1195.600 832.000 ;
        RECT 4.000 826.560 1196.000 830.600 ;
        RECT 4.400 825.160 1196.000 826.560 ;
        RECT 4.000 821.120 1196.000 825.160 ;
        RECT 4.000 819.720 1195.600 821.120 ;
        RECT 4.000 816.360 1196.000 819.720 ;
        RECT 4.400 814.960 1196.000 816.360 ;
        RECT 4.000 810.240 1196.000 814.960 ;
        RECT 4.000 808.840 1195.600 810.240 ;
        RECT 4.000 805.480 1196.000 808.840 ;
        RECT 4.400 804.080 1196.000 805.480 ;
        RECT 4.000 798.680 1196.000 804.080 ;
        RECT 4.000 797.280 1195.600 798.680 ;
        RECT 4.000 795.280 1196.000 797.280 ;
        RECT 4.400 793.880 1196.000 795.280 ;
        RECT 4.000 787.800 1196.000 793.880 ;
        RECT 4.000 786.400 1195.600 787.800 ;
        RECT 4.000 784.400 1196.000 786.400 ;
        RECT 4.400 783.000 1196.000 784.400 ;
        RECT 4.000 776.920 1196.000 783.000 ;
        RECT 4.000 775.520 1195.600 776.920 ;
        RECT 4.000 774.200 1196.000 775.520 ;
        RECT 4.400 772.800 1196.000 774.200 ;
        RECT 4.000 766.040 1196.000 772.800 ;
        RECT 4.000 764.640 1195.600 766.040 ;
        RECT 4.000 763.320 1196.000 764.640 ;
        RECT 4.400 761.920 1196.000 763.320 ;
        RECT 4.000 755.160 1196.000 761.920 ;
        RECT 4.000 753.760 1195.600 755.160 ;
        RECT 4.000 753.120 1196.000 753.760 ;
        RECT 4.400 751.720 1196.000 753.120 ;
        RECT 4.000 743.600 1196.000 751.720 ;
        RECT 4.000 742.240 1195.600 743.600 ;
        RECT 4.400 742.200 1195.600 742.240 ;
        RECT 4.400 740.840 1196.000 742.200 ;
        RECT 4.000 732.720 1196.000 740.840 ;
        RECT 4.000 732.040 1195.600 732.720 ;
        RECT 4.400 731.320 1195.600 732.040 ;
        RECT 4.400 730.640 1196.000 731.320 ;
        RECT 4.000 721.840 1196.000 730.640 ;
        RECT 4.000 721.160 1195.600 721.840 ;
        RECT 4.400 720.440 1195.600 721.160 ;
        RECT 4.400 719.760 1196.000 720.440 ;
        RECT 4.000 710.960 1196.000 719.760 ;
        RECT 4.400 709.560 1195.600 710.960 ;
        RECT 4.000 700.080 1196.000 709.560 ;
        RECT 4.400 698.680 1195.600 700.080 ;
        RECT 4.000 689.880 1196.000 698.680 ;
        RECT 4.400 688.520 1196.000 689.880 ;
        RECT 4.400 688.480 1195.600 688.520 ;
        RECT 4.000 687.120 1195.600 688.480 ;
        RECT 4.000 679.000 1196.000 687.120 ;
        RECT 4.400 677.640 1196.000 679.000 ;
        RECT 4.400 677.600 1195.600 677.640 ;
        RECT 4.000 676.240 1195.600 677.600 ;
        RECT 4.000 668.800 1196.000 676.240 ;
        RECT 4.400 667.400 1196.000 668.800 ;
        RECT 4.000 666.760 1196.000 667.400 ;
        RECT 4.000 665.360 1195.600 666.760 ;
        RECT 4.000 657.920 1196.000 665.360 ;
        RECT 4.400 656.520 1196.000 657.920 ;
        RECT 4.000 655.880 1196.000 656.520 ;
        RECT 4.000 654.480 1195.600 655.880 ;
        RECT 4.000 647.720 1196.000 654.480 ;
        RECT 4.400 646.320 1196.000 647.720 ;
        RECT 4.000 645.000 1196.000 646.320 ;
        RECT 4.000 643.600 1195.600 645.000 ;
        RECT 4.000 636.840 1196.000 643.600 ;
        RECT 4.400 635.440 1196.000 636.840 ;
        RECT 4.000 633.440 1196.000 635.440 ;
        RECT 4.000 632.040 1195.600 633.440 ;
        RECT 4.000 626.640 1196.000 632.040 ;
        RECT 4.400 625.240 1196.000 626.640 ;
        RECT 4.000 622.560 1196.000 625.240 ;
        RECT 4.000 621.160 1195.600 622.560 ;
        RECT 4.000 615.760 1196.000 621.160 ;
        RECT 4.400 614.360 1196.000 615.760 ;
        RECT 4.000 611.680 1196.000 614.360 ;
        RECT 4.000 610.280 1195.600 611.680 ;
        RECT 4.000 605.560 1196.000 610.280 ;
        RECT 4.400 604.160 1196.000 605.560 ;
        RECT 4.000 600.800 1196.000 604.160 ;
        RECT 4.000 599.400 1195.600 600.800 ;
        RECT 4.000 595.360 1196.000 599.400 ;
        RECT 4.400 593.960 1196.000 595.360 ;
        RECT 4.000 589.920 1196.000 593.960 ;
        RECT 4.000 588.520 1195.600 589.920 ;
        RECT 4.000 584.480 1196.000 588.520 ;
        RECT 4.400 583.080 1196.000 584.480 ;
        RECT 4.000 579.040 1196.000 583.080 ;
        RECT 4.000 577.640 1195.600 579.040 ;
        RECT 4.000 574.280 1196.000 577.640 ;
        RECT 4.400 572.880 1196.000 574.280 ;
        RECT 4.000 567.480 1196.000 572.880 ;
        RECT 4.000 566.080 1195.600 567.480 ;
        RECT 4.000 563.400 1196.000 566.080 ;
        RECT 4.400 562.000 1196.000 563.400 ;
        RECT 4.000 556.600 1196.000 562.000 ;
        RECT 4.000 555.200 1195.600 556.600 ;
        RECT 4.000 553.200 1196.000 555.200 ;
        RECT 4.400 551.800 1196.000 553.200 ;
        RECT 4.000 545.720 1196.000 551.800 ;
        RECT 4.000 544.320 1195.600 545.720 ;
        RECT 4.000 542.320 1196.000 544.320 ;
        RECT 4.400 540.920 1196.000 542.320 ;
        RECT 4.000 534.840 1196.000 540.920 ;
        RECT 4.000 533.440 1195.600 534.840 ;
        RECT 4.000 532.120 1196.000 533.440 ;
        RECT 4.400 530.720 1196.000 532.120 ;
        RECT 4.000 523.960 1196.000 530.720 ;
        RECT 4.000 522.560 1195.600 523.960 ;
        RECT 4.000 521.240 1196.000 522.560 ;
        RECT 4.400 519.840 1196.000 521.240 ;
        RECT 4.000 512.400 1196.000 519.840 ;
        RECT 4.000 511.040 1195.600 512.400 ;
        RECT 4.400 511.000 1195.600 511.040 ;
        RECT 4.400 509.640 1196.000 511.000 ;
        RECT 4.000 501.520 1196.000 509.640 ;
        RECT 4.000 500.160 1195.600 501.520 ;
        RECT 4.400 500.120 1195.600 500.160 ;
        RECT 4.400 498.760 1196.000 500.120 ;
        RECT 4.000 490.640 1196.000 498.760 ;
        RECT 4.000 489.960 1195.600 490.640 ;
        RECT 4.400 489.240 1195.600 489.960 ;
        RECT 4.400 488.560 1196.000 489.240 ;
        RECT 4.000 479.760 1196.000 488.560 ;
        RECT 4.000 479.080 1195.600 479.760 ;
        RECT 4.400 478.360 1195.600 479.080 ;
        RECT 4.400 477.680 1196.000 478.360 ;
        RECT 4.000 468.880 1196.000 477.680 ;
        RECT 4.400 467.480 1195.600 468.880 ;
        RECT 4.000 458.000 1196.000 467.480 ;
        RECT 4.400 457.320 1196.000 458.000 ;
        RECT 4.400 456.600 1195.600 457.320 ;
        RECT 4.000 455.920 1195.600 456.600 ;
        RECT 4.000 447.800 1196.000 455.920 ;
        RECT 4.400 446.440 1196.000 447.800 ;
        RECT 4.400 446.400 1195.600 446.440 ;
        RECT 4.000 445.040 1195.600 446.400 ;
        RECT 4.000 436.920 1196.000 445.040 ;
        RECT 4.400 435.560 1196.000 436.920 ;
        RECT 4.400 435.520 1195.600 435.560 ;
        RECT 4.000 434.160 1195.600 435.520 ;
        RECT 4.000 426.720 1196.000 434.160 ;
        RECT 4.400 425.320 1196.000 426.720 ;
        RECT 4.000 424.680 1196.000 425.320 ;
        RECT 4.000 423.280 1195.600 424.680 ;
        RECT 4.000 415.840 1196.000 423.280 ;
        RECT 4.400 414.440 1196.000 415.840 ;
        RECT 4.000 413.800 1196.000 414.440 ;
        RECT 4.000 412.400 1195.600 413.800 ;
        RECT 4.000 405.640 1196.000 412.400 ;
        RECT 4.400 404.240 1196.000 405.640 ;
        RECT 4.000 402.240 1196.000 404.240 ;
        RECT 4.000 400.840 1195.600 402.240 ;
        RECT 4.000 394.760 1196.000 400.840 ;
        RECT 4.400 393.360 1196.000 394.760 ;
        RECT 4.000 391.360 1196.000 393.360 ;
        RECT 4.000 389.960 1195.600 391.360 ;
        RECT 4.000 384.560 1196.000 389.960 ;
        RECT 4.400 383.160 1196.000 384.560 ;
        RECT 4.000 380.480 1196.000 383.160 ;
        RECT 4.000 379.080 1195.600 380.480 ;
        RECT 4.000 373.680 1196.000 379.080 ;
        RECT 4.400 372.280 1196.000 373.680 ;
        RECT 4.000 369.600 1196.000 372.280 ;
        RECT 4.000 368.200 1195.600 369.600 ;
        RECT 4.000 363.480 1196.000 368.200 ;
        RECT 4.400 362.080 1196.000 363.480 ;
        RECT 4.000 358.720 1196.000 362.080 ;
        RECT 4.000 357.320 1195.600 358.720 ;
        RECT 4.000 352.600 1196.000 357.320 ;
        RECT 4.400 351.200 1196.000 352.600 ;
        RECT 4.000 347.160 1196.000 351.200 ;
        RECT 4.000 345.760 1195.600 347.160 ;
        RECT 4.000 342.400 1196.000 345.760 ;
        RECT 4.400 341.000 1196.000 342.400 ;
        RECT 4.000 336.280 1196.000 341.000 ;
        RECT 4.000 334.880 1195.600 336.280 ;
        RECT 4.000 331.520 1196.000 334.880 ;
        RECT 4.400 330.120 1196.000 331.520 ;
        RECT 4.000 325.400 1196.000 330.120 ;
        RECT 4.000 324.000 1195.600 325.400 ;
        RECT 4.000 321.320 1196.000 324.000 ;
        RECT 4.400 319.920 1196.000 321.320 ;
        RECT 4.000 314.520 1196.000 319.920 ;
        RECT 4.000 313.120 1195.600 314.520 ;
        RECT 4.000 310.440 1196.000 313.120 ;
        RECT 4.400 309.040 1196.000 310.440 ;
        RECT 4.000 303.640 1196.000 309.040 ;
        RECT 4.000 302.240 1195.600 303.640 ;
        RECT 4.000 300.240 1196.000 302.240 ;
        RECT 4.400 298.840 1196.000 300.240 ;
        RECT 4.000 292.760 1196.000 298.840 ;
        RECT 4.000 291.360 1195.600 292.760 ;
        RECT 4.000 290.040 1196.000 291.360 ;
        RECT 4.400 288.640 1196.000 290.040 ;
        RECT 4.000 281.200 1196.000 288.640 ;
        RECT 4.000 279.800 1195.600 281.200 ;
        RECT 4.000 279.160 1196.000 279.800 ;
        RECT 4.400 277.760 1196.000 279.160 ;
        RECT 4.000 270.320 1196.000 277.760 ;
        RECT 4.000 268.960 1195.600 270.320 ;
        RECT 4.400 268.920 1195.600 268.960 ;
        RECT 4.400 267.560 1196.000 268.920 ;
        RECT 4.000 259.440 1196.000 267.560 ;
        RECT 4.000 258.080 1195.600 259.440 ;
        RECT 4.400 258.040 1195.600 258.080 ;
        RECT 4.400 256.680 1196.000 258.040 ;
        RECT 4.000 248.560 1196.000 256.680 ;
        RECT 4.000 247.880 1195.600 248.560 ;
        RECT 4.400 247.160 1195.600 247.880 ;
        RECT 4.400 246.480 1196.000 247.160 ;
        RECT 4.000 237.680 1196.000 246.480 ;
        RECT 4.000 237.000 1195.600 237.680 ;
        RECT 4.400 236.280 1195.600 237.000 ;
        RECT 4.400 235.600 1196.000 236.280 ;
        RECT 4.000 226.800 1196.000 235.600 ;
        RECT 4.400 226.120 1196.000 226.800 ;
        RECT 4.400 225.400 1195.600 226.120 ;
        RECT 4.000 224.720 1195.600 225.400 ;
        RECT 4.000 215.920 1196.000 224.720 ;
        RECT 4.400 215.240 1196.000 215.920 ;
        RECT 4.400 214.520 1195.600 215.240 ;
        RECT 4.000 213.840 1195.600 214.520 ;
        RECT 4.000 205.720 1196.000 213.840 ;
        RECT 4.400 204.360 1196.000 205.720 ;
        RECT 4.400 204.320 1195.600 204.360 ;
        RECT 4.000 202.960 1195.600 204.320 ;
        RECT 4.000 194.840 1196.000 202.960 ;
        RECT 4.400 193.480 1196.000 194.840 ;
        RECT 4.400 193.440 1195.600 193.480 ;
        RECT 4.000 192.080 1195.600 193.440 ;
        RECT 4.000 184.640 1196.000 192.080 ;
        RECT 4.400 183.240 1196.000 184.640 ;
        RECT 4.000 182.600 1196.000 183.240 ;
        RECT 4.000 181.200 1195.600 182.600 ;
        RECT 4.000 173.760 1196.000 181.200 ;
        RECT 4.400 172.360 1196.000 173.760 ;
        RECT 4.000 171.040 1196.000 172.360 ;
        RECT 4.000 169.640 1195.600 171.040 ;
        RECT 4.000 163.560 1196.000 169.640 ;
        RECT 4.400 162.160 1196.000 163.560 ;
        RECT 4.000 160.160 1196.000 162.160 ;
        RECT 4.000 158.760 1195.600 160.160 ;
        RECT 4.000 152.680 1196.000 158.760 ;
        RECT 4.400 151.280 1196.000 152.680 ;
        RECT 4.000 149.280 1196.000 151.280 ;
        RECT 4.000 147.880 1195.600 149.280 ;
        RECT 4.000 142.480 1196.000 147.880 ;
        RECT 4.400 141.080 1196.000 142.480 ;
        RECT 4.000 138.400 1196.000 141.080 ;
        RECT 4.000 137.000 1195.600 138.400 ;
        RECT 4.000 131.600 1196.000 137.000 ;
        RECT 4.400 130.200 1196.000 131.600 ;
        RECT 4.000 127.520 1196.000 130.200 ;
        RECT 4.000 126.120 1195.600 127.520 ;
        RECT 4.000 121.400 1196.000 126.120 ;
        RECT 4.400 120.000 1196.000 121.400 ;
        RECT 4.000 115.960 1196.000 120.000 ;
        RECT 4.000 114.560 1195.600 115.960 ;
        RECT 4.000 110.520 1196.000 114.560 ;
        RECT 4.400 109.120 1196.000 110.520 ;
        RECT 4.000 105.080 1196.000 109.120 ;
        RECT 4.000 103.680 1195.600 105.080 ;
        RECT 4.000 100.320 1196.000 103.680 ;
        RECT 4.400 98.920 1196.000 100.320 ;
        RECT 4.000 94.200 1196.000 98.920 ;
        RECT 4.000 92.800 1195.600 94.200 ;
        RECT 4.000 89.440 1196.000 92.800 ;
        RECT 4.400 88.040 1196.000 89.440 ;
        RECT 4.000 83.320 1196.000 88.040 ;
        RECT 4.000 81.920 1195.600 83.320 ;
        RECT 4.000 79.240 1196.000 81.920 ;
        RECT 4.400 77.840 1196.000 79.240 ;
        RECT 4.000 72.440 1196.000 77.840 ;
        RECT 4.000 71.040 1195.600 72.440 ;
        RECT 4.000 68.360 1196.000 71.040 ;
        RECT 4.400 66.960 1196.000 68.360 ;
        RECT 4.000 60.880 1196.000 66.960 ;
        RECT 4.000 59.480 1195.600 60.880 ;
        RECT 4.000 58.160 1196.000 59.480 ;
        RECT 4.400 56.760 1196.000 58.160 ;
        RECT 4.000 50.000 1196.000 56.760 ;
        RECT 4.000 48.600 1195.600 50.000 ;
        RECT 4.000 47.280 1196.000 48.600 ;
        RECT 4.400 45.880 1196.000 47.280 ;
        RECT 4.000 39.120 1196.000 45.880 ;
        RECT 4.000 37.720 1195.600 39.120 ;
        RECT 4.000 37.080 1196.000 37.720 ;
        RECT 4.400 35.680 1196.000 37.080 ;
        RECT 4.000 28.240 1196.000 35.680 ;
        RECT 4.000 26.840 1195.600 28.240 ;
        RECT 4.000 26.200 1196.000 26.840 ;
        RECT 4.400 24.800 1196.000 26.200 ;
        RECT 4.000 17.360 1196.000 24.800 ;
        RECT 4.000 16.000 1195.600 17.360 ;
        RECT 4.400 15.960 1195.600 16.000 ;
        RECT 4.400 14.600 1196.000 15.960 ;
        RECT 4.000 6.480 1196.000 14.600 ;
        RECT 4.000 5.800 1195.600 6.480 ;
        RECT 4.400 5.080 1195.600 5.800 ;
        RECT 4.400 4.400 1196.000 5.080 ;
        RECT 4.000 4.255 1196.000 4.400 ;
      LAYER met4 ;
        RECT 6.735 10.640 20.640 1188.880 ;
        RECT 23.040 10.640 97.440 1188.880 ;
        RECT 99.840 10.640 1186.505 1188.880 ;
  END
END hs32_core1
END LIBRARY

