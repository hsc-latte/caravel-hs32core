VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2712.230 1200.780 2712.550 1200.840 ;
        RECT 2728.790 1200.780 2729.110 1200.840 ;
        RECT 2712.230 1200.640 2729.110 1200.780 ;
        RECT 2712.230 1200.580 2712.550 1200.640 ;
        RECT 2728.790 1200.580 2729.110 1200.640 ;
        RECT 2728.790 89.660 2729.110 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 2728.790 89.520 2899.310 89.660 ;
        RECT 2728.790 89.460 2729.110 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 2712.260 1200.580 2712.520 1200.840 ;
        RECT 2728.820 1200.580 2729.080 1200.840 ;
        RECT 2728.820 89.460 2729.080 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 2712.250 1205.115 2712.530 1205.485 ;
        RECT 2712.320 1200.870 2712.460 1205.115 ;
        RECT 2712.260 1200.550 2712.520 1200.870 ;
        RECT 2728.820 1200.550 2729.080 1200.870 ;
        RECT 2728.880 89.750 2729.020 1200.550 ;
        RECT 2728.820 89.430 2729.080 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2712.250 1205.160 2712.530 1205.440 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2712.225 1205.450 2712.555 1205.465 ;
        RECT 2699.740 1205.400 2712.555 1205.450 ;
        RECT 2696.000 1205.150 2712.555 1205.400 ;
        RECT 2696.000 1204.800 2700.000 1205.150 ;
        RECT 2712.225 1205.135 2712.555 1205.150 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2722.810 2429.200 2723.130 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 2722.810 2429.060 2901.150 2429.200 ;
        RECT 2722.810 2429.000 2723.130 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 2713.150 1524.460 2713.470 1524.520 ;
        RECT 2722.810 1524.460 2723.130 1524.520 ;
        RECT 2713.150 1524.320 2723.130 1524.460 ;
        RECT 2713.150 1524.260 2713.470 1524.320 ;
        RECT 2722.810 1524.260 2723.130 1524.320 ;
      LAYER via ;
        RECT 2722.840 2429.000 2723.100 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 2713.180 1524.260 2713.440 1524.520 ;
        RECT 2722.840 1524.260 2723.100 1524.520 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 2722.840 2428.970 2723.100 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 2722.900 1524.550 2723.040 2428.970 ;
        RECT 2713.180 1524.230 2713.440 1524.550 ;
        RECT 2722.840 1524.230 2723.100 1524.550 ;
        RECT 2713.240 1521.005 2713.380 1524.230 ;
        RECT 2713.170 1520.635 2713.450 1521.005 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
        RECT 2713.170 1520.680 2713.450 1520.960 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2713.145 1520.970 2713.475 1520.985 ;
        RECT 2699.740 1520.920 2713.475 1520.970 ;
        RECT 2696.000 1520.670 2713.475 1520.920 ;
        RECT 2696.000 1520.320 2700.000 1520.670 ;
        RECT 2713.145 1520.655 2713.475 1520.670 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2722.350 2663.800 2722.670 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 2722.350 2663.660 2901.150 2663.800 ;
        RECT 2722.350 2663.600 2722.670 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 2713.150 1549.960 2713.470 1550.020 ;
        RECT 2722.350 1549.960 2722.670 1550.020 ;
        RECT 2713.150 1549.820 2722.670 1549.960 ;
        RECT 2713.150 1549.760 2713.470 1549.820 ;
        RECT 2722.350 1549.760 2722.670 1549.820 ;
      LAYER via ;
        RECT 2722.380 2663.600 2722.640 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 2713.180 1549.760 2713.440 1550.020 ;
        RECT 2722.380 1549.760 2722.640 1550.020 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 2722.380 2663.570 2722.640 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 2713.170 1551.915 2713.450 1552.285 ;
        RECT 2713.240 1550.050 2713.380 1551.915 ;
        RECT 2722.440 1550.050 2722.580 2663.570 ;
        RECT 2713.180 1549.730 2713.440 1550.050 ;
        RECT 2722.380 1549.730 2722.640 1550.050 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
        RECT 2713.170 1551.960 2713.450 1552.240 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2713.145 1552.250 2713.475 1552.265 ;
        RECT 2699.740 1552.200 2713.475 1552.250 ;
        RECT 2696.000 1551.950 2713.475 1552.200 ;
        RECT 2696.000 1551.600 2700.000 1551.950 ;
        RECT 2713.145 1551.935 2713.475 1551.950 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2721.890 2898.400 2722.210 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 2721.890 2898.260 2901.150 2898.400 ;
        RECT 2721.890 2898.200 2722.210 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
        RECT 2713.150 1584.640 2713.470 1584.700 ;
        RECT 2721.890 1584.640 2722.210 1584.700 ;
        RECT 2713.150 1584.500 2722.210 1584.640 ;
        RECT 2713.150 1584.440 2713.470 1584.500 ;
        RECT 2721.890 1584.440 2722.210 1584.500 ;
      LAYER via ;
        RECT 2721.920 2898.200 2722.180 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
        RECT 2713.180 1584.440 2713.440 1584.700 ;
        RECT 2721.920 1584.440 2722.180 1584.700 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 2721.920 2898.170 2722.180 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 2721.980 1584.730 2722.120 2898.170 ;
        RECT 2713.180 1584.410 2713.440 1584.730 ;
        RECT 2721.920 1584.410 2722.180 1584.730 ;
        RECT 2713.240 1584.245 2713.380 1584.410 ;
        RECT 2713.170 1583.875 2713.450 1584.245 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
        RECT 2713.170 1583.920 2713.450 1584.200 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
        RECT 2713.145 1584.210 2713.475 1584.225 ;
        RECT 2699.740 1584.160 2713.475 1584.210 ;
        RECT 2696.000 1583.910 2713.475 1584.160 ;
        RECT 2696.000 1583.560 2700.000 1583.910 ;
        RECT 2713.145 1583.895 2713.475 1583.910 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2728.790 3133.000 2729.110 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 2728.790 3132.860 2901.150 3133.000 ;
        RECT 2728.790 3132.800 2729.110 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
        RECT 2713.150 1621.020 2713.470 1621.080 ;
        RECT 2728.790 1621.020 2729.110 1621.080 ;
        RECT 2713.150 1620.880 2729.110 1621.020 ;
        RECT 2713.150 1620.820 2713.470 1620.880 ;
        RECT 2728.790 1620.820 2729.110 1620.880 ;
      LAYER via ;
        RECT 2728.820 3132.800 2729.080 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
        RECT 2713.180 1620.820 2713.440 1621.080 ;
        RECT 2728.820 1620.820 2729.080 1621.080 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 2728.820 3132.770 2729.080 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 2728.880 1621.110 2729.020 3132.770 ;
        RECT 2713.180 1620.790 2713.440 1621.110 ;
        RECT 2728.820 1620.790 2729.080 1621.110 ;
        RECT 2713.240 1615.525 2713.380 1620.790 ;
        RECT 2713.170 1615.155 2713.450 1615.525 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
        RECT 2713.170 1615.200 2713.450 1615.480 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
        RECT 2713.145 1615.490 2713.475 1615.505 ;
        RECT 2699.740 1615.440 2713.475 1615.490 ;
        RECT 2696.000 1615.190 2713.475 1615.440 ;
        RECT 2696.000 1614.840 2700.000 1615.190 ;
        RECT 2713.145 1615.175 2713.475 1615.190 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2735.690 3367.600 2736.010 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 2735.690 3367.460 2901.150 3367.600 ;
        RECT 2735.690 3367.400 2736.010 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
        RECT 2713.150 1644.480 2713.470 1644.540 ;
        RECT 2735.690 1644.480 2736.010 1644.540 ;
        RECT 2713.150 1644.340 2736.010 1644.480 ;
        RECT 2713.150 1644.280 2713.470 1644.340 ;
        RECT 2735.690 1644.280 2736.010 1644.340 ;
      LAYER via ;
        RECT 2735.720 3367.400 2735.980 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
        RECT 2713.180 1644.280 2713.440 1644.540 ;
        RECT 2735.720 1644.280 2735.980 1644.540 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 2735.720 3367.370 2735.980 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 2713.170 1647.115 2713.450 1647.485 ;
        RECT 2713.240 1644.570 2713.380 1647.115 ;
        RECT 2735.780 1644.570 2735.920 3367.370 ;
        RECT 2713.180 1644.250 2713.440 1644.570 ;
        RECT 2735.720 1644.250 2735.980 1644.570 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
        RECT 2713.170 1647.160 2713.450 1647.440 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
        RECT 2713.145 1647.450 2713.475 1647.465 ;
        RECT 2699.740 1647.400 2713.475 1647.450 ;
        RECT 2696.000 1647.150 2713.475 1647.400 ;
        RECT 2696.000 1646.800 2700.000 1647.150 ;
        RECT 2713.145 1647.135 2713.475 1647.150 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2749.490 3501.560 2749.810 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 2749.490 3501.420 2798.570 3501.560 ;
        RECT 2749.490 3501.360 2749.810 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
        RECT 2713.150 1681.200 2713.470 1681.260 ;
        RECT 2749.490 1681.200 2749.810 1681.260 ;
        RECT 2713.150 1681.060 2749.810 1681.200 ;
        RECT 2713.150 1681.000 2713.470 1681.060 ;
        RECT 2749.490 1681.000 2749.810 1681.060 ;
      LAYER via ;
        RECT 2749.520 3501.360 2749.780 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
        RECT 2713.180 1681.000 2713.440 1681.260 ;
        RECT 2749.520 1681.000 2749.780 1681.260 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 2749.520 3501.330 2749.780 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 2749.580 1681.290 2749.720 3501.330 ;
        RECT 2713.180 1680.970 2713.440 1681.290 ;
        RECT 2749.520 1680.970 2749.780 1681.290 ;
        RECT 2713.240 1678.765 2713.380 1680.970 ;
        RECT 2713.170 1678.395 2713.450 1678.765 ;
      LAYER via2 ;
        RECT 2713.170 1678.440 2713.450 1678.720 ;
      LAYER met3 ;
        RECT 2713.145 1678.730 2713.475 1678.745 ;
        RECT 2699.740 1678.680 2713.475 1678.730 ;
        RECT 2696.000 1678.430 2713.475 1678.680 ;
        RECT 2696.000 1678.080 2700.000 1678.430 ;
        RECT 2713.145 1678.415 2713.475 1678.430 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2473.950 3499.180 2474.270 3499.240 ;
        RECT 2476.710 3499.180 2477.030 3499.240 ;
        RECT 2473.950 3499.040 2477.030 3499.180 ;
        RECT 2473.950 3498.980 2474.270 3499.040 ;
        RECT 2476.710 3498.980 2477.030 3499.040 ;
        RECT 2476.710 3054.120 2477.030 3054.180 ;
        RECT 2706.710 3054.120 2707.030 3054.180 ;
        RECT 2476.710 3053.980 2707.030 3054.120 ;
        RECT 2476.710 3053.920 2477.030 3053.980 ;
        RECT 2706.710 3053.920 2707.030 3053.980 ;
      LAYER via ;
        RECT 2473.980 3498.980 2474.240 3499.240 ;
        RECT 2476.740 3498.980 2477.000 3499.240 ;
        RECT 2476.740 3053.920 2477.000 3054.180 ;
        RECT 2706.740 3053.920 2707.000 3054.180 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3499.270 2474.180 3517.600 ;
        RECT 2473.980 3498.950 2474.240 3499.270 ;
        RECT 2476.740 3498.950 2477.000 3499.270 ;
        RECT 2476.800 3054.210 2476.940 3498.950 ;
        RECT 2476.740 3053.890 2477.000 3054.210 ;
        RECT 2706.740 3053.890 2707.000 3054.210 ;
        RECT 2706.800 1710.725 2706.940 3053.890 ;
        RECT 2706.730 1710.355 2707.010 1710.725 ;
      LAYER via2 ;
        RECT 2706.730 1710.400 2707.010 1710.680 ;
      LAYER met3 ;
        RECT 2706.705 1710.690 2707.035 1710.705 ;
        RECT 2699.740 1710.640 2707.035 1710.690 ;
        RECT 2696.000 1710.390 2707.035 1710.640 ;
        RECT 2696.000 1710.040 2700.000 1710.390 ;
        RECT 2706.705 1710.375 2707.035 1710.390 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2149.190 3498.500 2149.510 3498.560 ;
        RECT 2152.410 3498.500 2152.730 3498.560 ;
        RECT 2149.190 3498.360 2152.730 3498.500 ;
        RECT 2149.190 3498.300 2149.510 3498.360 ;
        RECT 2152.410 3498.300 2152.730 3498.360 ;
        RECT 2152.410 3053.440 2152.730 3053.500 ;
        RECT 2707.170 3053.440 2707.490 3053.500 ;
        RECT 2152.410 3053.300 2707.490 3053.440 ;
        RECT 2152.410 3053.240 2152.730 3053.300 ;
        RECT 2707.170 3053.240 2707.490 3053.300 ;
      LAYER via ;
        RECT 2149.220 3498.300 2149.480 3498.560 ;
        RECT 2152.440 3498.300 2152.700 3498.560 ;
        RECT 2152.440 3053.240 2152.700 3053.500 ;
        RECT 2707.200 3053.240 2707.460 3053.500 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3498.590 2149.420 3517.600 ;
        RECT 2149.220 3498.270 2149.480 3498.590 ;
        RECT 2152.440 3498.270 2152.700 3498.590 ;
        RECT 2152.500 3053.530 2152.640 3498.270 ;
        RECT 2152.440 3053.210 2152.700 3053.530 ;
        RECT 2707.200 3053.210 2707.460 3053.530 ;
        RECT 2707.260 1742.005 2707.400 3053.210 ;
        RECT 2707.190 1741.635 2707.470 1742.005 ;
      LAYER via2 ;
        RECT 2707.190 1741.680 2707.470 1741.960 ;
      LAYER met3 ;
        RECT 2707.165 1741.970 2707.495 1741.985 ;
        RECT 2699.740 1741.920 2707.495 1741.970 ;
        RECT 2696.000 1741.670 2707.495 1741.920 ;
        RECT 2696.000 1741.320 2700.000 1741.670 ;
        RECT 2707.165 1741.655 2707.495 1741.670 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1824.890 3498.500 1825.210 3498.560 ;
        RECT 1828.110 3498.500 1828.430 3498.560 ;
        RECT 1824.890 3498.360 1828.430 3498.500 ;
        RECT 1824.890 3498.300 1825.210 3498.360 ;
        RECT 1828.110 3498.300 1828.430 3498.360 ;
        RECT 1828.110 3053.100 1828.430 3053.160 ;
        RECT 2707.630 3053.100 2707.950 3053.160 ;
        RECT 1828.110 3052.960 2707.950 3053.100 ;
        RECT 1828.110 3052.900 1828.430 3052.960 ;
        RECT 2707.630 3052.900 2707.950 3052.960 ;
      LAYER via ;
        RECT 1824.920 3498.300 1825.180 3498.560 ;
        RECT 1828.140 3498.300 1828.400 3498.560 ;
        RECT 1828.140 3052.900 1828.400 3053.160 ;
        RECT 2707.660 3052.900 2707.920 3053.160 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3498.590 1825.120 3517.600 ;
        RECT 1824.920 3498.270 1825.180 3498.590 ;
        RECT 1828.140 3498.270 1828.400 3498.590 ;
        RECT 1828.200 3053.190 1828.340 3498.270 ;
        RECT 1828.140 3052.870 1828.400 3053.190 ;
        RECT 2707.660 3052.870 2707.920 3053.190 ;
        RECT 2707.720 1773.965 2707.860 3052.870 ;
        RECT 2707.650 1773.595 2707.930 1773.965 ;
      LAYER via2 ;
        RECT 2707.650 1773.640 2707.930 1773.920 ;
      LAYER met3 ;
        RECT 2707.625 1773.930 2707.955 1773.945 ;
        RECT 2699.740 1773.880 2707.955 1773.930 ;
        RECT 2696.000 1773.630 2707.955 1773.880 ;
        RECT 2696.000 1773.280 2700.000 1773.630 ;
        RECT 2707.625 1773.615 2707.955 1773.630 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 2398.940 1504.130 2399.000 ;
        RECT 2709.470 2398.940 2709.790 2399.000 ;
        RECT 1503.810 2398.800 2709.790 2398.940 ;
        RECT 1503.810 2398.740 1504.130 2398.800 ;
        RECT 2709.470 2398.740 2709.790 2398.800 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 2398.740 1504.100 2399.000 ;
        RECT 2709.500 2398.740 2709.760 2399.000 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 2399.030 1504.040 3498.270 ;
        RECT 1503.840 2398.710 1504.100 2399.030 ;
        RECT 2709.500 2398.710 2709.760 2399.030 ;
        RECT 2709.560 1805.245 2709.700 2398.710 ;
        RECT 2709.490 1804.875 2709.770 1805.245 ;
      LAYER via2 ;
        RECT 2709.490 1804.920 2709.770 1805.200 ;
      LAYER met3 ;
        RECT 2709.465 1805.210 2709.795 1805.225 ;
        RECT 2699.740 1805.160 2709.795 1805.210 ;
        RECT 2696.000 1804.910 2709.795 1805.160 ;
        RECT 2696.000 1804.560 2700.000 1804.910 ;
        RECT 2709.465 1804.895 2709.795 1804.910 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1235.460 2713.470 1235.520 ;
        RECT 2735.690 1235.460 2736.010 1235.520 ;
        RECT 2713.150 1235.320 2736.010 1235.460 ;
        RECT 2713.150 1235.260 2713.470 1235.320 ;
        RECT 2735.690 1235.260 2736.010 1235.320 ;
        RECT 2735.690 324.260 2736.010 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 2735.690 324.120 2899.310 324.260 ;
        RECT 2735.690 324.060 2736.010 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 2713.180 1235.260 2713.440 1235.520 ;
        RECT 2735.720 1235.260 2735.980 1235.520 ;
        RECT 2735.720 324.060 2735.980 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 2713.170 1236.395 2713.450 1236.765 ;
        RECT 2713.240 1235.550 2713.380 1236.395 ;
        RECT 2713.180 1235.230 2713.440 1235.550 ;
        RECT 2735.720 1235.230 2735.980 1235.550 ;
        RECT 2735.780 324.350 2735.920 1235.230 ;
        RECT 2735.720 324.030 2735.980 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2713.170 1236.440 2713.450 1236.720 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2713.145 1236.730 2713.475 1236.745 ;
        RECT 2699.740 1236.680 2713.475 1236.730 ;
        RECT 2696.000 1236.430 2713.475 1236.680 ;
        RECT 2696.000 1236.080 2700.000 1236.430 ;
        RECT 2713.145 1236.415 2713.475 1236.430 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3503.260 1176.150 3503.320 ;
        RECT 1179.510 3503.260 1179.830 3503.320 ;
        RECT 1175.830 3503.120 1179.830 3503.260 ;
        RECT 1175.830 3503.060 1176.150 3503.120 ;
        RECT 1179.510 3503.060 1179.830 3503.120 ;
        RECT 1179.510 2398.600 1179.830 2398.660 ;
        RECT 2709.930 2398.600 2710.250 2398.660 ;
        RECT 1179.510 2398.460 2710.250 2398.600 ;
        RECT 1179.510 2398.400 1179.830 2398.460 ;
        RECT 2709.930 2398.400 2710.250 2398.460 ;
      LAYER via ;
        RECT 1175.860 3503.060 1176.120 3503.320 ;
        RECT 1179.540 3503.060 1179.800 3503.320 ;
        RECT 1179.540 2398.400 1179.800 2398.660 ;
        RECT 2709.960 2398.400 2710.220 2398.660 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3503.350 1176.060 3517.600 ;
        RECT 1175.860 3503.030 1176.120 3503.350 ;
        RECT 1179.540 3503.030 1179.800 3503.350 ;
        RECT 1179.600 2398.690 1179.740 3503.030 ;
        RECT 1179.540 2398.370 1179.800 2398.690 ;
        RECT 2709.960 2398.370 2710.220 2398.690 ;
        RECT 2710.020 1836.525 2710.160 2398.370 ;
        RECT 2709.950 1836.155 2710.230 1836.525 ;
      LAYER via2 ;
        RECT 2709.950 1836.200 2710.230 1836.480 ;
      LAYER met3 ;
        RECT 2709.925 1836.490 2710.255 1836.505 ;
        RECT 2699.740 1836.440 2710.255 1836.490 ;
        RECT 2696.000 1836.190 2710.255 1836.440 ;
        RECT 2696.000 1835.840 2700.000 1836.190 ;
        RECT 2709.925 1836.175 2710.255 1836.190 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3498.500 851.850 3498.560 ;
        RECT 855.210 3498.500 855.530 3498.560 ;
        RECT 851.530 3498.360 855.530 3498.500 ;
        RECT 851.530 3498.300 851.850 3498.360 ;
        RECT 855.210 3498.300 855.530 3498.360 ;
        RECT 855.210 2398.260 855.530 2398.320 ;
        RECT 2710.390 2398.260 2710.710 2398.320 ;
        RECT 855.210 2398.120 2710.710 2398.260 ;
        RECT 855.210 2398.060 855.530 2398.120 ;
        RECT 2710.390 2398.060 2710.710 2398.120 ;
      LAYER via ;
        RECT 851.560 3498.300 851.820 3498.560 ;
        RECT 855.240 3498.300 855.500 3498.560 ;
        RECT 855.240 2398.060 855.500 2398.320 ;
        RECT 2710.420 2398.060 2710.680 2398.320 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3498.590 851.760 3517.600 ;
        RECT 851.560 3498.270 851.820 3498.590 ;
        RECT 855.240 3498.270 855.500 3498.590 ;
        RECT 855.300 2398.350 855.440 3498.270 ;
        RECT 855.240 2398.030 855.500 2398.350 ;
        RECT 2710.420 2398.030 2710.680 2398.350 ;
        RECT 2710.480 1868.485 2710.620 2398.030 ;
        RECT 2710.410 1868.115 2710.690 1868.485 ;
      LAYER via2 ;
        RECT 2710.410 1868.160 2710.690 1868.440 ;
      LAYER met3 ;
        RECT 2710.385 1868.450 2710.715 1868.465 ;
        RECT 2699.740 1868.400 2710.715 1868.450 ;
        RECT 2696.000 1868.150 2710.715 1868.400 ;
        RECT 2696.000 1867.800 2700.000 1868.150 ;
        RECT 2710.385 1868.135 2710.715 1868.150 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 2397.920 531.230 2397.980 ;
        RECT 2710.850 2397.920 2711.170 2397.980 ;
        RECT 530.910 2397.780 2711.170 2397.920 ;
        RECT 530.910 2397.720 531.230 2397.780 ;
        RECT 2710.850 2397.720 2711.170 2397.780 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 2397.720 531.200 2397.980 ;
        RECT 2710.880 2397.720 2711.140 2397.980 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 2398.010 531.140 3498.270 ;
        RECT 530.940 2397.690 531.200 2398.010 ;
        RECT 2710.880 2397.690 2711.140 2398.010 ;
        RECT 2710.940 1899.765 2711.080 2397.690 ;
        RECT 2710.870 1899.395 2711.150 1899.765 ;
      LAYER via2 ;
        RECT 2710.870 1899.440 2711.150 1899.720 ;
      LAYER met3 ;
        RECT 2710.845 1899.730 2711.175 1899.745 ;
        RECT 2699.740 1899.680 2711.175 1899.730 ;
        RECT 2696.000 1899.430 2711.175 1899.680 ;
        RECT 2696.000 1899.080 2700.000 1899.430 ;
        RECT 2710.845 1899.415 2711.175 1899.430 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.560 202.790 3501.620 ;
        RECT 2705.330 3501.560 2705.650 3501.620 ;
        RECT 202.470 3501.420 2705.650 3501.560 ;
        RECT 202.470 3501.360 202.790 3501.420 ;
        RECT 2705.330 3501.360 2705.650 3501.420 ;
      LAYER via ;
        RECT 202.500 3501.360 202.760 3501.620 ;
        RECT 2705.360 3501.360 2705.620 3501.620 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.650 202.700 3517.600 ;
        RECT 202.500 3501.330 202.760 3501.650 ;
        RECT 2705.360 3501.330 2705.620 3501.650 ;
        RECT 2705.420 1931.725 2705.560 3501.330 ;
        RECT 2705.350 1931.355 2705.630 1931.725 ;
      LAYER via2 ;
        RECT 2705.350 1931.400 2705.630 1931.680 ;
      LAYER met3 ;
        RECT 2705.325 1931.690 2705.655 1931.705 ;
        RECT 2699.740 1931.640 2705.655 1931.690 ;
        RECT 2696.000 1931.390 2705.655 1931.640 ;
        RECT 2696.000 1931.040 2700.000 1931.390 ;
        RECT 2705.325 1931.375 2705.655 1931.390 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 2705.790 3408.740 2706.110 3408.800 ;
        RECT 17.550 3408.600 2706.110 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 2705.790 3408.540 2706.110 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 2705.820 3408.540 2706.080 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 2705.820 3408.510 2706.080 3408.830 ;
        RECT 2705.880 1963.005 2706.020 3408.510 ;
        RECT 2705.810 1962.635 2706.090 1963.005 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
        RECT 2705.810 1962.680 2706.090 1962.960 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
        RECT 2705.785 1962.970 2706.115 1962.985 ;
        RECT 2699.740 1962.920 2706.115 1962.970 ;
        RECT 2696.000 1962.670 2706.115 1962.920 ;
        RECT 2696.000 1962.320 2700.000 1962.670 ;
        RECT 2705.785 1962.655 2706.115 1962.670 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.005 17.320 3124.075 ;
        RECT 17.110 3118.635 17.390 3119.005 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
        RECT 17.110 3118.680 17.390 3118.960 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
        RECT 17.085 3118.970 17.415 3118.985 ;
        RECT 2694.030 3118.970 2694.410 3118.980 ;
        RECT 17.085 3118.670 2694.410 3118.970 ;
        RECT 17.085 3118.655 17.415 3118.670 ;
        RECT 2694.030 3118.660 2694.410 3118.670 ;
        RECT 2696.790 2075.170 2697.170 2075.180 ;
        RECT 2696.790 2074.870 2699.890 2075.170 ;
        RECT 2696.790 2074.860 2697.170 2074.870 ;
        RECT 2696.790 2069.050 2697.170 2069.060 ;
        RECT 2699.590 2069.050 2699.890 2074.870 ;
        RECT 2696.790 2068.750 2699.890 2069.050 ;
        RECT 2696.790 2068.740 2697.170 2068.750 ;
        RECT 2696.790 1997.340 2697.170 1997.660 ;
        RECT 2696.830 1994.880 2697.130 1997.340 ;
        RECT 2696.000 1994.280 2700.000 1994.880 ;
      LAYER via3 ;
        RECT 2694.060 3118.660 2694.380 3118.980 ;
        RECT 2696.820 2074.860 2697.140 2075.180 ;
        RECT 2696.820 2068.740 2697.140 2069.060 ;
        RECT 2696.820 1997.340 2697.140 1997.660 ;
      LAYER met4 ;
        RECT 2694.055 3118.655 2694.385 3118.985 ;
        RECT 2694.070 2188.050 2694.370 3118.655 ;
        RECT 2693.150 2187.750 2694.370 2188.050 ;
        RECT 2693.150 2181.250 2693.450 2187.750 ;
        RECT 2693.150 2180.950 2694.370 2181.250 ;
        RECT 2694.070 2082.650 2694.370 2180.950 ;
        RECT 2694.070 2082.350 2696.210 2082.650 ;
        RECT 2695.910 2075.170 2696.210 2082.350 ;
        RECT 2696.815 2075.170 2697.145 2075.185 ;
        RECT 2695.910 2074.870 2697.145 2075.170 ;
        RECT 2696.815 2074.855 2697.145 2074.870 ;
        RECT 2696.815 2069.050 2697.145 2069.065 ;
        RECT 2695.910 2068.750 2697.145 2069.050 ;
        RECT 2695.910 2065.650 2696.210 2068.750 ;
        RECT 2696.815 2068.735 2697.145 2068.750 ;
        RECT 2694.070 2065.350 2696.210 2065.650 ;
        RECT 2694.070 2018.730 2694.370 2065.350 ;
        RECT 2694.070 2018.430 2695.290 2018.730 ;
        RECT 2694.990 1997.650 2695.290 2018.430 ;
        RECT 2696.815 1997.650 2697.145 1997.665 ;
        RECT 2694.990 1997.350 2697.145 1997.650 ;
        RECT 2696.815 1997.335 2697.145 1997.350 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 2397.580 17.870 2397.640 ;
        RECT 2702.570 2397.580 2702.890 2397.640 ;
        RECT 17.550 2397.440 2702.890 2397.580 ;
        RECT 17.550 2397.380 17.870 2397.440 ;
        RECT 2702.570 2397.380 2702.890 2397.440 ;
      LAYER via ;
        RECT 17.580 2397.380 17.840 2397.640 ;
        RECT 2702.600 2397.380 2702.860 2397.640 ;
      LAYER met2 ;
        RECT 17.570 2836.435 17.850 2836.805 ;
        RECT 17.640 2397.670 17.780 2836.435 ;
        RECT 17.580 2397.350 17.840 2397.670 ;
        RECT 2702.600 2397.350 2702.860 2397.670 ;
        RECT 2702.660 2026.245 2702.800 2397.350 ;
        RECT 2702.590 2025.875 2702.870 2026.245 ;
      LAYER via2 ;
        RECT 17.570 2836.480 17.850 2836.760 ;
        RECT 2702.590 2025.920 2702.870 2026.200 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 17.545 2836.770 17.875 2836.785 ;
        RECT -4.800 2836.470 17.875 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 17.545 2836.455 17.875 2836.470 ;
        RECT 2702.565 2026.210 2702.895 2026.225 ;
        RECT 2699.740 2026.160 2702.895 2026.210 ;
        RECT 2696.000 2025.910 2702.895 2026.160 ;
        RECT 2696.000 2025.560 2700.000 2025.910 ;
        RECT 2702.565 2025.895 2702.895 2025.910 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2546.500 16.490 2546.560 ;
        RECT 2697.510 2546.500 2697.830 2546.560 ;
        RECT 16.170 2546.360 2697.830 2546.500 ;
        RECT 16.170 2546.300 16.490 2546.360 ;
        RECT 2697.510 2546.300 2697.830 2546.360 ;
      LAYER via ;
        RECT 16.200 2546.300 16.460 2546.560 ;
        RECT 2697.540 2546.300 2697.800 2546.560 ;
      LAYER met2 ;
        RECT 16.190 2549.475 16.470 2549.845 ;
        RECT 16.260 2546.590 16.400 2549.475 ;
        RECT 16.200 2546.270 16.460 2546.590 ;
        RECT 2697.540 2546.270 2697.800 2546.590 ;
        RECT 2697.600 2060.925 2697.740 2546.270 ;
        RECT 2697.530 2060.555 2697.810 2060.925 ;
      LAYER via2 ;
        RECT 16.190 2549.520 16.470 2549.800 ;
        RECT 2697.530 2060.600 2697.810 2060.880 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 16.165 2549.810 16.495 2549.825 ;
        RECT -4.800 2549.510 16.495 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 16.165 2549.495 16.495 2549.510 ;
        RECT 2697.505 2060.890 2697.835 2060.905 ;
        RECT 2697.505 2060.575 2698.050 2060.890 ;
        RECT 2697.750 2058.120 2698.050 2060.575 ;
        RECT 2696.000 2057.520 2700.000 2058.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1299.110 2392.820 1299.430 2392.880 ;
        RECT 2703.490 2392.820 2703.810 2392.880 ;
        RECT 1299.110 2392.680 2703.810 2392.820 ;
        RECT 1299.110 2392.620 1299.430 2392.680 ;
        RECT 2703.490 2392.620 2703.810 2392.680 ;
        RECT 17.090 2262.940 17.410 2263.000 ;
        RECT 1299.110 2262.940 1299.430 2263.000 ;
        RECT 17.090 2262.800 1299.430 2262.940 ;
        RECT 17.090 2262.740 17.410 2262.800 ;
        RECT 1299.110 2262.740 1299.430 2262.800 ;
      LAYER via ;
        RECT 1299.140 2392.620 1299.400 2392.880 ;
        RECT 2703.520 2392.620 2703.780 2392.880 ;
        RECT 17.120 2262.740 17.380 2263.000 ;
        RECT 1299.140 2262.740 1299.400 2263.000 ;
      LAYER met2 ;
        RECT 1299.140 2392.590 1299.400 2392.910 ;
        RECT 2703.520 2392.590 2703.780 2392.910 ;
        RECT 1299.200 2263.030 1299.340 2392.590 ;
        RECT 17.120 2262.710 17.380 2263.030 ;
        RECT 1299.140 2262.710 1299.400 2263.030 ;
        RECT 17.180 2262.205 17.320 2262.710 ;
        RECT 17.110 2261.835 17.390 2262.205 ;
        RECT 2703.580 2089.485 2703.720 2392.590 ;
        RECT 2703.510 2089.115 2703.790 2089.485 ;
      LAYER via2 ;
        RECT 17.110 2261.880 17.390 2262.160 ;
        RECT 2703.510 2089.160 2703.790 2089.440 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 17.085 2262.170 17.415 2262.185 ;
        RECT -4.800 2261.870 17.415 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 17.085 2261.855 17.415 2261.870 ;
        RECT 2703.485 2089.450 2703.815 2089.465 ;
        RECT 2699.740 2089.400 2703.815 2089.450 ;
        RECT 2696.000 2089.150 2703.815 2089.400 ;
        RECT 2696.000 2088.800 2700.000 2089.150 ;
        RECT 2703.485 2089.135 2703.815 2089.150 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1303.710 2392.480 1304.030 2392.540 ;
        RECT 2713.610 2392.480 2713.930 2392.540 ;
        RECT 1303.710 2392.340 2713.930 2392.480 ;
        RECT 1303.710 2392.280 1304.030 2392.340 ;
        RECT 2713.610 2392.280 2713.930 2392.340 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 1303.710 1980.060 1304.030 1980.120 ;
        RECT 15.710 1979.920 1304.030 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 1303.710 1979.860 1304.030 1979.920 ;
      LAYER via ;
        RECT 1303.740 2392.280 1304.000 2392.540 ;
        RECT 2713.640 2392.280 2713.900 2392.540 ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 1303.740 1979.860 1304.000 1980.120 ;
      LAYER met2 ;
        RECT 1303.740 2392.250 1304.000 2392.570 ;
        RECT 2713.640 2392.250 2713.900 2392.570 ;
        RECT 1303.800 1980.150 1303.940 2392.250 ;
        RECT 2713.700 2120.765 2713.840 2392.250 ;
        RECT 2713.630 2120.395 2713.910 2120.765 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 1303.740 1979.830 1304.000 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 2713.630 2120.440 2713.910 2120.720 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT 2713.605 2120.730 2713.935 2120.745 ;
        RECT 2699.740 2120.680 2713.935 2120.730 ;
        RECT 2696.000 2120.430 2713.935 2120.680 ;
        RECT 2696.000 2120.080 2700.000 2120.430 ;
        RECT 2713.605 2120.415 2713.935 2120.430 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1263.000 2713.470 1263.060 ;
        RECT 2749.490 1263.000 2749.810 1263.060 ;
        RECT 2713.150 1262.860 2749.810 1263.000 ;
        RECT 2713.150 1262.800 2713.470 1262.860 ;
        RECT 2749.490 1262.800 2749.810 1262.860 ;
        RECT 2749.490 558.860 2749.810 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 2749.490 558.720 2899.310 558.860 ;
        RECT 2749.490 558.660 2749.810 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 2713.180 1262.800 2713.440 1263.060 ;
        RECT 2749.520 1262.800 2749.780 1263.060 ;
        RECT 2749.520 558.660 2749.780 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 2713.170 1267.675 2713.450 1268.045 ;
        RECT 2713.240 1263.090 2713.380 1267.675 ;
        RECT 2713.180 1262.770 2713.440 1263.090 ;
        RECT 2749.520 1262.770 2749.780 1263.090 ;
        RECT 2749.580 558.950 2749.720 1262.770 ;
        RECT 2749.520 558.630 2749.780 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2713.170 1267.720 2713.450 1268.000 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2713.145 1268.010 2713.475 1268.025 ;
        RECT 2699.740 1267.960 2713.475 1268.010 ;
        RECT 2696.000 1267.710 2713.475 1267.960 ;
        RECT 2696.000 1267.360 2700.000 1267.710 ;
        RECT 2713.145 1267.695 2713.475 1267.710 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1302.330 2392.140 1302.650 2392.200 ;
        RECT 2713.150 2392.140 2713.470 2392.200 ;
        RECT 1302.330 2392.000 2713.470 2392.140 ;
        RECT 1302.330 2391.940 1302.650 2392.000 ;
        RECT 2713.150 2391.940 2713.470 2392.000 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 1302.330 1690.380 1302.650 1690.440 ;
        RECT 17.090 1690.240 1302.650 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 1302.330 1690.180 1302.650 1690.240 ;
      LAYER via ;
        RECT 1302.360 2391.940 1302.620 2392.200 ;
        RECT 2713.180 2391.940 2713.440 2392.200 ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 1302.360 1690.180 1302.620 1690.440 ;
      LAYER met2 ;
        RECT 1302.360 2391.910 1302.620 2392.230 ;
        RECT 2713.180 2391.910 2713.440 2392.230 ;
        RECT 1302.420 1690.470 1302.560 2391.910 ;
        RECT 2713.240 2152.725 2713.380 2391.910 ;
        RECT 2713.170 2152.355 2713.450 2152.725 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 1302.360 1690.150 1302.620 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 2713.170 2152.400 2713.450 2152.680 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT 2713.145 2152.690 2713.475 2152.705 ;
        RECT 2699.740 2152.640 2713.475 2152.690 ;
        RECT 2696.000 2152.390 2713.475 2152.640 ;
        RECT 2696.000 2152.040 2700.000 2152.390 ;
        RECT 2713.145 2152.375 2713.475 2152.390 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1300.950 2390.100 1301.270 2390.160 ;
        RECT 2716.370 2390.100 2716.690 2390.160 ;
        RECT 1300.950 2389.960 2716.690 2390.100 ;
        RECT 1300.950 2389.900 1301.270 2389.960 ;
        RECT 2716.370 2389.900 2716.690 2389.960 ;
        RECT 17.090 1476.520 17.410 1476.580 ;
        RECT 1300.950 1476.520 1301.270 1476.580 ;
        RECT 17.090 1476.380 1301.270 1476.520 ;
        RECT 17.090 1476.320 17.410 1476.380 ;
        RECT 1300.950 1476.320 1301.270 1476.380 ;
      LAYER via ;
        RECT 1300.980 2389.900 1301.240 2390.160 ;
        RECT 2716.400 2389.900 2716.660 2390.160 ;
        RECT 17.120 1476.320 17.380 1476.580 ;
        RECT 1300.980 1476.320 1301.240 1476.580 ;
      LAYER met2 ;
        RECT 1300.980 2389.870 1301.240 2390.190 ;
        RECT 2716.400 2389.870 2716.660 2390.190 ;
        RECT 1301.040 1476.610 1301.180 2389.870 ;
        RECT 2716.460 2184.005 2716.600 2389.870 ;
        RECT 2716.390 2183.635 2716.670 2184.005 ;
        RECT 17.120 1476.290 17.380 1476.610 ;
        RECT 1300.980 1476.290 1301.240 1476.610 ;
        RECT 17.180 1472.045 17.320 1476.290 ;
        RECT 17.110 1471.675 17.390 1472.045 ;
      LAYER via2 ;
        RECT 2716.390 2183.680 2716.670 2183.960 ;
        RECT 17.110 1471.720 17.390 1472.000 ;
      LAYER met3 ;
        RECT 2716.365 2183.970 2716.695 2183.985 ;
        RECT 2699.740 2183.920 2716.695 2183.970 ;
        RECT 2696.000 2183.670 2716.695 2183.920 ;
        RECT 2696.000 2183.320 2700.000 2183.670 ;
        RECT 2716.365 2183.655 2716.695 2183.670 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.085 1472.010 17.415 1472.025 ;
        RECT -4.800 1471.710 17.415 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.085 1471.695 17.415 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2697.530 2031.995 2697.810 2032.365 ;
        RECT 2697.600 2028.965 2697.740 2031.995 ;
        RECT 2697.530 2028.595 2697.810 2028.965 ;
        RECT 2697.530 2010.915 2697.810 2011.285 ;
        RECT 2697.600 1956.885 2697.740 2010.915 ;
        RECT 2697.530 1956.515 2697.810 1956.885 ;
        RECT 2697.530 1942.915 2697.810 1943.285 ;
        RECT 2697.600 1866.445 2697.740 1942.915 ;
        RECT 2697.530 1866.075 2697.810 1866.445 ;
        RECT 2696.610 1463.515 2696.890 1463.885 ;
        RECT 2696.680 1460.485 2696.820 1463.515 ;
        RECT 2696.610 1460.115 2696.890 1460.485 ;
        RECT 2696.610 1432.915 2696.890 1433.285 ;
        RECT 2696.680 1325.165 2696.820 1432.915 ;
        RECT 2696.610 1324.795 2696.890 1325.165 ;
        RECT 17.570 1256.115 17.850 1256.485 ;
        RECT 17.640 1204.125 17.780 1256.115 ;
        RECT 17.570 1203.755 17.850 1204.125 ;
      LAYER via2 ;
        RECT 2697.530 2032.040 2697.810 2032.320 ;
        RECT 2697.530 2028.640 2697.810 2028.920 ;
        RECT 2697.530 2010.960 2697.810 2011.240 ;
        RECT 2697.530 1956.560 2697.810 1956.840 ;
        RECT 2697.530 1942.960 2697.810 1943.240 ;
        RECT 2697.530 1866.120 2697.810 1866.400 ;
        RECT 2696.610 1463.560 2696.890 1463.840 ;
        RECT 2696.610 1460.160 2696.890 1460.440 ;
        RECT 2696.610 1432.960 2696.890 1433.240 ;
        RECT 2696.610 1324.840 2696.890 1325.120 ;
        RECT 17.570 1256.160 17.850 1256.440 ;
        RECT 17.570 1203.800 17.850 1204.080 ;
      LAYER met3 ;
        RECT 2696.000 2215.280 2700.000 2215.880 ;
        RECT 2696.830 2213.220 2697.130 2215.280 ;
        RECT 2696.790 2212.900 2697.170 2213.220 ;
        RECT 2697.505 2032.340 2697.835 2032.345 ;
        RECT 2697.505 2032.330 2698.090 2032.340 ;
        RECT 2697.280 2032.030 2698.090 2032.330 ;
        RECT 2697.505 2032.020 2698.090 2032.030 ;
        RECT 2697.505 2032.015 2697.835 2032.020 ;
        RECT 2696.790 2028.930 2697.170 2028.940 ;
        RECT 2697.505 2028.930 2697.835 2028.945 ;
        RECT 2696.790 2028.630 2697.835 2028.930 ;
        RECT 2696.790 2028.620 2697.170 2028.630 ;
        RECT 2697.505 2028.615 2697.835 2028.630 ;
        RECT 2696.790 2011.250 2697.170 2011.260 ;
        RECT 2697.505 2011.250 2697.835 2011.265 ;
        RECT 2696.790 2010.950 2697.835 2011.250 ;
        RECT 2696.790 2010.940 2697.170 2010.950 ;
        RECT 2697.505 2010.935 2697.835 2010.950 ;
        RECT 2696.790 1956.850 2697.170 1956.860 ;
        RECT 2697.505 1956.850 2697.835 1956.865 ;
        RECT 2696.790 1956.550 2697.835 1956.850 ;
        RECT 2696.790 1956.540 2697.170 1956.550 ;
        RECT 2697.505 1956.535 2697.835 1956.550 ;
        RECT 2696.790 1943.250 2697.170 1943.260 ;
        RECT 2697.505 1943.250 2697.835 1943.265 ;
        RECT 2696.790 1942.950 2697.835 1943.250 ;
        RECT 2696.790 1942.940 2697.170 1942.950 ;
        RECT 2697.505 1942.935 2697.835 1942.950 ;
        RECT 2697.505 1866.410 2697.835 1866.425 ;
        RECT 2698.630 1866.410 2699.010 1866.420 ;
        RECT 2697.505 1866.110 2699.010 1866.410 ;
        RECT 2697.505 1866.095 2697.835 1866.110 ;
        RECT 2698.630 1866.100 2699.010 1866.110 ;
        RECT 2696.790 1820.850 2697.170 1820.860 ;
        RECT 2698.630 1820.850 2699.010 1820.860 ;
        RECT 2696.790 1820.550 2699.010 1820.850 ;
        RECT 2696.790 1820.540 2697.170 1820.550 ;
        RECT 2698.630 1820.540 2699.010 1820.550 ;
        RECT 2696.585 1463.860 2696.915 1463.865 ;
        RECT 2696.585 1463.850 2697.170 1463.860 ;
        RECT 2696.360 1463.550 2697.170 1463.850 ;
        RECT 2696.585 1463.540 2697.170 1463.550 ;
        RECT 2696.585 1463.535 2696.915 1463.540 ;
        RECT 2696.585 1460.460 2696.915 1460.465 ;
        RECT 2696.585 1460.450 2697.170 1460.460 ;
        RECT 2696.585 1460.150 2697.370 1460.450 ;
        RECT 2696.585 1460.140 2697.170 1460.150 ;
        RECT 2696.585 1460.135 2696.915 1460.140 ;
        RECT 2696.585 1433.260 2696.915 1433.265 ;
        RECT 2696.585 1433.250 2697.170 1433.260 ;
        RECT 2696.585 1432.950 2697.370 1433.250 ;
        RECT 2696.585 1432.940 2697.170 1432.950 ;
        RECT 2696.585 1432.935 2696.915 1432.940 ;
        RECT 2696.585 1325.140 2696.915 1325.145 ;
        RECT 2696.585 1325.130 2697.170 1325.140 ;
        RECT 2696.360 1324.830 2697.170 1325.130 ;
        RECT 2696.585 1324.820 2697.170 1324.830 ;
        RECT 2696.585 1324.815 2696.915 1324.820 ;
        RECT 2696.790 1284.020 2697.170 1284.340 ;
        RECT 2696.830 1283.660 2697.130 1284.020 ;
        RECT 2696.790 1283.340 2697.170 1283.660 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 17.545 1256.450 17.875 1256.465 ;
        RECT -4.800 1256.150 17.875 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 17.545 1256.135 17.875 1256.150 ;
        RECT 17.545 1204.090 17.875 1204.105 ;
        RECT 2694.950 1204.090 2695.330 1204.100 ;
        RECT 17.545 1203.790 2695.330 1204.090 ;
        RECT 17.545 1203.775 17.875 1203.790 ;
        RECT 2694.950 1203.780 2695.330 1203.790 ;
      LAYER via3 ;
        RECT 2696.820 2212.900 2697.140 2213.220 ;
        RECT 2697.740 2032.020 2698.060 2032.340 ;
        RECT 2696.820 2028.620 2697.140 2028.940 ;
        RECT 2696.820 2010.940 2697.140 2011.260 ;
        RECT 2696.820 1956.540 2697.140 1956.860 ;
        RECT 2696.820 1942.940 2697.140 1943.260 ;
        RECT 2698.660 1866.100 2698.980 1866.420 ;
        RECT 2696.820 1820.540 2697.140 1820.860 ;
        RECT 2698.660 1820.540 2698.980 1820.860 ;
        RECT 2696.820 1463.540 2697.140 1463.860 ;
        RECT 2696.820 1460.140 2697.140 1460.460 ;
        RECT 2696.820 1432.940 2697.140 1433.260 ;
        RECT 2696.820 1324.820 2697.140 1325.140 ;
        RECT 2696.820 1284.020 2697.140 1284.340 ;
        RECT 2696.820 1283.340 2697.140 1283.660 ;
        RECT 2694.980 1203.780 2695.300 1204.100 ;
      LAYER met4 ;
        RECT 2696.815 2212.895 2697.145 2213.225 ;
        RECT 2696.830 2211.850 2697.130 2212.895 ;
        RECT 2694.990 2211.550 2697.130 2211.850 ;
        RECT 2694.990 2143.850 2695.290 2211.550 ;
        RECT 2694.990 2143.550 2696.210 2143.850 ;
        RECT 2695.910 2086.730 2696.210 2143.550 ;
        RECT 2695.910 2086.430 2698.050 2086.730 ;
        RECT 2697.750 2032.345 2698.050 2086.430 ;
        RECT 2697.735 2032.015 2698.065 2032.345 ;
        RECT 2696.815 2028.615 2697.145 2028.945 ;
        RECT 2696.830 2011.265 2697.130 2028.615 ;
        RECT 2696.815 2010.935 2697.145 2011.265 ;
        RECT 2696.815 1956.850 2697.145 1956.865 ;
        RECT 2695.910 1956.550 2697.145 1956.850 ;
        RECT 2695.910 1943.250 2696.210 1956.550 ;
        RECT 2696.815 1956.535 2697.145 1956.550 ;
        RECT 2696.815 1943.250 2697.145 1943.265 ;
        RECT 2695.910 1942.950 2697.145 1943.250 ;
        RECT 2696.815 1942.935 2697.145 1942.950 ;
        RECT 2698.655 1866.095 2698.985 1866.425 ;
        RECT 2698.670 1820.865 2698.970 1866.095 ;
        RECT 2696.815 1820.850 2697.145 1820.865 ;
        RECT 2695.910 1820.550 2697.145 1820.850 ;
        RECT 2695.910 1650.850 2696.210 1820.550 ;
        RECT 2696.815 1820.535 2697.145 1820.550 ;
        RECT 2698.655 1820.535 2698.985 1820.865 ;
        RECT 2694.990 1650.550 2696.210 1650.850 ;
        RECT 2694.990 1610.050 2695.290 1650.550 ;
        RECT 2694.990 1609.750 2696.210 1610.050 ;
        RECT 2695.910 1606.650 2696.210 1609.750 ;
        RECT 2694.070 1606.350 2696.210 1606.650 ;
        RECT 2694.070 1565.850 2694.370 1606.350 ;
        RECT 2694.070 1565.550 2695.290 1565.850 ;
        RECT 2694.990 1504.650 2695.290 1565.550 ;
        RECT 2694.070 1504.350 2695.290 1504.650 ;
        RECT 2694.070 1491.050 2694.370 1504.350 ;
        RECT 2694.070 1490.750 2696.210 1491.050 ;
        RECT 2695.910 1463.850 2696.210 1490.750 ;
        RECT 2696.815 1463.850 2697.145 1463.865 ;
        RECT 2695.910 1463.550 2697.145 1463.850 ;
        RECT 2696.815 1463.535 2697.145 1463.550 ;
        RECT 2696.815 1460.450 2697.145 1460.465 ;
        RECT 2694.990 1460.150 2697.145 1460.450 ;
        RECT 2694.990 1433.250 2695.290 1460.150 ;
        RECT 2696.815 1460.135 2697.145 1460.150 ;
        RECT 2696.815 1433.250 2697.145 1433.265 ;
        RECT 2694.990 1432.950 2697.145 1433.250 ;
        RECT 2696.815 1432.935 2697.145 1432.950 ;
        RECT 2696.815 1324.815 2697.145 1325.145 ;
        RECT 2696.830 1284.345 2697.130 1324.815 ;
        RECT 2696.815 1284.015 2697.145 1284.345 ;
        RECT 2696.815 1283.650 2697.145 1283.665 ;
        RECT 2695.910 1283.350 2697.145 1283.650 ;
        RECT 2695.910 1253.050 2696.210 1283.350 ;
        RECT 2696.815 1283.335 2697.145 1283.350 ;
        RECT 2694.990 1252.750 2696.210 1253.050 ;
        RECT 2694.990 1204.105 2695.290 1252.750 ;
        RECT 2694.975 1203.775 2695.305 1204.105 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 1041.660 17.410 1041.720 ;
        RECT 2708.090 1041.660 2708.410 1041.720 ;
        RECT 17.090 1041.520 2708.410 1041.660 ;
        RECT 17.090 1041.460 17.410 1041.520 ;
        RECT 2708.090 1041.460 2708.410 1041.520 ;
      LAYER via ;
        RECT 17.120 1041.460 17.380 1041.720 ;
        RECT 2708.120 1041.460 2708.380 1041.720 ;
      LAYER met2 ;
        RECT 2708.110 2246.875 2708.390 2247.245 ;
        RECT 2708.180 1041.750 2708.320 2246.875 ;
        RECT 17.120 1041.430 17.380 1041.750 ;
        RECT 2708.120 1041.430 2708.380 1041.750 ;
        RECT 17.180 1040.925 17.320 1041.430 ;
        RECT 17.110 1040.555 17.390 1040.925 ;
      LAYER via2 ;
        RECT 2708.110 2246.920 2708.390 2247.200 ;
        RECT 17.110 1040.600 17.390 1040.880 ;
      LAYER met3 ;
        RECT 2708.085 2247.210 2708.415 2247.225 ;
        RECT 2699.740 2247.160 2708.415 2247.210 ;
        RECT 2696.000 2246.910 2708.415 2247.160 ;
        RECT 2696.000 2246.560 2700.000 2246.910 ;
        RECT 2708.085 2246.895 2708.415 2246.910 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.085 1040.890 17.415 1040.905 ;
        RECT -4.800 1040.590 17.415 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.085 1040.575 17.415 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2703.050 1995.275 2703.330 1995.645 ;
        RECT 2703.120 1977.285 2703.260 1995.275 ;
        RECT 2703.050 1976.915 2703.330 1977.285 ;
        RECT 2691.550 1113.995 2691.830 1114.365 ;
        RECT 2691.620 1027.325 2691.760 1113.995 ;
        RECT 2691.550 1026.955 2691.830 1027.325 ;
        RECT 19.870 1005.195 20.150 1005.565 ;
        RECT 19.940 825.365 20.080 1005.195 ;
        RECT 19.870 824.995 20.150 825.365 ;
      LAYER via2 ;
        RECT 2703.050 1995.320 2703.330 1995.600 ;
        RECT 2703.050 1976.960 2703.330 1977.240 ;
        RECT 2691.550 1114.040 2691.830 1114.320 ;
        RECT 2691.550 1027.000 2691.830 1027.280 ;
        RECT 19.870 1005.240 20.150 1005.520 ;
        RECT 19.870 825.040 20.150 825.320 ;
      LAYER met3 ;
        RECT 2696.000 2278.520 2700.000 2279.120 ;
        RECT 2696.830 2276.460 2697.130 2278.520 ;
        RECT 2696.790 2276.140 2697.170 2276.460 ;
        RECT 2696.790 2256.050 2697.170 2256.060 ;
        RECT 2698.630 2256.050 2699.010 2256.060 ;
        RECT 2696.790 2255.750 2699.010 2256.050 ;
        RECT 2696.790 2255.740 2697.170 2255.750 ;
        RECT 2698.630 2255.740 2699.010 2255.750 ;
        RECT 2698.630 2212.530 2699.010 2212.540 ;
        RECT 2697.750 2212.230 2699.010 2212.530 ;
        RECT 2696.790 2211.170 2697.170 2211.180 ;
        RECT 2697.750 2211.170 2698.050 2212.230 ;
        RECT 2698.630 2212.220 2699.010 2212.230 ;
        RECT 2696.790 2210.870 2698.050 2211.170 ;
        RECT 2696.790 2210.860 2697.170 2210.870 ;
        RECT 2696.790 2072.450 2697.170 2072.460 ;
        RECT 2698.630 2072.450 2699.010 2072.460 ;
        RECT 2696.790 2072.150 2699.010 2072.450 ;
        RECT 2696.790 2072.140 2697.170 2072.150 ;
        RECT 2698.630 2072.140 2699.010 2072.150 ;
        RECT 2697.710 1995.610 2698.090 1995.620 ;
        RECT 2703.025 1995.610 2703.355 1995.625 ;
        RECT 2697.710 1995.310 2703.355 1995.610 ;
        RECT 2697.710 1995.300 2698.090 1995.310 ;
        RECT 2703.025 1995.295 2703.355 1995.310 ;
        RECT 2696.790 1977.250 2697.170 1977.260 ;
        RECT 2703.025 1977.250 2703.355 1977.265 ;
        RECT 2696.790 1976.950 2703.355 1977.250 ;
        RECT 2696.790 1976.940 2697.170 1976.950 ;
        RECT 2703.025 1976.935 2703.355 1976.950 ;
        RECT 2696.790 1942.570 2697.170 1942.580 ;
        RECT 2698.630 1942.570 2699.010 1942.580 ;
        RECT 2696.790 1942.270 2699.010 1942.570 ;
        RECT 2696.790 1942.260 2697.170 1942.270 ;
        RECT 2698.630 1942.260 2699.010 1942.270 ;
        RECT 2696.790 1917.410 2697.170 1917.420 ;
        RECT 2698.630 1917.410 2699.010 1917.420 ;
        RECT 2696.790 1917.110 2699.010 1917.410 ;
        RECT 2696.790 1917.100 2697.170 1917.110 ;
        RECT 2698.630 1917.100 2699.010 1917.110 ;
        RECT 2696.790 1882.050 2697.170 1882.060 ;
        RECT 2698.630 1882.050 2699.010 1882.060 ;
        RECT 2696.790 1881.750 2699.010 1882.050 ;
        RECT 2696.790 1881.740 2697.170 1881.750 ;
        RECT 2698.630 1881.740 2699.010 1881.750 ;
        RECT 2696.790 1873.210 2697.170 1873.220 ;
        RECT 2698.630 1873.210 2699.010 1873.220 ;
        RECT 2696.790 1872.910 2699.010 1873.210 ;
        RECT 2696.790 1872.900 2697.170 1872.910 ;
        RECT 2698.630 1872.900 2699.010 1872.910 ;
        RECT 2692.190 1138.810 2692.570 1138.820 ;
        RECT 2693.110 1138.810 2693.490 1138.820 ;
        RECT 2692.190 1138.510 2693.490 1138.810 ;
        RECT 2692.190 1138.500 2692.570 1138.510 ;
        RECT 2693.110 1138.500 2693.490 1138.510 ;
        RECT 2691.525 1114.330 2691.855 1114.345 ;
        RECT 2693.110 1114.330 2693.490 1114.340 ;
        RECT 2691.525 1114.030 2693.490 1114.330 ;
        RECT 2691.525 1114.015 2691.855 1114.030 ;
        RECT 2693.110 1114.020 2693.490 1114.030 ;
        RECT 2691.525 1027.300 2691.855 1027.305 ;
        RECT 2691.270 1027.290 2691.855 1027.300 ;
        RECT 2691.070 1026.990 2691.855 1027.290 ;
        RECT 2691.270 1026.980 2691.855 1026.990 ;
        RECT 2691.525 1026.975 2691.855 1026.980 ;
        RECT 19.845 1005.530 20.175 1005.545 ;
        RECT 2691.270 1005.530 2691.650 1005.540 ;
        RECT 19.845 1005.230 2691.650 1005.530 ;
        RECT 19.845 1005.215 20.175 1005.230 ;
        RECT 2691.270 1005.220 2691.650 1005.230 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 19.845 825.330 20.175 825.345 ;
        RECT -4.800 825.030 20.175 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 19.845 825.015 20.175 825.030 ;
      LAYER via3 ;
        RECT 2696.820 2276.140 2697.140 2276.460 ;
        RECT 2696.820 2255.740 2697.140 2256.060 ;
        RECT 2698.660 2255.740 2698.980 2256.060 ;
        RECT 2696.820 2210.860 2697.140 2211.180 ;
        RECT 2698.660 2212.220 2698.980 2212.540 ;
        RECT 2696.820 2072.140 2697.140 2072.460 ;
        RECT 2698.660 2072.140 2698.980 2072.460 ;
        RECT 2697.740 1995.300 2698.060 1995.620 ;
        RECT 2696.820 1976.940 2697.140 1977.260 ;
        RECT 2696.820 1942.260 2697.140 1942.580 ;
        RECT 2698.660 1942.260 2698.980 1942.580 ;
        RECT 2696.820 1917.100 2697.140 1917.420 ;
        RECT 2698.660 1917.100 2698.980 1917.420 ;
        RECT 2696.820 1881.740 2697.140 1882.060 ;
        RECT 2698.660 1881.740 2698.980 1882.060 ;
        RECT 2696.820 1872.900 2697.140 1873.220 ;
        RECT 2698.660 1872.900 2698.980 1873.220 ;
        RECT 2692.220 1138.500 2692.540 1138.820 ;
        RECT 2693.140 1138.500 2693.460 1138.820 ;
        RECT 2693.140 1114.020 2693.460 1114.340 ;
        RECT 2691.300 1026.980 2691.620 1027.300 ;
        RECT 2691.300 1005.220 2691.620 1005.540 ;
      LAYER met4 ;
        RECT 2696.815 2276.450 2697.145 2276.465 ;
        RECT 2695.910 2276.150 2697.145 2276.450 ;
        RECT 2695.910 2256.050 2696.210 2276.150 ;
        RECT 2696.815 2276.135 2697.145 2276.150 ;
        RECT 2696.815 2256.050 2697.145 2256.065 ;
        RECT 2695.910 2255.750 2697.145 2256.050 ;
        RECT 2696.815 2255.735 2697.145 2255.750 ;
        RECT 2698.655 2255.735 2698.985 2256.065 ;
        RECT 2698.670 2212.545 2698.970 2255.735 ;
        RECT 2698.655 2212.215 2698.985 2212.545 ;
        RECT 2696.815 2210.855 2697.145 2211.185 ;
        RECT 2696.830 2089.450 2697.130 2210.855 ;
        RECT 2696.830 2089.150 2698.970 2089.450 ;
        RECT 2698.670 2072.465 2698.970 2089.150 ;
        RECT 2696.815 2072.450 2697.145 2072.465 ;
        RECT 2693.150 2072.150 2697.145 2072.450 ;
        RECT 2693.150 2007.850 2693.450 2072.150 ;
        RECT 2696.815 2072.135 2697.145 2072.150 ;
        RECT 2698.655 2072.135 2698.985 2072.465 ;
        RECT 2693.150 2007.550 2694.370 2007.850 ;
        RECT 2694.070 1994.250 2694.370 2007.550 ;
        RECT 2697.735 1995.295 2698.065 1995.625 ;
        RECT 2697.750 1994.250 2698.050 1995.295 ;
        RECT 2694.070 1993.950 2698.050 1994.250 ;
        RECT 2696.815 1977.250 2697.145 1977.265 ;
        RECT 2694.070 1976.950 2697.145 1977.250 ;
        RECT 2694.070 1942.570 2694.370 1976.950 ;
        RECT 2696.815 1976.935 2697.145 1976.950 ;
        RECT 2696.815 1942.570 2697.145 1942.585 ;
        RECT 2694.070 1942.270 2697.145 1942.570 ;
        RECT 2696.815 1942.255 2697.145 1942.270 ;
        RECT 2698.655 1942.255 2698.985 1942.585 ;
        RECT 2698.670 1917.425 2698.970 1942.255 ;
        RECT 2696.815 1917.095 2697.145 1917.425 ;
        RECT 2698.655 1917.095 2698.985 1917.425 ;
        RECT 2696.830 1882.065 2697.130 1917.095 ;
        RECT 2696.815 1881.735 2697.145 1882.065 ;
        RECT 2698.655 1881.735 2698.985 1882.065 ;
        RECT 2698.670 1873.225 2698.970 1881.735 ;
        RECT 2696.815 1872.895 2697.145 1873.225 ;
        RECT 2698.655 1872.895 2698.985 1873.225 ;
        RECT 2696.830 1861.650 2697.130 1872.895 ;
        RECT 2694.070 1861.350 2697.130 1861.650 ;
        RECT 2694.070 1848.730 2694.370 1861.350 ;
        RECT 2693.150 1848.430 2694.370 1848.730 ;
        RECT 2693.150 1763.050 2693.450 1848.430 ;
        RECT 2693.150 1762.750 2694.370 1763.050 ;
        RECT 2694.070 1712.050 2694.370 1762.750 ;
        RECT 2692.230 1711.750 2694.370 1712.050 ;
        RECT 2692.230 1708.650 2692.530 1711.750 ;
        RECT 2691.310 1708.350 2692.530 1708.650 ;
        RECT 2691.310 1637.250 2691.610 1708.350 ;
        RECT 2691.310 1636.950 2693.450 1637.250 ;
        RECT 2693.150 1613.450 2693.450 1636.950 ;
        RECT 2691.310 1613.150 2693.450 1613.450 ;
        RECT 2691.310 1606.650 2691.610 1613.150 ;
        RECT 2691.310 1606.350 2692.530 1606.650 ;
        RECT 2692.230 1586.930 2692.530 1606.350 ;
        RECT 2690.390 1586.630 2692.530 1586.930 ;
        RECT 2690.390 1501.250 2690.690 1586.630 ;
        RECT 2689.470 1500.950 2690.690 1501.250 ;
        RECT 2689.470 1457.050 2689.770 1500.950 ;
        RECT 2689.470 1456.750 2691.610 1457.050 ;
        RECT 2691.310 1409.450 2691.610 1456.750 ;
        RECT 2691.310 1409.150 2694.370 1409.450 ;
        RECT 2694.070 1327.850 2694.370 1409.150 ;
        RECT 2694.070 1327.550 2695.290 1327.850 ;
        RECT 2694.990 1283.650 2695.290 1327.550 ;
        RECT 2694.070 1283.350 2695.290 1283.650 ;
        RECT 2694.070 1273.450 2694.370 1283.350 ;
        RECT 2694.070 1273.150 2695.290 1273.450 ;
        RECT 2694.990 1256.450 2695.290 1273.150 ;
        RECT 2692.230 1256.150 2695.290 1256.450 ;
        RECT 2692.230 1232.650 2692.530 1256.150 ;
        RECT 2692.230 1232.350 2694.370 1232.650 ;
        RECT 2694.070 1212.250 2694.370 1232.350 ;
        RECT 2692.230 1211.950 2694.370 1212.250 ;
        RECT 2692.230 1138.825 2692.530 1211.950 ;
        RECT 2692.215 1138.495 2692.545 1138.825 ;
        RECT 2693.135 1138.495 2693.465 1138.825 ;
        RECT 2693.150 1114.345 2693.450 1138.495 ;
        RECT 2693.135 1114.015 2693.465 1114.345 ;
        RECT 2691.295 1026.975 2691.625 1027.305 ;
        RECT 2691.310 1005.545 2691.610 1026.975 ;
        RECT 2691.295 1005.215 2691.625 1005.545 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 1004.515 17.390 1004.885 ;
        RECT 17.180 610.485 17.320 1004.515 ;
        RECT 17.110 610.115 17.390 610.485 ;
      LAYER via2 ;
        RECT 17.110 1004.560 17.390 1004.840 ;
        RECT 17.110 610.160 17.390 610.440 ;
      LAYER met3 ;
        RECT 2701.390 2310.450 2701.770 2310.460 ;
        RECT 2699.740 2310.400 2701.770 2310.450 ;
        RECT 2696.000 2310.150 2701.770 2310.400 ;
        RECT 2696.000 2309.800 2700.000 2310.150 ;
        RECT 2701.390 2310.140 2701.770 2310.150 ;
        RECT 17.085 1004.850 17.415 1004.865 ;
        RECT 2701.390 1004.850 2701.770 1004.860 ;
        RECT 17.085 1004.550 2701.770 1004.850 ;
        RECT 17.085 1004.535 17.415 1004.550 ;
        RECT 2701.390 1004.540 2701.770 1004.550 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 17.085 610.450 17.415 610.465 ;
        RECT -4.800 610.150 17.415 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 17.085 610.135 17.415 610.150 ;
      LAYER via3 ;
        RECT 2701.420 2310.140 2701.740 2310.460 ;
        RECT 2701.420 1004.540 2701.740 1004.860 ;
      LAYER met4 ;
        RECT 2701.415 2310.135 2701.745 2310.465 ;
        RECT 2701.430 1004.865 2701.730 2310.135 ;
        RECT 2701.415 1004.535 2701.745 1004.865 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.110 399.995 17.390 400.365 ;
        RECT 17.180 394.925 17.320 399.995 ;
        RECT 17.110 394.555 17.390 394.925 ;
      LAYER via2 ;
        RECT 17.110 400.040 17.390 400.320 ;
        RECT 17.110 394.600 17.390 394.880 ;
      LAYER met3 ;
        RECT 2714.270 2342.410 2714.650 2342.420 ;
        RECT 2699.740 2342.360 2714.650 2342.410 ;
        RECT 2696.000 2342.110 2714.650 2342.360 ;
        RECT 2696.000 2341.760 2700.000 2342.110 ;
        RECT 2714.270 2342.100 2714.650 2342.110 ;
        RECT 17.085 400.330 17.415 400.345 ;
        RECT 2714.270 400.330 2714.650 400.340 ;
        RECT 17.085 400.030 2714.650 400.330 ;
        RECT 17.085 400.015 17.415 400.030 ;
        RECT 2714.270 400.020 2714.650 400.030 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 17.085 394.890 17.415 394.905 ;
        RECT -4.800 394.590 17.415 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 17.085 394.575 17.415 394.590 ;
      LAYER via3 ;
        RECT 2714.300 2342.100 2714.620 2342.420 ;
        RECT 2714.300 400.020 2714.620 400.340 ;
      LAYER met4 ;
        RECT 2714.295 2342.095 2714.625 2342.425 ;
        RECT 2714.310 400.345 2714.610 2342.095 ;
        RECT 2714.295 400.015 2714.625 400.345 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2713.350 2373.690 2713.730 2373.700 ;
        RECT 2699.740 2373.640 2713.730 2373.690 ;
        RECT 2696.000 2373.390 2713.730 2373.640 ;
        RECT 2696.000 2373.040 2700.000 2373.390 ;
        RECT 2713.350 2373.380 2713.730 2373.390 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 2713.350 179.330 2713.730 179.340 ;
        RECT -4.800 179.030 2713.730 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 2713.350 179.020 2713.730 179.030 ;
      LAYER via3 ;
        RECT 2713.380 2373.380 2713.700 2373.700 ;
        RECT 2713.380 179.020 2713.700 179.340 ;
      LAYER met4 ;
        RECT 2713.375 2373.375 2713.705 2373.705 ;
        RECT 2713.390 179.345 2713.690 2373.375 ;
        RECT 2713.375 179.015 2713.705 179.345 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2715.910 793.460 2716.230 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 2715.910 793.320 2899.310 793.460 ;
        RECT 2715.910 793.260 2716.230 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 2715.940 793.260 2716.200 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 2715.470 1299.635 2715.750 1300.005 ;
        RECT 2715.540 1258.410 2715.680 1299.635 ;
        RECT 2715.540 1258.270 2716.140 1258.410 ;
        RECT 2716.000 793.550 2716.140 1258.270 ;
        RECT 2715.940 793.230 2716.200 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2715.470 1299.680 2715.750 1299.960 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2715.445 1299.970 2715.775 1299.985 ;
        RECT 2699.740 1299.920 2715.775 1299.970 ;
        RECT 2696.000 1299.670 2715.775 1299.920 ;
        RECT 2696.000 1299.320 2700.000 1299.670 ;
        RECT 2715.445 1299.655 2715.775 1299.670 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2716.830 1028.060 2717.150 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 2716.830 1027.920 2899.310 1028.060 ;
        RECT 2716.830 1027.860 2717.150 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 2716.860 1027.860 2717.120 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 2716.850 1330.915 2717.130 1331.285 ;
        RECT 2716.920 1028.150 2717.060 1330.915 ;
        RECT 2716.860 1027.830 2717.120 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2716.850 1330.960 2717.130 1331.240 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2716.825 1331.250 2717.155 1331.265 ;
        RECT 2699.740 1331.200 2717.155 1331.250 ;
        RECT 2696.000 1330.950 2717.155 1331.200 ;
        RECT 2696.000 1330.600 2700.000 1330.950 ;
        RECT 2716.825 1330.935 2717.155 1330.950 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2714.990 1262.660 2715.310 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 2714.990 1262.520 2899.310 1262.660 ;
        RECT 2714.990 1262.460 2715.310 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 2715.020 1262.460 2715.280 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 2715.010 1362.875 2715.290 1363.245 ;
        RECT 2715.080 1262.750 2715.220 1362.875 ;
        RECT 2715.020 1262.430 2715.280 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2715.010 1362.920 2715.290 1363.200 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2714.985 1363.210 2715.315 1363.225 ;
        RECT 2699.740 1363.160 2715.315 1363.210 ;
        RECT 2696.000 1362.910 2715.315 1363.160 ;
        RECT 2696.000 1362.560 2700.000 1362.910 ;
        RECT 2714.985 1362.895 2715.315 1362.910 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2705.790 1400.700 2706.110 1400.760 ;
        RECT 2903.590 1400.700 2903.910 1400.760 ;
        RECT 2705.790 1400.560 2903.910 1400.700 ;
        RECT 2705.790 1400.500 2706.110 1400.560 ;
        RECT 2903.590 1400.500 2903.910 1400.560 ;
      LAYER via ;
        RECT 2705.820 1400.500 2706.080 1400.760 ;
        RECT 2903.620 1400.500 2903.880 1400.760 ;
      LAYER met2 ;
        RECT 2903.610 1495.475 2903.890 1495.845 ;
        RECT 2903.680 1400.790 2903.820 1495.475 ;
        RECT 2705.820 1400.470 2706.080 1400.790 ;
        RECT 2903.620 1400.470 2903.880 1400.790 ;
        RECT 2705.880 1397.245 2706.020 1400.470 ;
        RECT 2705.810 1396.875 2706.090 1397.245 ;
      LAYER via2 ;
        RECT 2903.610 1495.520 2903.890 1495.800 ;
        RECT 2705.810 1396.920 2706.090 1397.200 ;
      LAYER met3 ;
        RECT 2903.585 1495.810 2903.915 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2903.585 1495.510 2924.800 1495.810 ;
        RECT 2903.585 1495.495 2903.915 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
        RECT 2705.785 1397.210 2706.115 1397.225 ;
        RECT 2698.670 1396.910 2706.115 1397.210 ;
        RECT 2698.670 1394.440 2698.970 1396.910 ;
        RECT 2705.785 1396.895 2706.115 1396.910 ;
        RECT 2696.000 1393.840 2700.000 1394.440 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1428.240 2713.470 1428.300 ;
        RECT 2902.210 1428.240 2902.530 1428.300 ;
        RECT 2713.150 1428.100 2902.530 1428.240 ;
        RECT 2713.150 1428.040 2713.470 1428.100 ;
        RECT 2902.210 1428.040 2902.530 1428.100 ;
      LAYER via ;
        RECT 2713.180 1428.040 2713.440 1428.300 ;
        RECT 2902.240 1428.040 2902.500 1428.300 ;
      LAYER met2 ;
        RECT 2902.230 1730.075 2902.510 1730.445 ;
        RECT 2902.300 1428.330 2902.440 1730.075 ;
        RECT 2713.180 1428.010 2713.440 1428.330 ;
        RECT 2902.240 1428.010 2902.500 1428.330 ;
        RECT 2713.240 1426.485 2713.380 1428.010 ;
        RECT 2713.170 1426.115 2713.450 1426.485 ;
      LAYER via2 ;
        RECT 2902.230 1730.120 2902.510 1730.400 ;
        RECT 2713.170 1426.160 2713.450 1426.440 ;
      LAYER met3 ;
        RECT 2902.205 1730.410 2902.535 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2902.205 1730.110 2924.800 1730.410 ;
        RECT 2902.205 1730.095 2902.535 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
        RECT 2713.145 1426.450 2713.475 1426.465 ;
        RECT 2699.740 1426.400 2713.475 1426.450 ;
        RECT 2696.000 1426.150 2713.475 1426.400 ;
        RECT 2696.000 1425.800 2700.000 1426.150 ;
        RECT 2713.145 1426.135 2713.475 1426.150 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2723.270 1960.000 2723.590 1960.060 ;
        RECT 2900.830 1960.000 2901.150 1960.060 ;
        RECT 2723.270 1959.860 2901.150 1960.000 ;
        RECT 2723.270 1959.800 2723.590 1959.860 ;
        RECT 2900.830 1959.800 2901.150 1959.860 ;
        RECT 2713.150 1456.460 2713.470 1456.520 ;
        RECT 2723.270 1456.460 2723.590 1456.520 ;
        RECT 2713.150 1456.320 2723.590 1456.460 ;
        RECT 2713.150 1456.260 2713.470 1456.320 ;
        RECT 2723.270 1456.260 2723.590 1456.320 ;
      LAYER via ;
        RECT 2723.300 1959.800 2723.560 1960.060 ;
        RECT 2900.860 1959.800 2901.120 1960.060 ;
        RECT 2713.180 1456.260 2713.440 1456.520 ;
        RECT 2723.300 1456.260 2723.560 1456.520 ;
      LAYER met2 ;
        RECT 2900.850 1964.675 2901.130 1965.045 ;
        RECT 2900.920 1960.090 2901.060 1964.675 ;
        RECT 2723.300 1959.770 2723.560 1960.090 ;
        RECT 2900.860 1959.770 2901.120 1960.090 ;
        RECT 2713.170 1457.395 2713.450 1457.765 ;
        RECT 2713.240 1456.550 2713.380 1457.395 ;
        RECT 2723.360 1456.550 2723.500 1959.770 ;
        RECT 2713.180 1456.230 2713.440 1456.550 ;
        RECT 2723.300 1456.230 2723.560 1456.550 ;
      LAYER via2 ;
        RECT 2900.850 1964.720 2901.130 1965.000 ;
        RECT 2713.170 1457.440 2713.450 1457.720 ;
      LAYER met3 ;
        RECT 2900.825 1965.010 2901.155 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2900.825 1964.710 2924.800 1965.010 ;
        RECT 2900.825 1964.695 2901.155 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
        RECT 2713.145 1457.730 2713.475 1457.745 ;
        RECT 2699.740 1457.680 2713.475 1457.730 ;
        RECT 2696.000 1457.430 2713.475 1457.680 ;
        RECT 2696.000 1457.080 2700.000 1457.430 ;
        RECT 2713.145 1457.415 2713.475 1457.430 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2770.650 2194.600 2770.970 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 2770.650 2194.460 2901.150 2194.600 ;
        RECT 2770.650 2194.400 2770.970 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 2713.150 1490.460 2713.470 1490.520 ;
        RECT 2770.650 1490.460 2770.970 1490.520 ;
        RECT 2713.150 1490.320 2770.970 1490.460 ;
        RECT 2713.150 1490.260 2713.470 1490.320 ;
        RECT 2770.650 1490.260 2770.970 1490.320 ;
      LAYER via ;
        RECT 2770.680 2194.400 2770.940 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 2713.180 1490.260 2713.440 1490.520 ;
        RECT 2770.680 1490.260 2770.940 1490.520 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 2770.680 2194.370 2770.940 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 2770.740 1490.550 2770.880 2194.370 ;
        RECT 2713.180 1490.230 2713.440 1490.550 ;
        RECT 2770.680 1490.230 2770.940 1490.550 ;
        RECT 2713.240 1489.725 2713.380 1490.230 ;
        RECT 2713.170 1489.355 2713.450 1489.725 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
        RECT 2713.170 1489.400 2713.450 1489.680 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
        RECT 2713.145 1489.690 2713.475 1489.705 ;
        RECT 2699.740 1489.640 2713.475 1489.690 ;
        RECT 2696.000 1489.390 2713.475 1489.640 ;
        RECT 2696.000 1489.040 2700.000 1489.390 ;
        RECT 2713.145 1489.375 2713.475 1489.390 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2712.230 1214.720 2712.550 1214.780 ;
        RECT 2770.190 1214.720 2770.510 1214.780 ;
        RECT 2712.230 1214.580 2770.510 1214.720 ;
        RECT 2712.230 1214.520 2712.550 1214.580 ;
        RECT 2770.190 1214.520 2770.510 1214.580 ;
        RECT 2770.190 206.960 2770.510 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 2770.190 206.820 2901.150 206.960 ;
        RECT 2770.190 206.760 2770.510 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 2712.260 1214.520 2712.520 1214.780 ;
        RECT 2770.220 1214.520 2770.480 1214.780 ;
        RECT 2770.220 206.760 2770.480 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 2712.250 1215.315 2712.530 1215.685 ;
        RECT 2712.320 1214.810 2712.460 1215.315 ;
        RECT 2712.260 1214.490 2712.520 1214.810 ;
        RECT 2770.220 1214.490 2770.480 1214.810 ;
        RECT 2770.280 207.050 2770.420 1214.490 ;
        RECT 2770.220 206.730 2770.480 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2712.250 1215.360 2712.530 1215.640 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2712.225 1215.650 2712.555 1215.665 ;
        RECT 2699.740 1215.600 2712.555 1215.650 ;
        RECT 2696.000 1215.350 2712.555 1215.600 ;
        RECT 2696.000 1215.000 2700.000 1215.350 ;
        RECT 2712.225 1215.335 2712.555 1215.350 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2777.090 2546.500 2777.410 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 2777.090 2546.360 2901.150 2546.500 ;
        RECT 2777.090 2546.300 2777.410 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
        RECT 2713.150 1531.600 2713.470 1531.660 ;
        RECT 2777.090 1531.600 2777.410 1531.660 ;
        RECT 2713.150 1531.460 2777.410 1531.600 ;
        RECT 2713.150 1531.400 2713.470 1531.460 ;
        RECT 2777.090 1531.400 2777.410 1531.460 ;
      LAYER via ;
        RECT 2777.120 2546.300 2777.380 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
        RECT 2713.180 1531.400 2713.440 1531.660 ;
        RECT 2777.120 1531.400 2777.380 1531.660 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 2777.120 2546.270 2777.380 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 2777.180 1531.690 2777.320 2546.270 ;
        RECT 2713.180 1531.370 2713.440 1531.690 ;
        RECT 2777.120 1531.370 2777.380 1531.690 ;
        RECT 2713.240 1531.205 2713.380 1531.370 ;
        RECT 2713.170 1530.835 2713.450 1531.205 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
        RECT 2713.170 1530.880 2713.450 1531.160 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
        RECT 2713.145 1531.170 2713.475 1531.185 ;
        RECT 2699.740 1531.120 2713.475 1531.170 ;
        RECT 2696.000 1530.870 2713.475 1531.120 ;
        RECT 2696.000 1530.520 2700.000 1530.870 ;
        RECT 2713.145 1530.855 2713.475 1530.870 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2783.990 2781.100 2784.310 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 2783.990 2780.960 2901.150 2781.100 ;
        RECT 2783.990 2780.900 2784.310 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
        RECT 2713.150 1566.280 2713.470 1566.340 ;
        RECT 2783.990 1566.280 2784.310 1566.340 ;
        RECT 2713.150 1566.140 2784.310 1566.280 ;
        RECT 2713.150 1566.080 2713.470 1566.140 ;
        RECT 2783.990 1566.080 2784.310 1566.140 ;
      LAYER via ;
        RECT 2784.020 2780.900 2784.280 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
        RECT 2713.180 1566.080 2713.440 1566.340 ;
        RECT 2784.020 1566.080 2784.280 1566.340 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 2784.020 2780.870 2784.280 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 2784.080 1566.370 2784.220 2780.870 ;
        RECT 2713.180 1566.050 2713.440 1566.370 ;
        RECT 2784.020 1566.050 2784.280 1566.370 ;
        RECT 2713.240 1563.165 2713.380 1566.050 ;
        RECT 2713.170 1562.795 2713.450 1563.165 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
        RECT 2713.170 1562.840 2713.450 1563.120 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
        RECT 2713.145 1563.130 2713.475 1563.145 ;
        RECT 2699.740 1563.080 2713.475 1563.130 ;
        RECT 2696.000 1562.830 2713.475 1563.080 ;
        RECT 2696.000 1562.480 2700.000 1562.830 ;
        RECT 2713.145 1562.815 2713.475 1562.830 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2790.890 3015.700 2791.210 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 2790.890 3015.560 2901.150 3015.700 ;
        RECT 2790.890 3015.500 2791.210 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
        RECT 2713.150 1600.620 2713.470 1600.680 ;
        RECT 2790.890 1600.620 2791.210 1600.680 ;
        RECT 2713.150 1600.480 2791.210 1600.620 ;
        RECT 2713.150 1600.420 2713.470 1600.480 ;
        RECT 2790.890 1600.420 2791.210 1600.480 ;
      LAYER via ;
        RECT 2790.920 3015.500 2791.180 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
        RECT 2713.180 1600.420 2713.440 1600.680 ;
        RECT 2790.920 1600.420 2791.180 1600.680 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 2790.920 3015.470 2791.180 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 2790.980 1600.710 2791.120 3015.470 ;
        RECT 2713.180 1600.390 2713.440 1600.710 ;
        RECT 2790.920 1600.390 2791.180 1600.710 ;
        RECT 2713.240 1594.445 2713.380 1600.390 ;
        RECT 2713.170 1594.075 2713.450 1594.445 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
        RECT 2713.170 1594.120 2713.450 1594.400 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
        RECT 2713.145 1594.410 2713.475 1594.425 ;
        RECT 2699.740 1594.360 2713.475 1594.410 ;
        RECT 2696.000 1594.110 2713.475 1594.360 ;
        RECT 2696.000 1593.760 2700.000 1594.110 ;
        RECT 2713.145 1594.095 2713.475 1594.110 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2804.690 3250.300 2805.010 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 2804.690 3250.160 2901.150 3250.300 ;
        RECT 2804.690 3250.100 2805.010 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 2713.150 1628.160 2713.470 1628.220 ;
        RECT 2804.690 1628.160 2805.010 1628.220 ;
        RECT 2713.150 1628.020 2805.010 1628.160 ;
        RECT 2713.150 1627.960 2713.470 1628.020 ;
        RECT 2804.690 1627.960 2805.010 1628.020 ;
      LAYER via ;
        RECT 2804.720 3250.100 2804.980 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 2713.180 1627.960 2713.440 1628.220 ;
        RECT 2804.720 1627.960 2804.980 1628.220 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 2804.720 3250.070 2804.980 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 2804.780 1628.250 2804.920 3250.070 ;
        RECT 2713.180 1627.930 2713.440 1628.250 ;
        RECT 2804.720 1627.930 2804.980 1628.250 ;
        RECT 2713.240 1626.405 2713.380 1627.930 ;
        RECT 2713.170 1626.035 2713.450 1626.405 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
        RECT 2713.170 1626.080 2713.450 1626.360 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
        RECT 2713.145 1626.370 2713.475 1626.385 ;
        RECT 2699.740 1626.320 2713.475 1626.370 ;
        RECT 2696.000 1626.070 2713.475 1626.320 ;
        RECT 2696.000 1625.720 2700.000 1626.070 ;
        RECT 2713.145 1626.055 2713.475 1626.070 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2818.490 3484.900 2818.810 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 2818.490 3484.760 2901.150 3484.900 ;
        RECT 2818.490 3484.700 2818.810 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 2713.150 1662.840 2713.470 1662.900 ;
        RECT 2818.490 1662.840 2818.810 1662.900 ;
        RECT 2713.150 1662.700 2818.810 1662.840 ;
        RECT 2713.150 1662.640 2713.470 1662.700 ;
        RECT 2818.490 1662.640 2818.810 1662.700 ;
      LAYER via ;
        RECT 2818.520 3484.700 2818.780 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 2713.180 1662.640 2713.440 1662.900 ;
        RECT 2818.520 1662.640 2818.780 1662.900 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 2818.520 3484.670 2818.780 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 2818.580 1662.930 2818.720 3484.670 ;
        RECT 2713.180 1662.610 2713.440 1662.930 ;
        RECT 2818.520 1662.610 2818.780 1662.930 ;
        RECT 2713.240 1657.685 2713.380 1662.610 ;
        RECT 2713.170 1657.315 2713.450 1657.685 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
        RECT 2713.170 1657.360 2713.450 1657.640 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
        RECT 2713.145 1657.650 2713.475 1657.665 ;
        RECT 2699.740 1657.600 2713.475 1657.650 ;
        RECT 2696.000 1657.350 2713.475 1657.600 ;
        RECT 2696.000 1657.000 2700.000 1657.350 ;
        RECT 2713.145 1657.335 2713.475 1657.350 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2635.870 3498.500 2636.190 3498.560 ;
        RECT 2642.310 3498.500 2642.630 3498.560 ;
        RECT 2635.870 3498.360 2642.630 3498.500 ;
        RECT 2635.870 3498.300 2636.190 3498.360 ;
        RECT 2642.310 3498.300 2642.630 3498.360 ;
        RECT 2642.310 2399.280 2642.630 2399.340 ;
        RECT 2709.010 2399.280 2709.330 2399.340 ;
        RECT 2642.310 2399.140 2709.330 2399.280 ;
        RECT 2642.310 2399.080 2642.630 2399.140 ;
        RECT 2709.010 2399.080 2709.330 2399.140 ;
      LAYER via ;
        RECT 2635.900 3498.300 2636.160 3498.560 ;
        RECT 2642.340 3498.300 2642.600 3498.560 ;
        RECT 2642.340 2399.080 2642.600 2399.340 ;
        RECT 2709.040 2399.080 2709.300 2399.340 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3498.590 2636.100 3517.600 ;
        RECT 2635.900 3498.270 2636.160 3498.590 ;
        RECT 2642.340 3498.270 2642.600 3498.590 ;
        RECT 2642.400 2399.370 2642.540 3498.270 ;
        RECT 2642.340 2399.050 2642.600 2399.370 ;
        RECT 2709.040 2399.050 2709.300 2399.370 ;
        RECT 2709.100 1689.645 2709.240 2399.050 ;
        RECT 2709.030 1689.275 2709.310 1689.645 ;
      LAYER via2 ;
        RECT 2709.030 1689.320 2709.310 1689.600 ;
      LAYER met3 ;
        RECT 2709.005 1689.610 2709.335 1689.625 ;
        RECT 2699.740 1689.560 2709.335 1689.610 ;
        RECT 2696.000 1689.310 2709.335 1689.560 ;
        RECT 2696.000 1688.960 2700.000 1689.310 ;
        RECT 2709.005 1689.295 2709.335 1689.310 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2311.570 3498.500 2311.890 3498.560 ;
        RECT 2318.010 3498.500 2318.330 3498.560 ;
        RECT 2311.570 3498.360 2318.330 3498.500 ;
        RECT 2311.570 3498.300 2311.890 3498.360 ;
        RECT 2318.010 3498.300 2318.330 3498.360 ;
        RECT 2318.010 3053.780 2318.330 3053.840 ;
        RECT 2696.590 3053.780 2696.910 3053.840 ;
        RECT 2318.010 3053.640 2696.910 3053.780 ;
        RECT 2318.010 3053.580 2318.330 3053.640 ;
        RECT 2696.590 3053.580 2696.910 3053.640 ;
        RECT 2696.590 1787.080 2696.910 1787.340 ;
        RECT 2696.680 1786.320 2696.820 1787.080 ;
        RECT 2696.590 1786.060 2696.910 1786.320 ;
      LAYER via ;
        RECT 2311.600 3498.300 2311.860 3498.560 ;
        RECT 2318.040 3498.300 2318.300 3498.560 ;
        RECT 2318.040 3053.580 2318.300 3053.840 ;
        RECT 2696.620 3053.580 2696.880 3053.840 ;
        RECT 2696.620 1787.080 2696.880 1787.340 ;
        RECT 2696.620 1786.060 2696.880 1786.320 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3498.590 2311.800 3517.600 ;
        RECT 2311.600 3498.270 2311.860 3498.590 ;
        RECT 2318.040 3498.270 2318.300 3498.590 ;
        RECT 2318.100 3053.870 2318.240 3498.270 ;
        RECT 2318.040 3053.550 2318.300 3053.870 ;
        RECT 2696.620 3053.550 2696.880 3053.870 ;
        RECT 2696.680 1787.370 2696.820 3053.550 ;
        RECT 2696.620 1787.050 2696.880 1787.370 ;
        RECT 2696.620 1786.030 2696.880 1786.350 ;
        RECT 2696.680 1721.605 2696.820 1786.030 ;
        RECT 2696.610 1721.235 2696.890 1721.605 ;
      LAYER via2 ;
        RECT 2696.610 1721.280 2696.890 1721.560 ;
      LAYER met3 ;
        RECT 2696.585 1721.570 2696.915 1721.585 ;
        RECT 2696.585 1721.255 2697.130 1721.570 ;
        RECT 2696.830 1720.840 2697.130 1721.255 ;
        RECT 2696.000 1720.240 2700.000 1720.840 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1987.270 3499.860 1987.590 3499.920 ;
        RECT 1993.710 3499.860 1994.030 3499.920 ;
        RECT 1987.270 3499.720 1994.030 3499.860 ;
        RECT 1987.270 3499.660 1987.590 3499.720 ;
        RECT 1993.710 3499.660 1994.030 3499.720 ;
        RECT 1993.710 2439.060 1994.030 2439.120 ;
        RECT 2697.050 2439.060 2697.370 2439.120 ;
        RECT 1993.710 2438.920 2697.370 2439.060 ;
        RECT 1993.710 2438.860 1994.030 2438.920 ;
        RECT 2697.050 2438.860 2697.370 2438.920 ;
      LAYER via ;
        RECT 1987.300 3499.660 1987.560 3499.920 ;
        RECT 1993.740 3499.660 1994.000 3499.920 ;
        RECT 1993.740 2438.860 1994.000 2439.120 ;
        RECT 2697.080 2438.860 2697.340 2439.120 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3499.950 1987.500 3517.600 ;
        RECT 1987.300 3499.630 1987.560 3499.950 ;
        RECT 1993.740 3499.630 1994.000 3499.950 ;
        RECT 1993.800 2439.150 1993.940 3499.630 ;
        RECT 1993.740 2438.830 1994.000 2439.150 ;
        RECT 2697.080 2438.830 2697.340 2439.150 ;
        RECT 2697.140 1753.565 2697.280 2438.830 ;
        RECT 2697.070 1753.195 2697.350 1753.565 ;
      LAYER via2 ;
        RECT 2697.070 1753.240 2697.350 1753.520 ;
      LAYER met3 ;
        RECT 2697.045 1753.530 2697.375 1753.545 ;
        RECT 2696.830 1753.215 2697.375 1753.530 ;
        RECT 2696.830 1752.800 2697.130 1753.215 ;
        RECT 2696.000 1752.200 2700.000 1752.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3503.600 1662.830 3503.660 ;
        RECT 2695.670 3503.600 2695.990 3503.660 ;
        RECT 1662.510 3503.460 2695.990 3503.600 ;
        RECT 1662.510 3503.400 1662.830 3503.460 ;
        RECT 2695.670 3503.400 2695.990 3503.460 ;
      LAYER via ;
        RECT 1662.540 3503.400 1662.800 3503.660 ;
        RECT 2695.700 3503.400 2695.960 3503.660 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3503.690 1662.740 3517.600 ;
        RECT 1662.540 3503.370 1662.800 3503.690 ;
        RECT 2695.700 3503.370 2695.960 3503.690 ;
        RECT 2695.760 1786.770 2695.900 3503.370 ;
        RECT 2696.610 1786.770 2696.890 1786.885 ;
        RECT 2695.760 1786.630 2696.890 1786.770 ;
        RECT 2696.610 1786.515 2696.890 1786.630 ;
      LAYER via2 ;
        RECT 2696.610 1786.560 2696.890 1786.840 ;
      LAYER met3 ;
        RECT 2696.585 1786.850 2696.915 1786.865 ;
        RECT 2696.585 1786.550 2698.050 1786.850 ;
        RECT 2696.585 1786.535 2696.915 1786.550 ;
        RECT 2697.750 1784.080 2698.050 1786.550 ;
        RECT 2696.000 1783.480 2700.000 1784.080 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3101.380 1338.530 3101.440 ;
        RECT 2701.650 3101.380 2701.970 3101.440 ;
        RECT 1338.210 3101.240 2701.970 3101.380 ;
        RECT 1338.210 3101.180 1338.530 3101.240 ;
        RECT 2701.650 3101.180 2701.970 3101.240 ;
      LAYER via ;
        RECT 1338.240 3101.180 1338.500 3101.440 ;
        RECT 2701.680 3101.180 2701.940 3101.440 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3101.470 1338.440 3517.600 ;
        RECT 1338.240 3101.150 1338.500 3101.470 ;
        RECT 2701.680 3101.150 2701.940 3101.470 ;
        RECT 2701.740 1815.445 2701.880 3101.150 ;
        RECT 2701.670 1815.075 2701.950 1815.445 ;
      LAYER via2 ;
        RECT 2701.670 1815.120 2701.950 1815.400 ;
      LAYER met3 ;
        RECT 2701.645 1815.410 2701.975 1815.425 ;
        RECT 2699.740 1815.360 2701.975 1815.410 ;
        RECT 2696.000 1815.110 2701.975 1815.360 ;
        RECT 2696.000 1814.760 2700.000 1815.110 ;
        RECT 2701.645 1815.095 2701.975 1815.110 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1242.260 2713.470 1242.320 ;
        RECT 2777.090 1242.260 2777.410 1242.320 ;
        RECT 2713.150 1242.120 2777.410 1242.260 ;
        RECT 2713.150 1242.060 2713.470 1242.120 ;
        RECT 2777.090 1242.060 2777.410 1242.120 ;
        RECT 2777.090 441.560 2777.410 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 2777.090 441.420 2901.150 441.560 ;
        RECT 2777.090 441.360 2777.410 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 2713.180 1242.060 2713.440 1242.320 ;
        RECT 2777.120 1242.060 2777.380 1242.320 ;
        RECT 2777.120 441.360 2777.380 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 2713.170 1246.595 2713.450 1246.965 ;
        RECT 2713.240 1242.350 2713.380 1246.595 ;
        RECT 2713.180 1242.030 2713.440 1242.350 ;
        RECT 2777.120 1242.030 2777.380 1242.350 ;
        RECT 2777.180 441.650 2777.320 1242.030 ;
        RECT 2777.120 441.330 2777.380 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2713.170 1246.640 2713.450 1246.920 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2713.145 1246.930 2713.475 1246.945 ;
        RECT 2699.740 1246.880 2713.475 1246.930 ;
        RECT 2696.000 1246.630 2713.475 1246.880 ;
        RECT 2696.000 1246.280 2700.000 1246.630 ;
        RECT 2713.145 1246.615 2713.475 1246.630 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3502.580 1014.230 3502.640 ;
        RECT 2699.350 3502.580 2699.670 3502.640 ;
        RECT 1013.910 3502.440 2699.670 3502.580 ;
        RECT 1013.910 3502.380 1014.230 3502.440 ;
        RECT 2699.350 3502.380 2699.670 3502.440 ;
      LAYER via ;
        RECT 1013.940 3502.380 1014.200 3502.640 ;
        RECT 2699.380 3502.380 2699.640 3502.640 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3502.670 1014.140 3517.600 ;
        RECT 1013.940 3502.350 1014.200 3502.670 ;
        RECT 2699.380 3502.350 2699.640 3502.670 ;
        RECT 2699.440 1848.085 2699.580 3502.350 ;
        RECT 2699.370 1847.715 2699.650 1848.085 ;
      LAYER via2 ;
        RECT 2699.370 1847.760 2699.650 1848.040 ;
      LAYER met3 ;
        RECT 2699.345 1848.050 2699.675 1848.065 ;
        RECT 2699.345 1847.735 2699.890 1848.050 ;
        RECT 2699.590 1847.320 2699.890 1847.735 ;
        RECT 2696.000 1846.720 2700.000 1847.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.885 689.380 3517.600 ;
        RECT 689.170 3503.515 689.450 3503.885 ;
      LAYER via2 ;
        RECT 689.170 3503.560 689.450 3503.840 ;
      LAYER met3 ;
        RECT 689.145 3503.850 689.475 3503.865 ;
        RECT 2691.270 3503.850 2691.650 3503.860 ;
        RECT 689.145 3503.550 2691.650 3503.850 ;
        RECT 689.145 3503.535 689.475 3503.550 ;
        RECT 2691.270 3503.540 2691.650 3503.550 ;
        RECT 2696.790 1881.060 2697.170 1881.380 ;
        RECT 2696.830 1878.600 2697.130 1881.060 ;
        RECT 2696.000 1878.000 2700.000 1878.600 ;
      LAYER via3 ;
        RECT 2691.300 3503.540 2691.620 3503.860 ;
        RECT 2696.820 1881.060 2697.140 1881.380 ;
      LAYER met4 ;
        RECT 2691.295 3503.535 2691.625 3503.865 ;
        RECT 2691.310 2137.050 2691.610 3503.535 ;
        RECT 2690.390 2136.750 2691.610 2137.050 ;
        RECT 2690.390 2130.250 2690.690 2136.750 ;
        RECT 2690.390 2129.950 2691.610 2130.250 ;
        RECT 2691.310 1997.650 2691.610 2129.950 ;
        RECT 2690.390 1997.350 2691.610 1997.650 ;
        RECT 2690.390 1994.250 2690.690 1997.350 ;
        RECT 2690.390 1993.950 2691.610 1994.250 ;
        RECT 2691.310 1888.850 2691.610 1993.950 ;
        RECT 2691.310 1888.550 2692.530 1888.850 ;
        RECT 2692.230 1881.370 2692.530 1888.550 ;
        RECT 2696.815 1881.370 2697.145 1881.385 ;
        RECT 2692.230 1881.070 2697.145 1881.370 ;
        RECT 2696.815 1881.055 2697.145 1881.070 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3501.900 365.170 3501.960 ;
        RECT 2700.730 3501.900 2701.050 3501.960 ;
        RECT 364.850 3501.760 2701.050 3501.900 ;
        RECT 364.850 3501.700 365.170 3501.760 ;
        RECT 2700.730 3501.700 2701.050 3501.760 ;
      LAYER via ;
        RECT 364.880 3501.700 365.140 3501.960 ;
        RECT 2700.760 3501.700 2701.020 3501.960 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3501.990 365.080 3517.600 ;
        RECT 364.880 3501.670 365.140 3501.990 ;
        RECT 2700.760 3501.670 2701.020 3501.990 ;
        RECT 2700.820 1910.645 2700.960 3501.670 ;
        RECT 2700.750 1910.275 2701.030 1910.645 ;
      LAYER via2 ;
        RECT 2700.750 1910.320 2701.030 1910.600 ;
      LAYER met3 ;
        RECT 2700.725 1910.610 2701.055 1910.625 ;
        RECT 2699.740 1910.560 2701.055 1910.610 ;
        RECT 2696.000 1910.310 2701.055 1910.560 ;
        RECT 2696.000 1909.960 2700.000 1910.310 ;
        RECT 2700.725 1910.295 2701.055 1910.310 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 2699.550 3501.810 2699.930 3501.820 ;
        RECT 40.545 3501.510 2699.930 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 2699.550 3501.500 2699.930 3501.510 ;
        RECT 2699.550 1942.260 2699.930 1942.580 ;
        RECT 2699.590 1941.840 2699.890 1942.260 ;
        RECT 2696.000 1941.240 2700.000 1941.840 ;
      LAYER via3 ;
        RECT 2699.580 3501.500 2699.900 3501.820 ;
        RECT 2699.580 1942.260 2699.900 1942.580 ;
      LAYER met4 ;
        RECT 2699.575 3501.495 2699.905 3501.825 ;
        RECT 2699.590 1942.585 2699.890 3501.495 ;
        RECT 2699.575 1942.255 2699.905 1942.585 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 2701.190 3263.900 2701.510 3263.960 ;
        RECT 15.250 3263.760 2701.510 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 2701.190 3263.700 2701.510 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 2701.220 3263.700 2701.480 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 2701.220 3263.670 2701.480 3263.990 ;
        RECT 2701.280 1973.885 2701.420 3263.670 ;
        RECT 2701.210 1973.515 2701.490 1973.885 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
        RECT 2701.210 1973.560 2701.490 1973.840 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
        RECT 2701.185 1973.850 2701.515 1973.865 ;
        RECT 2699.740 1973.800 2701.515 1973.850 ;
        RECT 2696.000 1973.550 2701.515 1973.800 ;
        RECT 2696.000 1973.200 2700.000 1973.550 ;
        RECT 2701.185 1973.535 2701.515 1973.550 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 2391.120 17.410 2391.180 ;
        RECT 2714.070 2391.120 2714.390 2391.180 ;
        RECT 17.090 2390.980 2714.390 2391.120 ;
        RECT 17.090 2390.920 17.410 2390.980 ;
        RECT 2714.070 2390.920 2714.390 2390.980 ;
      LAYER via ;
        RECT 17.120 2390.920 17.380 2391.180 ;
        RECT 2714.100 2390.920 2714.360 2391.180 ;
      LAYER met2 ;
        RECT 17.110 2979.915 17.390 2980.285 ;
        RECT 17.180 2391.210 17.320 2979.915 ;
        RECT 17.120 2390.890 17.380 2391.210 ;
        RECT 2714.100 2390.890 2714.360 2391.210 ;
        RECT 2714.160 2005.165 2714.300 2390.890 ;
        RECT 2714.090 2004.795 2714.370 2005.165 ;
      LAYER via2 ;
        RECT 17.110 2979.960 17.390 2980.240 ;
        RECT 2714.090 2004.840 2714.370 2005.120 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 17.085 2980.250 17.415 2980.265 ;
        RECT -4.800 2979.950 17.415 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 17.085 2979.935 17.415 2979.950 ;
        RECT 2714.065 2005.130 2714.395 2005.145 ;
        RECT 2699.740 2005.080 2714.395 2005.130 ;
        RECT 2696.000 2004.830 2714.395 2005.080 ;
        RECT 2696.000 2004.480 2700.000 2004.830 ;
        RECT 2714.065 2004.815 2714.395 2004.830 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2391.460 18.790 2391.520 ;
        RECT 2714.530 2391.460 2714.850 2391.520 ;
        RECT 18.470 2391.320 2714.850 2391.460 ;
        RECT 18.470 2391.260 18.790 2391.320 ;
        RECT 2714.530 2391.260 2714.850 2391.320 ;
      LAYER via ;
        RECT 18.500 2391.260 18.760 2391.520 ;
        RECT 2714.560 2391.260 2714.820 2391.520 ;
      LAYER met2 ;
        RECT 18.490 2692.955 18.770 2693.325 ;
        RECT 18.560 2391.550 18.700 2692.955 ;
        RECT 18.500 2391.230 18.760 2391.550 ;
        RECT 2714.560 2391.230 2714.820 2391.550 ;
        RECT 2714.620 2037.125 2714.760 2391.230 ;
        RECT 2714.550 2036.755 2714.830 2037.125 ;
      LAYER via2 ;
        RECT 18.490 2693.000 18.770 2693.280 ;
        RECT 2714.550 2036.800 2714.830 2037.080 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 18.465 2693.290 18.795 2693.305 ;
        RECT -4.800 2692.990 18.795 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 18.465 2692.975 18.795 2692.990 ;
        RECT 2714.525 2037.090 2714.855 2037.105 ;
        RECT 2699.740 2037.040 2714.855 2037.090 ;
        RECT 2696.000 2036.790 2714.855 2037.040 ;
        RECT 2696.000 2036.440 2700.000 2036.790 ;
        RECT 2714.525 2036.775 2714.855 2036.790 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2401.320 16.030 2401.380 ;
        RECT 2703.030 2401.320 2703.350 2401.380 ;
        RECT 15.710 2401.180 2703.350 2401.320 ;
        RECT 15.710 2401.120 16.030 2401.180 ;
        RECT 2703.030 2401.120 2703.350 2401.180 ;
      LAYER via ;
        RECT 15.740 2401.120 16.000 2401.380 ;
        RECT 2703.060 2401.120 2703.320 2401.380 ;
      LAYER met2 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
        RECT 15.800 2401.410 15.940 2405.315 ;
        RECT 15.740 2401.090 16.000 2401.410 ;
        RECT 2703.060 2401.090 2703.320 2401.410 ;
        RECT 2703.120 2068.405 2703.260 2401.090 ;
        RECT 2703.050 2068.035 2703.330 2068.405 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
        RECT 2703.050 2068.080 2703.330 2068.360 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
        RECT 2703.025 2068.370 2703.355 2068.385 ;
        RECT 2699.740 2068.320 2703.355 2068.370 ;
        RECT 2696.000 2068.070 2703.355 2068.320 ;
        RECT 2696.000 2067.720 2700.000 2068.070 ;
        RECT 2703.025 2068.055 2703.355 2068.070 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1300.030 2390.440 1300.350 2390.500 ;
        RECT 2715.450 2390.440 2715.770 2390.500 ;
        RECT 1300.030 2390.300 2715.770 2390.440 ;
        RECT 1300.030 2390.240 1300.350 2390.300 ;
        RECT 2715.450 2390.240 2715.770 2390.300 ;
        RECT 16.170 2125.240 16.490 2125.300 ;
        RECT 1300.030 2125.240 1300.350 2125.300 ;
        RECT 16.170 2125.100 1300.350 2125.240 ;
        RECT 16.170 2125.040 16.490 2125.100 ;
        RECT 1300.030 2125.040 1300.350 2125.100 ;
      LAYER via ;
        RECT 1300.060 2390.240 1300.320 2390.500 ;
        RECT 2715.480 2390.240 2715.740 2390.500 ;
        RECT 16.200 2125.040 16.460 2125.300 ;
        RECT 1300.060 2125.040 1300.320 2125.300 ;
      LAYER met2 ;
        RECT 1300.060 2390.210 1300.320 2390.530 ;
        RECT 2715.480 2390.210 2715.740 2390.530 ;
        RECT 1300.120 2125.330 1300.260 2390.210 ;
        RECT 16.200 2125.010 16.460 2125.330 ;
        RECT 1300.060 2125.010 1300.320 2125.330 ;
        RECT 16.260 2118.725 16.400 2125.010 ;
        RECT 16.190 2118.355 16.470 2118.725 ;
        RECT 2715.540 2100.365 2715.680 2390.210 ;
        RECT 2715.470 2099.995 2715.750 2100.365 ;
      LAYER via2 ;
        RECT 16.190 2118.400 16.470 2118.680 ;
        RECT 2715.470 2100.040 2715.750 2100.320 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.165 2118.690 16.495 2118.705 ;
        RECT -4.800 2118.390 16.495 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.165 2118.375 16.495 2118.390 ;
        RECT 2715.445 2100.330 2715.775 2100.345 ;
        RECT 2699.740 2100.280 2715.775 2100.330 ;
        RECT 2696.000 2100.030 2715.775 2100.280 ;
        RECT 2696.000 2099.680 2700.000 2100.030 ;
        RECT 2715.445 2100.015 2715.775 2100.030 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1302.790 2395.540 1303.110 2395.600 ;
        RECT 2703.950 2395.540 2704.270 2395.600 ;
        RECT 1302.790 2395.400 2704.270 2395.540 ;
        RECT 1302.790 2395.340 1303.110 2395.400 ;
        RECT 2703.950 2395.340 2704.270 2395.400 ;
        RECT 15.710 1835.220 16.030 1835.280 ;
        RECT 1302.790 1835.220 1303.110 1835.280 ;
        RECT 15.710 1835.080 1303.110 1835.220 ;
        RECT 15.710 1835.020 16.030 1835.080 ;
        RECT 1302.790 1835.020 1303.110 1835.080 ;
      LAYER via ;
        RECT 1302.820 2395.340 1303.080 2395.600 ;
        RECT 2703.980 2395.340 2704.240 2395.600 ;
        RECT 15.740 1835.020 16.000 1835.280 ;
        RECT 1302.820 1835.020 1303.080 1835.280 ;
      LAYER met2 ;
        RECT 1302.820 2395.310 1303.080 2395.630 ;
        RECT 2703.980 2395.310 2704.240 2395.630 ;
        RECT 1302.880 1835.310 1303.020 2395.310 ;
        RECT 2704.040 2131.645 2704.180 2395.310 ;
        RECT 2703.970 2131.275 2704.250 2131.645 ;
        RECT 15.740 1834.990 16.000 1835.310 ;
        RECT 1302.820 1834.990 1303.080 1835.310 ;
        RECT 15.800 1831.085 15.940 1834.990 ;
        RECT 15.730 1830.715 16.010 1831.085 ;
      LAYER via2 ;
        RECT 2703.970 2131.320 2704.250 2131.600 ;
        RECT 15.730 1830.760 16.010 1831.040 ;
      LAYER met3 ;
        RECT 2703.945 2131.610 2704.275 2131.625 ;
        RECT 2699.740 2131.560 2704.275 2131.610 ;
        RECT 2696.000 2131.310 2704.275 2131.560 ;
        RECT 2696.000 2130.960 2700.000 2131.310 ;
        RECT 2703.945 2131.295 2704.275 2131.310 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 15.705 1831.050 16.035 1831.065 ;
        RECT -4.800 1830.750 16.035 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 15.705 1830.735 16.035 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1276.600 2713.470 1276.660 ;
        RECT 2783.990 1276.600 2784.310 1276.660 ;
        RECT 2713.150 1276.460 2784.310 1276.600 ;
        RECT 2713.150 1276.400 2713.470 1276.460 ;
        RECT 2783.990 1276.400 2784.310 1276.460 ;
        RECT 2783.990 676.160 2784.310 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2783.990 676.020 2901.150 676.160 ;
        RECT 2783.990 675.960 2784.310 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 2713.180 1276.400 2713.440 1276.660 ;
        RECT 2784.020 1276.400 2784.280 1276.660 ;
        RECT 2784.020 675.960 2784.280 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 2713.170 1278.555 2713.450 1278.925 ;
        RECT 2713.240 1276.690 2713.380 1278.555 ;
        RECT 2713.180 1276.370 2713.440 1276.690 ;
        RECT 2784.020 1276.370 2784.280 1276.690 ;
        RECT 2784.080 676.250 2784.220 1276.370 ;
        RECT 2784.020 675.930 2784.280 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2713.170 1278.600 2713.450 1278.880 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2713.145 1278.890 2713.475 1278.905 ;
        RECT 2699.740 1278.840 2713.475 1278.890 ;
        RECT 2696.000 1278.590 2713.475 1278.840 ;
        RECT 2696.000 1278.240 2700.000 1278.590 ;
        RECT 2713.145 1278.575 2713.475 1278.590 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1301.410 2391.800 1301.730 2391.860 ;
        RECT 2717.750 2391.800 2718.070 2391.860 ;
        RECT 1301.410 2391.660 2718.070 2391.800 ;
        RECT 1301.410 2391.600 1301.730 2391.660 ;
        RECT 2717.750 2391.600 2718.070 2391.660 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 1301.410 1545.540 1301.730 1545.600 ;
        RECT 16.630 1545.400 1301.730 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 1301.410 1545.340 1301.730 1545.400 ;
      LAYER via ;
        RECT 1301.440 2391.600 1301.700 2391.860 ;
        RECT 2717.780 2391.600 2718.040 2391.860 ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 1301.440 1545.340 1301.700 1545.600 ;
      LAYER met2 ;
        RECT 1301.440 2391.570 1301.700 2391.890 ;
        RECT 2717.780 2391.570 2718.040 2391.890 ;
        RECT 1301.500 1545.630 1301.640 2391.570 ;
        RECT 2717.840 2162.925 2717.980 2391.570 ;
        RECT 2717.770 2162.555 2718.050 2162.925 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 1301.440 1545.310 1301.700 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 2717.770 2162.600 2718.050 2162.880 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT 2717.745 2162.890 2718.075 2162.905 ;
        RECT 2699.740 2162.840 2718.075 2162.890 ;
        RECT 2696.000 2162.590 2718.075 2162.840 ;
        RECT 2696.000 2162.240 2700.000 2162.590 ;
        RECT 2717.745 2162.575 2718.075 2162.590 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2712.230 1216.080 2712.550 1216.140 ;
        RECT 2713.610 1216.080 2713.930 1216.140 ;
        RECT 2712.230 1215.940 2713.930 1216.080 ;
        RECT 2712.230 1215.880 2712.550 1215.940 ;
        RECT 2713.610 1215.880 2713.930 1215.940 ;
        RECT 17.090 1205.540 17.410 1205.600 ;
        RECT 2713.610 1205.540 2713.930 1205.600 ;
        RECT 17.090 1205.400 2713.930 1205.540 ;
        RECT 17.090 1205.340 17.410 1205.400 ;
        RECT 2713.610 1205.340 2713.930 1205.400 ;
      LAYER via ;
        RECT 2712.260 1215.880 2712.520 1216.140 ;
        RECT 2713.640 1215.880 2713.900 1216.140 ;
        RECT 17.120 1205.340 17.380 1205.600 ;
        RECT 2713.640 1205.340 2713.900 1205.600 ;
      LAYER met2 ;
        RECT 2712.250 2194.515 2712.530 2194.885 ;
        RECT 17.110 1328.195 17.390 1328.565 ;
        RECT 17.180 1205.630 17.320 1328.195 ;
        RECT 2712.320 1216.170 2712.460 2194.515 ;
        RECT 2712.260 1215.850 2712.520 1216.170 ;
        RECT 2713.640 1215.850 2713.900 1216.170 ;
        RECT 2713.700 1205.630 2713.840 1215.850 ;
        RECT 17.120 1205.310 17.380 1205.630 ;
        RECT 2713.640 1205.310 2713.900 1205.630 ;
      LAYER via2 ;
        RECT 2712.250 2194.560 2712.530 2194.840 ;
        RECT 17.110 1328.240 17.390 1328.520 ;
      LAYER met3 ;
        RECT 2712.225 2194.850 2712.555 2194.865 ;
        RECT 2699.740 2194.800 2712.555 2194.850 ;
        RECT 2696.000 2194.550 2712.555 2194.800 ;
        RECT 2696.000 2194.200 2700.000 2194.550 ;
        RECT 2712.225 2194.535 2712.555 2194.550 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 17.085 1328.530 17.415 1328.545 ;
        RECT -4.800 1328.230 17.415 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 17.085 1328.215 17.415 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 2711.770 1117.820 2712.090 1117.880 ;
        RECT 15.710 1117.680 2712.090 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 2711.770 1117.620 2712.090 1117.680 ;
      LAYER via ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 2711.800 1117.620 2712.060 1117.880 ;
      LAYER met2 ;
        RECT 2711.790 2225.795 2712.070 2226.165 ;
        RECT 2711.860 1117.910 2712.000 2225.795 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 2711.800 1117.590 2712.060 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 2711.790 2225.840 2712.070 2226.120 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT 2711.765 2226.130 2712.095 2226.145 ;
        RECT 2699.740 2226.080 2712.095 2226.130 ;
        RECT 2696.000 2225.830 2712.095 2226.080 ;
        RECT 2696.000 2225.480 2700.000 2225.830 ;
        RECT 2711.765 2225.815 2712.095 2225.830 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 1003.920 17.870 1003.980 ;
        RECT 2712.690 1003.920 2713.010 1003.980 ;
        RECT 17.550 1003.780 2713.010 1003.920 ;
        RECT 17.550 1003.720 17.870 1003.780 ;
        RECT 2712.690 1003.720 2713.010 1003.780 ;
      LAYER via ;
        RECT 17.580 1003.720 17.840 1003.980 ;
        RECT 2712.720 1003.720 2712.980 1003.980 ;
      LAYER met2 ;
        RECT 2712.710 2257.755 2712.990 2258.125 ;
        RECT 2712.780 1004.010 2712.920 2257.755 ;
        RECT 17.580 1003.690 17.840 1004.010 ;
        RECT 2712.720 1003.690 2712.980 1004.010 ;
        RECT 17.640 897.445 17.780 1003.690 ;
        RECT 17.570 897.075 17.850 897.445 ;
      LAYER via2 ;
        RECT 2712.710 2257.800 2712.990 2258.080 ;
        RECT 17.570 897.120 17.850 897.400 ;
      LAYER met3 ;
        RECT 2712.685 2258.090 2713.015 2258.105 ;
        RECT 2699.740 2258.040 2713.015 2258.090 ;
        RECT 2696.000 2257.790 2713.015 2258.040 ;
        RECT 2696.000 2257.440 2700.000 2257.790 ;
        RECT 2712.685 2257.775 2713.015 2257.790 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 17.545 897.410 17.875 897.425 ;
        RECT -4.800 897.110 17.875 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 17.545 897.095 17.875 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.030 1003.155 18.310 1003.525 ;
        RECT 18.100 681.885 18.240 1003.155 ;
        RECT 18.030 681.515 18.310 681.885 ;
      LAYER via2 ;
        RECT 18.030 1003.200 18.310 1003.480 ;
        RECT 18.030 681.560 18.310 681.840 ;
      LAYER met3 ;
        RECT 2716.110 2289.370 2716.490 2289.380 ;
        RECT 2699.740 2289.320 2716.490 2289.370 ;
        RECT 2696.000 2289.070 2716.490 2289.320 ;
        RECT 2696.000 2288.720 2700.000 2289.070 ;
        RECT 2716.110 2289.060 2716.490 2289.070 ;
        RECT 18.005 1003.490 18.335 1003.505 ;
        RECT 2716.110 1003.490 2716.490 1003.500 ;
        RECT 18.005 1003.190 2716.490 1003.490 ;
        RECT 18.005 1003.175 18.335 1003.190 ;
        RECT 2716.110 1003.180 2716.490 1003.190 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 18.005 681.850 18.335 681.865 ;
        RECT -4.800 681.550 18.335 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 18.005 681.535 18.335 681.550 ;
      LAYER via3 ;
        RECT 2716.140 2289.060 2716.460 2289.380 ;
        RECT 2716.140 1003.180 2716.460 1003.500 ;
      LAYER met4 ;
        RECT 2716.135 2289.055 2716.465 2289.385 ;
        RECT 2716.150 1003.505 2716.450 2289.055 ;
        RECT 2716.135 1003.175 2716.465 1003.505 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2698.890 1697.520 2699.210 1697.580 ;
        RECT 2699.810 1697.520 2700.130 1697.580 ;
        RECT 2698.890 1697.380 2700.130 1697.520 ;
        RECT 2698.890 1697.320 2699.210 1697.380 ;
        RECT 2699.810 1697.320 2700.130 1697.380 ;
        RECT 724.570 468.420 724.890 468.480 ;
        RECT 772.410 468.420 772.730 468.480 ;
        RECT 724.570 468.280 772.730 468.420 ;
        RECT 724.570 468.220 724.890 468.280 ;
        RECT 772.410 468.220 772.730 468.280 ;
        RECT 193.270 467.740 193.590 467.800 ;
        RECT 240.650 467.740 240.970 467.800 ;
        RECT 193.270 467.600 240.970 467.740 ;
        RECT 193.270 467.540 193.590 467.600 ;
        RECT 240.650 467.540 240.970 467.600 ;
      LAYER via ;
        RECT 2698.920 1697.320 2699.180 1697.580 ;
        RECT 2699.840 1697.320 2700.100 1697.580 ;
        RECT 724.600 468.220 724.860 468.480 ;
        RECT 772.440 468.220 772.700 468.480 ;
        RECT 193.300 467.540 193.560 467.800 ;
        RECT 240.680 467.540 240.940 467.800 ;
      LAYER met2 ;
        RECT 2699.830 1744.355 2700.110 1744.725 ;
        RECT 2699.900 1697.610 2700.040 1744.355 ;
        RECT 2698.920 1697.290 2699.180 1697.610 ;
        RECT 2699.840 1697.290 2700.100 1697.610 ;
        RECT 2698.980 1656.325 2699.120 1697.290 ;
        RECT 2698.910 1655.955 2699.190 1656.325 ;
        RECT 2699.370 1459.435 2699.650 1459.805 ;
        RECT 2699.440 1395.885 2699.580 1459.435 ;
        RECT 2699.370 1395.515 2699.650 1395.885 ;
        RECT 2698.910 1366.955 2699.190 1367.325 ;
        RECT 2698.980 1325.165 2699.120 1366.955 ;
        RECT 2698.910 1324.795 2699.190 1325.165 ;
        RECT 2699.830 1079.995 2700.110 1080.365 ;
        RECT 2699.900 1015.085 2700.040 1079.995 ;
        RECT 2699.830 1014.715 2700.110 1015.085 ;
        RECT 2699.830 965.755 2700.110 966.125 ;
        RECT 2699.900 918.525 2700.040 965.755 ;
        RECT 2699.830 918.155 2700.110 918.525 ;
        RECT 2700.750 835.195 2701.030 835.565 ;
        RECT 2700.820 821.285 2700.960 835.195 ;
        RECT 2700.750 820.915 2701.030 821.285 ;
        RECT 2699.830 812.755 2700.110 813.125 ;
        RECT 2699.900 766.205 2700.040 812.755 ;
        RECT 2699.830 765.835 2700.110 766.205 ;
        RECT 2699.830 738.635 2700.110 739.005 ;
        RECT 2699.900 724.725 2700.040 738.635 ;
        RECT 2699.830 724.355 2700.110 724.725 ;
        RECT 2699.830 603.315 2700.110 603.685 ;
        RECT 2699.900 579.885 2700.040 603.315 ;
        RECT 2699.830 579.515 2700.110 579.885 ;
        RECT 362.110 469.355 362.390 469.725 ;
        RECT 458.710 469.355 458.990 469.725 ;
        RECT 555.310 469.355 555.590 469.725 ;
        RECT 651.910 469.355 652.190 469.725 ;
        RECT 362.180 468.365 362.320 469.355 ;
        RECT 458.780 468.365 458.920 469.355 ;
        RECT 555.380 468.365 555.520 469.355 ;
        RECT 651.980 468.365 652.120 469.355 ;
        RECT 772.430 468.675 772.710 469.045 ;
        RECT 772.500 468.510 772.640 468.675 ;
        RECT 724.600 468.365 724.860 468.510 ;
        RECT 240.670 467.995 240.950 468.365 ;
        RECT 362.110 467.995 362.390 468.365 ;
        RECT 458.710 467.995 458.990 468.365 ;
        RECT 555.310 467.995 555.590 468.365 ;
        RECT 651.910 467.995 652.190 468.365 ;
        RECT 700.210 467.995 700.490 468.365 ;
        RECT 724.590 467.995 724.870 468.365 ;
        RECT 772.440 468.190 772.700 468.510 ;
        RECT 240.740 467.830 240.880 467.995 ;
        RECT 193.300 467.685 193.560 467.830 ;
        RECT 193.290 467.315 193.570 467.685 ;
        RECT 240.680 467.510 240.940 467.830 ;
        RECT 700.280 466.325 700.420 467.995 ;
        RECT 700.210 465.955 700.490 466.325 ;
      LAYER via2 ;
        RECT 2699.830 1744.400 2700.110 1744.680 ;
        RECT 2698.910 1656.000 2699.190 1656.280 ;
        RECT 2699.370 1459.480 2699.650 1459.760 ;
        RECT 2699.370 1395.560 2699.650 1395.840 ;
        RECT 2698.910 1367.000 2699.190 1367.280 ;
        RECT 2698.910 1324.840 2699.190 1325.120 ;
        RECT 2699.830 1080.040 2700.110 1080.320 ;
        RECT 2699.830 1014.760 2700.110 1015.040 ;
        RECT 2699.830 965.800 2700.110 966.080 ;
        RECT 2699.830 918.200 2700.110 918.480 ;
        RECT 2700.750 835.240 2701.030 835.520 ;
        RECT 2700.750 820.960 2701.030 821.240 ;
        RECT 2699.830 812.800 2700.110 813.080 ;
        RECT 2699.830 765.880 2700.110 766.160 ;
        RECT 2699.830 738.680 2700.110 738.960 ;
        RECT 2699.830 724.400 2700.110 724.680 ;
        RECT 2699.830 603.360 2700.110 603.640 ;
        RECT 2699.830 579.560 2700.110 579.840 ;
        RECT 362.110 469.400 362.390 469.680 ;
        RECT 458.710 469.400 458.990 469.680 ;
        RECT 555.310 469.400 555.590 469.680 ;
        RECT 651.910 469.400 652.190 469.680 ;
        RECT 772.430 468.720 772.710 469.000 ;
        RECT 240.670 468.040 240.950 468.320 ;
        RECT 362.110 468.040 362.390 468.320 ;
        RECT 458.710 468.040 458.990 468.320 ;
        RECT 555.310 468.040 555.590 468.320 ;
        RECT 651.910 468.040 652.190 468.320 ;
        RECT 700.210 468.040 700.490 468.320 ;
        RECT 724.590 468.040 724.870 468.320 ;
        RECT 193.290 467.360 193.570 467.640 ;
        RECT 700.210 466.000 700.490 466.280 ;
      LAYER met3 ;
        RECT 2696.000 2320.680 2700.000 2321.280 ;
        RECT 2698.670 2318.620 2698.970 2320.680 ;
        RECT 2698.630 2318.300 2699.010 2318.620 ;
        RECT 2698.630 2260.130 2699.010 2260.140 ;
        RECT 2702.310 2260.130 2702.690 2260.140 ;
        RECT 2698.630 2259.830 2702.690 2260.130 ;
        RECT 2698.630 2259.820 2699.010 2259.830 ;
        RECT 2702.310 2259.820 2702.690 2259.830 ;
        RECT 2698.630 2211.850 2699.010 2211.860 ;
        RECT 2702.310 2211.850 2702.690 2211.860 ;
        RECT 2698.630 2211.550 2702.690 2211.850 ;
        RECT 2698.630 2211.540 2699.010 2211.550 ;
        RECT 2702.310 2211.540 2702.690 2211.550 ;
        RECT 2698.630 2163.570 2699.010 2163.580 ;
        RECT 2702.310 2163.570 2702.690 2163.580 ;
        RECT 2698.630 2163.270 2702.690 2163.570 ;
        RECT 2698.630 2163.260 2699.010 2163.270 ;
        RECT 2702.310 2163.260 2702.690 2163.270 ;
        RECT 2698.630 2067.010 2699.010 2067.020 ;
        RECT 2702.310 2067.010 2702.690 2067.020 ;
        RECT 2698.630 2066.710 2702.690 2067.010 ;
        RECT 2698.630 2066.700 2699.010 2066.710 ;
        RECT 2702.310 2066.700 2702.690 2066.710 ;
        RECT 2698.630 2018.730 2699.010 2018.740 ;
        RECT 2702.310 2018.730 2702.690 2018.740 ;
        RECT 2698.630 2018.430 2702.690 2018.730 ;
        RECT 2698.630 2018.420 2699.010 2018.430 ;
        RECT 2702.310 2018.420 2702.690 2018.430 ;
        RECT 2698.630 1905.170 2699.010 1905.180 ;
        RECT 2702.310 1905.170 2702.690 1905.180 ;
        RECT 2698.630 1904.870 2702.690 1905.170 ;
        RECT 2698.630 1904.860 2699.010 1904.870 ;
        RECT 2702.310 1904.860 2702.690 1904.870 ;
        RECT 2698.630 1745.060 2699.010 1745.380 ;
        RECT 2698.670 1744.690 2698.970 1745.060 ;
        RECT 2699.805 1744.690 2700.135 1744.705 ;
        RECT 2698.670 1744.390 2700.135 1744.690 ;
        RECT 2699.805 1744.375 2700.135 1744.390 ;
        RECT 2698.885 1656.290 2699.215 1656.305 ;
        RECT 2699.550 1656.290 2699.930 1656.300 ;
        RECT 2698.885 1655.990 2699.930 1656.290 ;
        RECT 2698.885 1655.975 2699.215 1655.990 ;
        RECT 2699.550 1655.980 2699.930 1655.990 ;
        RECT 2699.550 1511.820 2699.930 1512.140 ;
        RECT 2699.590 1510.770 2699.890 1511.820 ;
        RECT 2700.470 1510.770 2700.850 1510.780 ;
        RECT 2699.590 1510.470 2700.850 1510.770 ;
        RECT 2700.470 1510.460 2700.850 1510.470 ;
        RECT 2699.345 1459.770 2699.675 1459.785 ;
        RECT 2700.470 1459.770 2700.850 1459.780 ;
        RECT 2699.345 1459.470 2700.850 1459.770 ;
        RECT 2699.345 1459.455 2699.675 1459.470 ;
        RECT 2700.470 1459.460 2700.850 1459.470 ;
        RECT 2699.345 1395.850 2699.675 1395.865 ;
        RECT 2700.470 1395.850 2700.850 1395.860 ;
        RECT 2699.345 1395.550 2700.850 1395.850 ;
        RECT 2699.345 1395.535 2699.675 1395.550 ;
        RECT 2700.470 1395.540 2700.850 1395.550 ;
        RECT 2698.885 1367.290 2699.215 1367.305 ;
        RECT 2700.470 1367.290 2700.850 1367.300 ;
        RECT 2698.885 1366.990 2700.850 1367.290 ;
        RECT 2698.885 1366.975 2699.215 1366.990 ;
        RECT 2700.470 1366.980 2700.850 1366.990 ;
        RECT 2698.885 1325.140 2699.215 1325.145 ;
        RECT 2698.630 1325.130 2699.215 1325.140 ;
        RECT 2698.430 1324.830 2699.215 1325.130 ;
        RECT 2698.630 1324.820 2699.215 1324.830 ;
        RECT 2698.885 1324.815 2699.215 1324.820 ;
        RECT 2698.630 1318.330 2699.010 1318.340 ;
        RECT 2698.630 1318.030 2699.890 1318.330 ;
        RECT 2698.630 1318.020 2699.010 1318.030 ;
        RECT 2699.590 1317.660 2699.890 1318.030 ;
        RECT 2699.550 1317.340 2699.930 1317.660 ;
        RECT 2699.805 1080.330 2700.135 1080.345 ;
        RECT 2700.470 1080.330 2700.850 1080.340 ;
        RECT 2699.805 1080.030 2700.850 1080.330 ;
        RECT 2699.805 1080.015 2700.135 1080.030 ;
        RECT 2700.470 1080.020 2700.850 1080.030 ;
        RECT 2699.805 1015.060 2700.135 1015.065 ;
        RECT 2699.550 1015.050 2700.135 1015.060 ;
        RECT 2699.350 1014.750 2700.135 1015.050 ;
        RECT 2699.550 1014.740 2700.135 1014.750 ;
        RECT 2699.805 1014.735 2700.135 1014.740 ;
        RECT 2699.550 980.060 2699.930 980.380 ;
        RECT 2699.590 979.010 2699.890 980.060 ;
        RECT 2700.470 979.010 2700.850 979.020 ;
        RECT 2699.590 978.710 2700.850 979.010 ;
        RECT 2700.470 978.700 2700.850 978.710 ;
        RECT 2699.805 966.090 2700.135 966.105 ;
        RECT 2700.470 966.090 2700.850 966.100 ;
        RECT 2699.805 965.790 2700.850 966.090 ;
        RECT 2699.805 965.775 2700.135 965.790 ;
        RECT 2700.470 965.780 2700.850 965.790 ;
        RECT 2699.805 918.500 2700.135 918.505 ;
        RECT 2699.550 918.490 2700.135 918.500 ;
        RECT 2699.350 918.190 2700.135 918.490 ;
        RECT 2699.550 918.180 2700.135 918.190 ;
        RECT 2699.805 918.175 2700.135 918.180 ;
        RECT 2699.550 883.500 2699.930 883.820 ;
        RECT 2699.590 882.450 2699.890 883.500 ;
        RECT 2700.470 882.450 2700.850 882.460 ;
        RECT 2699.590 882.150 2700.850 882.450 ;
        RECT 2700.470 882.140 2700.850 882.150 ;
        RECT 2700.725 835.540 2701.055 835.545 ;
        RECT 2700.470 835.530 2701.055 835.540 ;
        RECT 2700.470 835.230 2701.280 835.530 ;
        RECT 2700.470 835.220 2701.055 835.230 ;
        RECT 2700.725 835.215 2701.055 835.220 ;
        RECT 2700.725 821.260 2701.055 821.265 ;
        RECT 2700.470 821.250 2701.055 821.260 ;
        RECT 2700.270 820.950 2701.055 821.250 ;
        RECT 2700.470 820.940 2701.055 820.950 ;
        RECT 2700.725 820.935 2701.055 820.940 ;
        RECT 2699.550 813.460 2699.930 813.780 ;
        RECT 2699.590 813.105 2699.890 813.460 ;
        RECT 2699.590 812.790 2700.135 813.105 ;
        RECT 2699.805 812.775 2700.135 812.790 ;
        RECT 2699.805 766.170 2700.135 766.185 ;
        RECT 2700.470 766.170 2700.850 766.180 ;
        RECT 2699.805 765.870 2700.850 766.170 ;
        RECT 2699.805 765.855 2700.135 765.870 ;
        RECT 2700.470 765.860 2700.850 765.870 ;
        RECT 2699.805 738.970 2700.135 738.985 ;
        RECT 2700.470 738.970 2700.850 738.980 ;
        RECT 2699.805 738.670 2700.850 738.970 ;
        RECT 2699.805 738.655 2700.135 738.670 ;
        RECT 2700.470 738.660 2700.850 738.670 ;
        RECT 2698.630 724.690 2699.010 724.700 ;
        RECT 2699.805 724.690 2700.135 724.705 ;
        RECT 2698.630 724.390 2700.135 724.690 ;
        RECT 2698.630 724.380 2699.010 724.390 ;
        RECT 2699.805 724.375 2700.135 724.390 ;
        RECT 2699.805 603.660 2700.135 603.665 ;
        RECT 2699.550 603.650 2700.135 603.660 ;
        RECT 2699.350 603.350 2700.135 603.650 ;
        RECT 2699.550 603.340 2700.135 603.350 ;
        RECT 2699.805 603.335 2700.135 603.340 ;
        RECT 2699.805 579.850 2700.135 579.865 ;
        RECT 2700.470 579.850 2700.850 579.860 ;
        RECT 2699.805 579.550 2700.850 579.850 ;
        RECT 2699.805 579.535 2700.135 579.550 ;
        RECT 2700.470 579.540 2700.850 579.550 ;
        RECT 337.910 469.690 338.290 469.700 ;
        RECT 362.085 469.690 362.415 469.705 ;
        RECT 337.910 469.390 362.415 469.690 ;
        RECT 337.910 469.380 338.290 469.390 ;
        RECT 362.085 469.375 362.415 469.390 ;
        RECT 434.510 469.690 434.890 469.700 ;
        RECT 458.685 469.690 459.015 469.705 ;
        RECT 434.510 469.390 459.015 469.690 ;
        RECT 434.510 469.380 434.890 469.390 ;
        RECT 458.685 469.375 459.015 469.390 ;
        RECT 531.110 469.690 531.490 469.700 ;
        RECT 555.285 469.690 555.615 469.705 ;
        RECT 531.110 469.390 555.615 469.690 ;
        RECT 531.110 469.380 531.490 469.390 ;
        RECT 555.285 469.375 555.615 469.390 ;
        RECT 627.710 469.690 628.090 469.700 ;
        RECT 651.885 469.690 652.215 469.705 ;
        RECT 627.710 469.390 652.215 469.690 ;
        RECT 627.710 469.380 628.090 469.390 ;
        RECT 651.885 469.375 652.215 469.390 ;
        RECT 48.110 469.010 48.490 469.020 ;
        RECT 772.405 469.010 772.735 469.025 ;
        RECT 48.110 468.710 96.290 469.010 ;
        RECT 48.110 468.700 48.490 468.710 ;
        RECT 95.990 467.650 96.290 468.710 ;
        RECT 109.790 468.710 111.010 469.010 ;
        RECT 109.790 467.650 110.090 468.710 ;
        RECT 110.710 468.330 111.010 468.710 ;
        RECT 302.990 468.710 304.210 469.010 ;
        RECT 144.710 468.330 145.090 468.340 ;
        RECT 110.710 468.030 145.090 468.330 ;
        RECT 144.710 468.020 145.090 468.030 ;
        RECT 240.645 468.330 240.975 468.345 ;
        RECT 241.310 468.330 241.690 468.340 ;
        RECT 240.645 468.030 241.690 468.330 ;
        RECT 240.645 468.015 240.975 468.030 ;
        RECT 241.310 468.020 241.690 468.030 ;
        RECT 193.265 467.650 193.595 467.665 ;
        RECT 95.990 467.350 110.090 467.650 ;
        RECT 192.590 467.350 193.595 467.650 ;
        RECT 48.110 466.970 48.490 466.980 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 24.230 466.670 48.490 466.970 ;
        RECT 24.230 466.290 24.530 466.670 ;
        RECT 48.110 466.660 48.490 466.670 ;
        RECT -4.800 465.990 24.530 466.290 ;
        RECT 144.710 466.290 145.090 466.300 ;
        RECT 192.590 466.290 192.890 467.350 ;
        RECT 193.265 467.335 193.595 467.350 ;
        RECT 289.150 467.650 289.530 467.660 ;
        RECT 302.990 467.650 303.290 468.710 ;
        RECT 303.910 468.330 304.210 468.710 ;
        RECT 399.590 468.710 400.810 469.010 ;
        RECT 337.910 468.330 338.290 468.340 ;
        RECT 303.910 468.030 338.290 468.330 ;
        RECT 337.910 468.020 338.290 468.030 ;
        RECT 362.085 468.330 362.415 468.345 ;
        RECT 362.085 468.030 386.090 468.330 ;
        RECT 362.085 468.015 362.415 468.030 ;
        RECT 289.150 467.350 303.290 467.650 ;
        RECT 385.790 467.650 386.090 468.030 ;
        RECT 399.590 467.650 399.890 468.710 ;
        RECT 400.510 468.330 400.810 468.710 ;
        RECT 496.190 468.710 497.410 469.010 ;
        RECT 434.510 468.330 434.890 468.340 ;
        RECT 400.510 468.030 434.890 468.330 ;
        RECT 434.510 468.020 434.890 468.030 ;
        RECT 458.685 468.330 459.015 468.345 ;
        RECT 458.685 468.030 482.690 468.330 ;
        RECT 458.685 468.015 459.015 468.030 ;
        RECT 385.790 467.350 399.890 467.650 ;
        RECT 482.390 467.650 482.690 468.030 ;
        RECT 496.190 467.650 496.490 468.710 ;
        RECT 497.110 468.330 497.410 468.710 ;
        RECT 592.790 468.710 594.010 469.010 ;
        RECT 531.110 468.330 531.490 468.340 ;
        RECT 497.110 468.030 531.490 468.330 ;
        RECT 531.110 468.020 531.490 468.030 ;
        RECT 555.285 468.330 555.615 468.345 ;
        RECT 555.285 468.030 579.290 468.330 ;
        RECT 555.285 468.015 555.615 468.030 ;
        RECT 482.390 467.350 496.490 467.650 ;
        RECT 578.990 467.650 579.290 468.030 ;
        RECT 592.790 467.650 593.090 468.710 ;
        RECT 593.710 468.330 594.010 468.710 ;
        RECT 772.405 468.710 807.450 469.010 ;
        RECT 772.405 468.695 772.735 468.710 ;
        RECT 627.710 468.330 628.090 468.340 ;
        RECT 593.710 468.030 628.090 468.330 ;
        RECT 627.710 468.020 628.090 468.030 ;
        RECT 651.885 468.330 652.215 468.345 ;
        RECT 700.185 468.330 700.515 468.345 ;
        RECT 724.565 468.330 724.895 468.345 ;
        RECT 651.885 468.030 675.890 468.330 ;
        RECT 651.885 468.015 652.215 468.030 ;
        RECT 578.990 467.350 593.090 467.650 ;
        RECT 675.590 467.650 675.890 468.030 ;
        RECT 700.185 468.030 724.895 468.330 ;
        RECT 700.185 468.015 700.515 468.030 ;
        RECT 724.565 468.015 724.895 468.030 ;
        RECT 807.150 467.650 807.450 468.710 ;
        RECT 854.990 468.710 904.050 469.010 ;
        RECT 854.990 467.650 855.290 468.710 ;
        RECT 675.590 467.350 676.810 467.650 ;
        RECT 807.150 467.350 855.290 467.650 ;
        RECT 903.750 467.650 904.050 468.710 ;
        RECT 951.590 468.710 1000.650 469.010 ;
        RECT 951.590 467.650 951.890 468.710 ;
        RECT 903.750 467.350 951.890 467.650 ;
        RECT 1000.350 467.650 1000.650 468.710 ;
        RECT 1048.190 468.710 1097.250 469.010 ;
        RECT 1048.190 467.650 1048.490 468.710 ;
        RECT 1000.350 467.350 1048.490 467.650 ;
        RECT 1096.950 467.650 1097.250 468.710 ;
        RECT 1144.790 468.710 1193.850 469.010 ;
        RECT 1144.790 467.650 1145.090 468.710 ;
        RECT 1096.950 467.350 1145.090 467.650 ;
        RECT 1193.550 467.650 1193.850 468.710 ;
        RECT 1241.390 468.710 1290.450 469.010 ;
        RECT 1241.390 467.650 1241.690 468.710 ;
        RECT 1193.550 467.350 1241.690 467.650 ;
        RECT 1290.150 467.650 1290.450 468.710 ;
        RECT 1337.990 468.710 1387.050 469.010 ;
        RECT 1337.990 467.650 1338.290 468.710 ;
        RECT 1290.150 467.350 1338.290 467.650 ;
        RECT 1386.750 467.650 1387.050 468.710 ;
        RECT 1434.590 468.710 1483.650 469.010 ;
        RECT 1434.590 467.650 1434.890 468.710 ;
        RECT 1386.750 467.350 1434.890 467.650 ;
        RECT 1483.350 467.650 1483.650 468.710 ;
        RECT 1531.190 468.710 1580.250 469.010 ;
        RECT 1531.190 467.650 1531.490 468.710 ;
        RECT 1483.350 467.350 1531.490 467.650 ;
        RECT 1579.950 467.650 1580.250 468.710 ;
        RECT 1627.790 468.710 1676.850 469.010 ;
        RECT 1627.790 467.650 1628.090 468.710 ;
        RECT 1579.950 467.350 1628.090 467.650 ;
        RECT 1676.550 467.650 1676.850 468.710 ;
        RECT 1724.390 468.710 1773.450 469.010 ;
        RECT 1724.390 467.650 1724.690 468.710 ;
        RECT 1676.550 467.350 1724.690 467.650 ;
        RECT 1773.150 467.650 1773.450 468.710 ;
        RECT 1820.990 468.710 1870.050 469.010 ;
        RECT 1820.990 467.650 1821.290 468.710 ;
        RECT 1773.150 467.350 1821.290 467.650 ;
        RECT 1869.750 467.650 1870.050 468.710 ;
        RECT 1917.590 468.710 1966.650 469.010 ;
        RECT 1917.590 467.650 1917.890 468.710 ;
        RECT 1869.750 467.350 1917.890 467.650 ;
        RECT 1966.350 467.650 1966.650 468.710 ;
        RECT 2014.190 468.710 2063.250 469.010 ;
        RECT 2014.190 467.650 2014.490 468.710 ;
        RECT 1966.350 467.350 2014.490 467.650 ;
        RECT 2062.950 467.650 2063.250 468.710 ;
        RECT 2110.790 468.710 2159.850 469.010 ;
        RECT 2110.790 467.650 2111.090 468.710 ;
        RECT 2062.950 467.350 2111.090 467.650 ;
        RECT 2159.550 467.650 2159.850 468.710 ;
        RECT 2207.390 468.710 2256.450 469.010 ;
        RECT 2207.390 467.650 2207.690 468.710 ;
        RECT 2159.550 467.350 2207.690 467.650 ;
        RECT 2256.150 467.650 2256.450 468.710 ;
        RECT 2303.990 468.710 2353.050 469.010 ;
        RECT 2303.990 467.650 2304.290 468.710 ;
        RECT 2256.150 467.350 2304.290 467.650 ;
        RECT 2352.750 467.650 2353.050 468.710 ;
        RECT 2400.590 468.710 2449.650 469.010 ;
        RECT 2400.590 467.650 2400.890 468.710 ;
        RECT 2352.750 467.350 2400.890 467.650 ;
        RECT 2449.350 467.650 2449.650 468.710 ;
        RECT 2497.190 468.710 2546.250 469.010 ;
        RECT 2497.190 467.650 2497.490 468.710 ;
        RECT 2449.350 467.350 2497.490 467.650 ;
        RECT 2545.950 467.650 2546.250 468.710 ;
        RECT 2593.790 468.710 2642.850 469.010 ;
        RECT 2593.790 467.650 2594.090 468.710 ;
        RECT 2545.950 467.350 2594.090 467.650 ;
        RECT 2642.550 467.650 2642.850 468.710 ;
        RECT 2700.470 467.650 2700.850 467.660 ;
        RECT 2642.550 467.350 2700.850 467.650 ;
        RECT 289.150 467.340 289.530 467.350 ;
        RECT 144.710 465.990 192.890 466.290 ;
        RECT 241.310 466.290 241.690 466.300 ;
        RECT 289.150 466.290 289.530 466.300 ;
        RECT 241.310 465.990 289.530 466.290 ;
        RECT 676.510 466.290 676.810 467.350 ;
        RECT 2700.470 467.340 2700.850 467.350 ;
        RECT 700.185 466.290 700.515 466.305 ;
        RECT 676.510 465.990 700.515 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 144.710 465.980 145.090 465.990 ;
        RECT 241.310 465.980 241.690 465.990 ;
        RECT 289.150 465.980 289.530 465.990 ;
        RECT 700.185 465.975 700.515 465.990 ;
      LAYER via3 ;
        RECT 2698.660 2318.300 2698.980 2318.620 ;
        RECT 2698.660 2259.820 2698.980 2260.140 ;
        RECT 2702.340 2259.820 2702.660 2260.140 ;
        RECT 2698.660 2211.540 2698.980 2211.860 ;
        RECT 2702.340 2211.540 2702.660 2211.860 ;
        RECT 2698.660 2163.260 2698.980 2163.580 ;
        RECT 2702.340 2163.260 2702.660 2163.580 ;
        RECT 2698.660 2066.700 2698.980 2067.020 ;
        RECT 2702.340 2066.700 2702.660 2067.020 ;
        RECT 2698.660 2018.420 2698.980 2018.740 ;
        RECT 2702.340 2018.420 2702.660 2018.740 ;
        RECT 2698.660 1904.860 2698.980 1905.180 ;
        RECT 2702.340 1904.860 2702.660 1905.180 ;
        RECT 2698.660 1745.060 2698.980 1745.380 ;
        RECT 2699.580 1655.980 2699.900 1656.300 ;
        RECT 2699.580 1511.820 2699.900 1512.140 ;
        RECT 2700.500 1510.460 2700.820 1510.780 ;
        RECT 2700.500 1459.460 2700.820 1459.780 ;
        RECT 2700.500 1395.540 2700.820 1395.860 ;
        RECT 2700.500 1366.980 2700.820 1367.300 ;
        RECT 2698.660 1324.820 2698.980 1325.140 ;
        RECT 2698.660 1318.020 2698.980 1318.340 ;
        RECT 2699.580 1317.340 2699.900 1317.660 ;
        RECT 2700.500 1080.020 2700.820 1080.340 ;
        RECT 2699.580 1014.740 2699.900 1015.060 ;
        RECT 2699.580 980.060 2699.900 980.380 ;
        RECT 2700.500 978.700 2700.820 979.020 ;
        RECT 2700.500 965.780 2700.820 966.100 ;
        RECT 2699.580 918.180 2699.900 918.500 ;
        RECT 2699.580 883.500 2699.900 883.820 ;
        RECT 2700.500 882.140 2700.820 882.460 ;
        RECT 2700.500 835.220 2700.820 835.540 ;
        RECT 2700.500 820.940 2700.820 821.260 ;
        RECT 2699.580 813.460 2699.900 813.780 ;
        RECT 2700.500 765.860 2700.820 766.180 ;
        RECT 2700.500 738.660 2700.820 738.980 ;
        RECT 2698.660 724.380 2698.980 724.700 ;
        RECT 2699.580 603.340 2699.900 603.660 ;
        RECT 2700.500 579.540 2700.820 579.860 ;
        RECT 337.940 469.380 338.260 469.700 ;
        RECT 434.540 469.380 434.860 469.700 ;
        RECT 531.140 469.380 531.460 469.700 ;
        RECT 627.740 469.380 628.060 469.700 ;
        RECT 48.140 468.700 48.460 469.020 ;
        RECT 144.740 468.020 145.060 468.340 ;
        RECT 241.340 468.020 241.660 468.340 ;
        RECT 48.140 466.660 48.460 466.980 ;
        RECT 144.740 465.980 145.060 466.300 ;
        RECT 289.180 467.340 289.500 467.660 ;
        RECT 337.940 468.020 338.260 468.340 ;
        RECT 434.540 468.020 434.860 468.340 ;
        RECT 531.140 468.020 531.460 468.340 ;
        RECT 627.740 468.020 628.060 468.340 ;
        RECT 241.340 465.980 241.660 466.300 ;
        RECT 289.180 465.980 289.500 466.300 ;
        RECT 2700.500 467.340 2700.820 467.660 ;
      LAYER met4 ;
        RECT 2698.655 2318.295 2698.985 2318.625 ;
        RECT 2698.670 2260.145 2698.970 2318.295 ;
        RECT 2698.655 2259.815 2698.985 2260.145 ;
        RECT 2702.335 2259.815 2702.665 2260.145 ;
        RECT 2702.350 2211.865 2702.650 2259.815 ;
        RECT 2698.655 2211.535 2698.985 2211.865 ;
        RECT 2702.335 2211.535 2702.665 2211.865 ;
        RECT 2698.670 2163.585 2698.970 2211.535 ;
        RECT 2698.655 2163.255 2698.985 2163.585 ;
        RECT 2702.335 2163.255 2702.665 2163.585 ;
        RECT 2702.350 2067.025 2702.650 2163.255 ;
        RECT 2698.655 2066.695 2698.985 2067.025 ;
        RECT 2702.335 2066.695 2702.665 2067.025 ;
        RECT 2698.670 2018.745 2698.970 2066.695 ;
        RECT 2698.655 2018.415 2698.985 2018.745 ;
        RECT 2702.335 2018.415 2702.665 2018.745 ;
        RECT 2702.350 1905.185 2702.650 2018.415 ;
        RECT 2698.655 1904.855 2698.985 1905.185 ;
        RECT 2702.335 1904.855 2702.665 1905.185 ;
        RECT 2698.670 1895.650 2698.970 1904.855 ;
        RECT 2698.670 1895.350 2699.890 1895.650 ;
        RECT 2699.590 1817.450 2699.890 1895.350 ;
        RECT 2698.670 1817.150 2699.890 1817.450 ;
        RECT 2698.670 1745.385 2698.970 1817.150 ;
        RECT 2698.655 1745.055 2698.985 1745.385 ;
        RECT 2699.575 1655.975 2699.905 1656.305 ;
        RECT 2699.590 1603.250 2699.890 1655.975 ;
        RECT 2699.590 1602.950 2700.810 1603.250 ;
        RECT 2700.510 1572.650 2700.810 1602.950 ;
        RECT 2699.590 1572.350 2700.810 1572.650 ;
        RECT 2699.590 1512.145 2699.890 1572.350 ;
        RECT 2699.575 1511.815 2699.905 1512.145 ;
        RECT 2700.495 1510.455 2700.825 1510.785 ;
        RECT 2700.510 1459.785 2700.810 1510.455 ;
        RECT 2700.495 1459.455 2700.825 1459.785 ;
        RECT 2700.495 1395.535 2700.825 1395.865 ;
        RECT 2700.510 1367.305 2700.810 1395.535 ;
        RECT 2700.495 1366.975 2700.825 1367.305 ;
        RECT 2698.655 1324.815 2698.985 1325.145 ;
        RECT 2698.670 1318.345 2698.970 1324.815 ;
        RECT 2698.655 1318.015 2698.985 1318.345 ;
        RECT 2699.575 1317.335 2699.905 1317.665 ;
        RECT 2699.590 1283.650 2699.890 1317.335 ;
        RECT 2699.590 1283.350 2700.810 1283.650 ;
        RECT 2700.510 1080.345 2700.810 1283.350 ;
        RECT 2700.495 1080.015 2700.825 1080.345 ;
        RECT 2699.575 1014.735 2699.905 1015.065 ;
        RECT 2699.590 980.385 2699.890 1014.735 ;
        RECT 2699.575 980.055 2699.905 980.385 ;
        RECT 2700.495 978.695 2700.825 979.025 ;
        RECT 2700.510 966.105 2700.810 978.695 ;
        RECT 2700.495 965.775 2700.825 966.105 ;
        RECT 2699.575 918.175 2699.905 918.505 ;
        RECT 2699.590 883.825 2699.890 918.175 ;
        RECT 2699.575 883.495 2699.905 883.825 ;
        RECT 2700.495 882.135 2700.825 882.465 ;
        RECT 2700.510 835.545 2700.810 882.135 ;
        RECT 2700.495 835.215 2700.825 835.545 ;
        RECT 2700.495 821.250 2700.825 821.265 ;
        RECT 2699.590 820.950 2700.825 821.250 ;
        RECT 2699.590 813.785 2699.890 820.950 ;
        RECT 2700.495 820.935 2700.825 820.950 ;
        RECT 2699.575 813.455 2699.905 813.785 ;
        RECT 2700.495 765.855 2700.825 766.185 ;
        RECT 2700.510 738.985 2700.810 765.855 ;
        RECT 2700.495 738.655 2700.825 738.985 ;
        RECT 2698.655 724.375 2698.985 724.705 ;
        RECT 2698.670 688.650 2698.970 724.375 ;
        RECT 2698.670 688.350 2700.810 688.650 ;
        RECT 2700.510 641.050 2700.810 688.350 ;
        RECT 2699.590 640.750 2700.810 641.050 ;
        RECT 2699.590 603.665 2699.890 640.750 ;
        RECT 2699.575 603.335 2699.905 603.665 ;
        RECT 2700.495 579.535 2700.825 579.865 ;
        RECT 337.935 469.375 338.265 469.705 ;
        RECT 434.535 469.375 434.865 469.705 ;
        RECT 531.135 469.375 531.465 469.705 ;
        RECT 627.735 469.375 628.065 469.705 ;
        RECT 48.135 468.695 48.465 469.025 ;
        RECT 48.150 466.985 48.450 468.695 ;
        RECT 337.950 468.345 338.250 469.375 ;
        RECT 434.550 468.345 434.850 469.375 ;
        RECT 531.150 468.345 531.450 469.375 ;
        RECT 627.750 468.345 628.050 469.375 ;
        RECT 144.735 468.015 145.065 468.345 ;
        RECT 241.335 468.015 241.665 468.345 ;
        RECT 337.935 468.015 338.265 468.345 ;
        RECT 434.535 468.015 434.865 468.345 ;
        RECT 531.135 468.015 531.465 468.345 ;
        RECT 627.735 468.015 628.065 468.345 ;
        RECT 48.135 466.655 48.465 466.985 ;
        RECT 144.750 466.305 145.050 468.015 ;
        RECT 241.350 466.305 241.650 468.015 ;
        RECT 2700.510 467.665 2700.810 579.535 ;
        RECT 289.175 467.335 289.505 467.665 ;
        RECT 2700.495 467.335 2700.825 467.665 ;
        RECT 289.190 466.305 289.490 467.335 ;
        RECT 144.735 465.975 145.065 466.305 ;
        RECT 241.335 465.975 241.665 466.305 ;
        RECT 289.175 465.975 289.505 466.305 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2703.030 2067.780 2703.350 2067.840 ;
        RECT 2703.950 2067.780 2704.270 2067.840 ;
        RECT 2703.030 2067.640 2704.270 2067.780 ;
        RECT 2703.030 2067.580 2703.350 2067.640 ;
        RECT 2703.950 2067.580 2704.270 2067.640 ;
      LAYER via ;
        RECT 2703.060 2067.580 2703.320 2067.840 ;
        RECT 2703.980 2067.580 2704.240 2067.840 ;
      LAYER met2 ;
        RECT 2703.970 2091.835 2704.250 2092.205 ;
        RECT 2704.040 2067.870 2704.180 2091.835 ;
        RECT 2703.060 2067.550 2703.320 2067.870 ;
        RECT 2703.980 2067.550 2704.240 2067.870 ;
        RECT 2703.120 2025.450 2703.260 2067.550 ;
        RECT 2702.660 2025.310 2703.260 2025.450 ;
        RECT 2702.660 1992.925 2702.800 2025.310 ;
        RECT 2702.590 1992.555 2702.870 1992.925 ;
        RECT 16.650 254.475 16.930 254.845 ;
        RECT 16.720 250.765 16.860 254.475 ;
        RECT 16.650 250.395 16.930 250.765 ;
      LAYER via2 ;
        RECT 2703.970 2091.880 2704.250 2092.160 ;
        RECT 2702.590 1992.600 2702.870 1992.880 ;
        RECT 16.650 254.520 16.930 254.800 ;
        RECT 16.650 250.440 16.930 250.720 ;
      LAYER met3 ;
        RECT 2696.000 2351.960 2700.000 2352.560 ;
        RECT 2697.750 2349.900 2698.050 2351.960 ;
        RECT 2697.710 2349.580 2698.090 2349.900 ;
        RECT 2697.710 2092.170 2698.090 2092.180 ;
        RECT 2703.945 2092.170 2704.275 2092.185 ;
        RECT 2697.710 2091.870 2704.275 2092.170 ;
        RECT 2697.710 2091.860 2698.090 2091.870 ;
        RECT 2703.945 2091.855 2704.275 2091.870 ;
        RECT 2697.710 1992.890 2698.090 1992.900 ;
        RECT 2702.565 1992.890 2702.895 1992.905 ;
        RECT 2697.710 1992.590 2702.895 1992.890 ;
        RECT 2697.710 1992.580 2698.090 1992.590 ;
        RECT 2702.565 1992.575 2702.895 1992.590 ;
        RECT 2697.710 1797.420 2698.090 1797.740 ;
        RECT 2697.750 1797.060 2698.050 1797.420 ;
        RECT 2697.710 1796.740 2698.090 1797.060 ;
        RECT 16.625 254.810 16.955 254.825 ;
        RECT 2697.710 254.810 2698.090 254.820 ;
        RECT 16.625 254.510 2698.090 254.810 ;
        RECT 16.625 254.495 16.955 254.510 ;
        RECT 2697.710 254.500 2698.090 254.510 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 16.625 250.730 16.955 250.745 ;
        RECT -4.800 250.430 16.955 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 16.625 250.415 16.955 250.430 ;
      LAYER via3 ;
        RECT 2697.740 2349.580 2698.060 2349.900 ;
        RECT 2697.740 2091.860 2698.060 2092.180 ;
        RECT 2697.740 1992.580 2698.060 1992.900 ;
        RECT 2697.740 1797.420 2698.060 1797.740 ;
        RECT 2697.740 1796.740 2698.060 1797.060 ;
        RECT 2697.740 254.500 2698.060 254.820 ;
      LAYER met4 ;
        RECT 2697.735 2349.575 2698.065 2349.905 ;
        RECT 2697.750 2092.185 2698.050 2349.575 ;
        RECT 2697.735 2091.855 2698.065 2092.185 ;
        RECT 2697.735 1992.575 2698.065 1992.905 ;
        RECT 2697.750 1797.745 2698.050 1992.575 ;
        RECT 2697.735 1797.415 2698.065 1797.745 ;
        RECT 2697.735 1796.735 2698.065 1797.065 ;
        RECT 2697.750 254.825 2698.050 1796.735 ;
        RECT 2697.735 254.495 2698.065 254.825 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.110 40.955 17.390 41.325 ;
        RECT 17.180 35.885 17.320 40.955 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 41.000 17.390 41.280 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT 2711.510 2384.570 2711.890 2384.580 ;
        RECT 2699.740 2384.520 2711.890 2384.570 ;
        RECT 2696.000 2384.270 2711.890 2384.520 ;
        RECT 2696.000 2383.920 2700.000 2384.270 ;
        RECT 2711.510 2384.260 2711.890 2384.270 ;
        RECT 17.085 41.290 17.415 41.305 ;
        RECT 2711.510 41.290 2711.890 41.300 ;
        RECT 17.085 40.990 2711.890 41.290 ;
        RECT 17.085 40.975 17.415 40.990 ;
        RECT 2711.510 40.980 2711.890 40.990 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
      LAYER via3 ;
        RECT 2711.540 2384.260 2711.860 2384.580 ;
        RECT 2711.540 40.980 2711.860 41.300 ;
      LAYER met4 ;
        RECT 2711.535 2384.255 2711.865 2384.585 ;
        RECT 2711.550 41.305 2711.850 2384.255 ;
        RECT 2711.535 40.975 2711.865 41.305 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2716.370 910.760 2716.690 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 2716.370 910.620 2901.150 910.760 ;
        RECT 2716.370 910.560 2716.690 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 2716.400 910.560 2716.660 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 2716.390 1309.835 2716.670 1310.205 ;
        RECT 2716.460 910.850 2716.600 1309.835 ;
        RECT 2716.400 910.530 2716.660 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2716.390 1309.880 2716.670 1310.160 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2716.365 1310.170 2716.695 1310.185 ;
        RECT 2699.740 1310.120 2716.695 1310.170 ;
        RECT 2696.000 1309.870 2716.695 1310.120 ;
        RECT 2696.000 1309.520 2700.000 1309.870 ;
        RECT 2716.365 1309.855 2716.695 1309.870 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2717.750 1145.360 2718.070 1145.420 ;
        RECT 2900.830 1145.360 2901.150 1145.420 ;
        RECT 2717.750 1145.220 2901.150 1145.360 ;
        RECT 2717.750 1145.160 2718.070 1145.220 ;
        RECT 2900.830 1145.160 2901.150 1145.220 ;
      LAYER via ;
        RECT 2717.780 1145.160 2718.040 1145.420 ;
        RECT 2900.860 1145.160 2901.120 1145.420 ;
      LAYER met2 ;
        RECT 2717.770 1341.795 2718.050 1342.165 ;
        RECT 2717.840 1145.450 2717.980 1341.795 ;
        RECT 2717.780 1145.130 2718.040 1145.450 ;
        RECT 2900.860 1145.130 2901.120 1145.450 ;
        RECT 2900.920 1144.285 2901.060 1145.130 ;
        RECT 2900.850 1143.915 2901.130 1144.285 ;
      LAYER via2 ;
        RECT 2717.770 1341.840 2718.050 1342.120 ;
        RECT 2900.850 1143.960 2901.130 1144.240 ;
      LAYER met3 ;
        RECT 2717.745 1342.130 2718.075 1342.145 ;
        RECT 2699.740 1342.080 2718.075 1342.130 ;
        RECT 2696.000 1341.830 2718.075 1342.080 ;
        RECT 2696.000 1341.480 2700.000 1341.830 ;
        RECT 2717.745 1341.815 2718.075 1341.830 ;
        RECT 2900.825 1144.250 2901.155 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2900.825 1143.950 2924.800 1144.250 ;
        RECT 2900.825 1143.935 2901.155 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1376.560 2713.470 1376.620 ;
        RECT 2900.830 1376.560 2901.150 1376.620 ;
        RECT 2713.150 1376.420 2901.150 1376.560 ;
        RECT 2713.150 1376.360 2713.470 1376.420 ;
        RECT 2900.830 1376.360 2901.150 1376.420 ;
      LAYER via ;
        RECT 2713.180 1376.360 2713.440 1376.620 ;
        RECT 2900.860 1376.360 2901.120 1376.620 ;
      LAYER met2 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
        RECT 2900.920 1376.650 2901.060 1378.515 ;
        RECT 2713.180 1376.330 2713.440 1376.650 ;
        RECT 2900.860 1376.330 2901.120 1376.650 ;
        RECT 2713.240 1373.445 2713.380 1376.330 ;
        RECT 2713.170 1373.075 2713.450 1373.445 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
        RECT 2713.170 1373.120 2713.450 1373.400 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
        RECT 2713.145 1373.410 2713.475 1373.425 ;
        RECT 2699.740 1373.360 2713.475 1373.410 ;
        RECT 2696.000 1373.110 2713.475 1373.360 ;
        RECT 2696.000 1372.760 2700.000 1373.110 ;
        RECT 2713.145 1373.095 2713.475 1373.110 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1407.500 2713.470 1407.560 ;
        RECT 2902.670 1407.500 2902.990 1407.560 ;
        RECT 2713.150 1407.360 2902.990 1407.500 ;
        RECT 2713.150 1407.300 2713.470 1407.360 ;
        RECT 2902.670 1407.300 2902.990 1407.360 ;
      LAYER via ;
        RECT 2713.180 1407.300 2713.440 1407.560 ;
        RECT 2902.700 1407.300 2902.960 1407.560 ;
      LAYER met2 ;
        RECT 2902.690 1613.115 2902.970 1613.485 ;
        RECT 2902.760 1407.590 2902.900 1613.115 ;
        RECT 2713.180 1407.270 2713.440 1407.590 ;
        RECT 2902.700 1407.270 2902.960 1407.590 ;
        RECT 2713.240 1405.405 2713.380 1407.270 ;
        RECT 2713.170 1405.035 2713.450 1405.405 ;
      LAYER via2 ;
        RECT 2902.690 1613.160 2902.970 1613.440 ;
        RECT 2713.170 1405.080 2713.450 1405.360 ;
      LAYER met3 ;
        RECT 2902.665 1613.450 2902.995 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2902.665 1613.150 2924.800 1613.450 ;
        RECT 2902.665 1613.135 2902.995 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2713.145 1405.370 2713.475 1405.385 ;
        RECT 2699.740 1405.320 2713.475 1405.370 ;
        RECT 2696.000 1405.070 2713.475 1405.320 ;
        RECT 2696.000 1404.720 2700.000 1405.070 ;
        RECT 2713.145 1405.055 2713.475 1405.070 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1441.840 2713.470 1441.900 ;
        RECT 2901.290 1441.840 2901.610 1441.900 ;
        RECT 2713.150 1441.700 2901.610 1441.840 ;
        RECT 2713.150 1441.640 2713.470 1441.700 ;
        RECT 2901.290 1441.640 2901.610 1441.700 ;
      LAYER via ;
        RECT 2713.180 1441.640 2713.440 1441.900 ;
        RECT 2901.320 1441.640 2901.580 1441.900 ;
      LAYER met2 ;
        RECT 2901.310 1847.715 2901.590 1848.085 ;
        RECT 2901.380 1441.930 2901.520 1847.715 ;
        RECT 2713.180 1441.610 2713.440 1441.930 ;
        RECT 2901.320 1441.610 2901.580 1441.930 ;
        RECT 2713.240 1436.685 2713.380 1441.610 ;
        RECT 2713.170 1436.315 2713.450 1436.685 ;
      LAYER via2 ;
        RECT 2901.310 1847.760 2901.590 1848.040 ;
        RECT 2713.170 1436.360 2713.450 1436.640 ;
      LAYER met3 ;
        RECT 2901.285 1848.050 2901.615 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2901.285 1847.750 2924.800 1848.050 ;
        RECT 2901.285 1847.735 2901.615 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
        RECT 2713.145 1436.650 2713.475 1436.665 ;
        RECT 2699.740 1436.600 2713.475 1436.650 ;
        RECT 2696.000 1436.350 2713.475 1436.600 ;
        RECT 2696.000 1436.000 2700.000 1436.350 ;
        RECT 2713.145 1436.335 2713.475 1436.350 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2825.850 2077.300 2826.170 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 2825.850 2077.160 2901.150 2077.300 ;
        RECT 2825.850 2077.100 2826.170 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
        RECT 2713.150 1469.720 2713.470 1469.780 ;
        RECT 2825.850 1469.720 2826.170 1469.780 ;
        RECT 2713.150 1469.580 2826.170 1469.720 ;
        RECT 2713.150 1469.520 2713.470 1469.580 ;
        RECT 2825.850 1469.520 2826.170 1469.580 ;
      LAYER via ;
        RECT 2825.880 2077.100 2826.140 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
        RECT 2713.180 1469.520 2713.440 1469.780 ;
        RECT 2825.880 1469.520 2826.140 1469.780 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 2825.880 2077.070 2826.140 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 2825.940 1469.810 2826.080 2077.070 ;
        RECT 2713.180 1469.490 2713.440 1469.810 ;
        RECT 2825.880 1469.490 2826.140 1469.810 ;
        RECT 2713.240 1468.645 2713.380 1469.490 ;
        RECT 2713.170 1468.275 2713.450 1468.645 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
        RECT 2713.170 1468.320 2713.450 1468.600 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
        RECT 2713.145 1468.610 2713.475 1468.625 ;
        RECT 2699.740 1468.560 2713.475 1468.610 ;
        RECT 2696.000 1468.310 2713.475 1468.560 ;
        RECT 2696.000 1467.960 2700.000 1468.310 ;
        RECT 2713.145 1468.295 2713.475 1468.310 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2839.190 2311.900 2839.510 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 2839.190 2311.760 2901.150 2311.900 ;
        RECT 2839.190 2311.700 2839.510 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 2713.150 1504.060 2713.470 1504.120 ;
        RECT 2839.190 1504.060 2839.510 1504.120 ;
        RECT 2713.150 1503.920 2839.510 1504.060 ;
        RECT 2713.150 1503.860 2713.470 1503.920 ;
        RECT 2839.190 1503.860 2839.510 1503.920 ;
      LAYER via ;
        RECT 2839.220 2311.700 2839.480 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 2713.180 1503.860 2713.440 1504.120 ;
        RECT 2839.220 1503.860 2839.480 1504.120 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 2839.220 2311.670 2839.480 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 2839.280 1504.150 2839.420 2311.670 ;
        RECT 2713.180 1503.830 2713.440 1504.150 ;
        RECT 2839.220 1503.830 2839.480 1504.150 ;
        RECT 2713.240 1499.925 2713.380 1503.830 ;
        RECT 2713.170 1499.555 2713.450 1499.925 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
        RECT 2713.170 1499.600 2713.450 1499.880 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
        RECT 2713.145 1499.890 2713.475 1499.905 ;
        RECT 2699.740 1499.840 2713.475 1499.890 ;
        RECT 2696.000 1499.590 2713.475 1499.840 ;
        RECT 2696.000 1499.240 2700.000 1499.590 ;
        RECT 2713.145 1499.575 2713.475 1499.590 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2710.850 1173.240 2711.170 1173.300 ;
        RECT 2714.070 1173.240 2714.390 1173.300 ;
        RECT 2710.850 1173.100 2714.390 1173.240 ;
        RECT 2710.850 1173.040 2711.170 1173.100 ;
        RECT 2714.070 1173.040 2714.390 1173.100 ;
        RECT 2713.150 1158.960 2713.470 1159.020 ;
        RECT 2714.070 1158.960 2714.390 1159.020 ;
        RECT 2713.150 1158.820 2714.390 1158.960 ;
        RECT 2713.150 1158.760 2713.470 1158.820 ;
        RECT 2714.070 1158.760 2714.390 1158.820 ;
        RECT 2713.150 1111.020 2713.470 1111.080 ;
        RECT 2714.530 1111.020 2714.850 1111.080 ;
        RECT 2713.150 1110.880 2714.850 1111.020 ;
        RECT 2713.150 1110.820 2713.470 1110.880 ;
        RECT 2714.530 1110.820 2714.850 1110.880 ;
        RECT 2714.530 1077.020 2714.850 1077.080 ;
        RECT 2714.160 1076.880 2714.850 1077.020 ;
        RECT 2714.160 1076.400 2714.300 1076.880 ;
        RECT 2714.530 1076.820 2714.850 1076.880 ;
        RECT 2714.070 1076.140 2714.390 1076.400 ;
        RECT 2713.610 1062.400 2713.930 1062.460 ;
        RECT 2714.070 1062.400 2714.390 1062.460 ;
        RECT 2713.610 1062.260 2714.390 1062.400 ;
        RECT 2713.610 1062.200 2713.930 1062.260 ;
        RECT 2714.070 1062.200 2714.390 1062.260 ;
        RECT 2713.610 1014.460 2713.930 1014.520 ;
        RECT 2714.530 1014.460 2714.850 1014.520 ;
        RECT 2713.610 1014.320 2714.850 1014.460 ;
        RECT 2713.610 1014.260 2713.930 1014.320 ;
        RECT 2714.530 1014.260 2714.850 1014.320 ;
        RECT 2714.530 980.460 2714.850 980.520 ;
        RECT 2714.160 980.320 2714.850 980.460 ;
        RECT 2714.160 979.840 2714.300 980.320 ;
        RECT 2714.530 980.260 2714.850 980.320 ;
        RECT 2714.070 979.580 2714.390 979.840 ;
        RECT 2714.070 869.620 2714.390 869.680 ;
        RECT 2714.990 869.620 2715.310 869.680 ;
        RECT 2714.070 869.480 2715.310 869.620 ;
        RECT 2714.070 869.420 2714.390 869.480 ;
        RECT 2714.990 869.420 2715.310 869.480 ;
        RECT 2714.070 814.200 2714.390 814.260 ;
        RECT 2714.990 814.200 2715.310 814.260 ;
        RECT 2714.070 814.060 2715.310 814.200 ;
        RECT 2714.070 814.000 2714.390 814.060 ;
        RECT 2714.990 814.000 2715.310 814.060 ;
        RECT 2714.070 766.260 2714.390 766.320 ;
        RECT 2714.990 766.260 2715.310 766.320 ;
        RECT 2714.070 766.120 2715.310 766.260 ;
        RECT 2714.070 766.060 2714.390 766.120 ;
        RECT 2714.990 766.060 2715.310 766.120 ;
        RECT 2714.990 717.640 2715.310 717.700 ;
        RECT 2715.910 717.640 2716.230 717.700 ;
        RECT 2714.990 717.500 2716.230 717.640 ;
        RECT 2714.990 717.440 2715.310 717.500 ;
        RECT 2715.910 717.440 2716.230 717.500 ;
        RECT 2714.990 669.700 2715.310 669.760 ;
        RECT 2715.910 669.700 2716.230 669.760 ;
        RECT 2714.990 669.560 2716.230 669.700 ;
        RECT 2714.990 669.500 2715.310 669.560 ;
        RECT 2715.910 669.500 2716.230 669.560 ;
        RECT 2714.990 620.740 2715.310 620.800 ;
        RECT 2716.830 620.740 2717.150 620.800 ;
        RECT 2714.990 620.600 2717.150 620.740 ;
        RECT 2714.990 620.540 2715.310 620.600 ;
        RECT 2716.830 620.540 2717.150 620.600 ;
        RECT 2714.990 496.980 2715.310 497.040 ;
        RECT 2715.910 496.980 2716.230 497.040 ;
        RECT 2714.990 496.840 2716.230 496.980 ;
        RECT 2714.990 496.780 2715.310 496.840 ;
        RECT 2715.910 496.780 2716.230 496.840 ;
        RECT 2714.070 483.040 2714.390 483.100 ;
        RECT 2714.530 483.040 2714.850 483.100 ;
        RECT 2714.070 482.900 2714.850 483.040 ;
        RECT 2714.070 482.840 2714.390 482.900 ;
        RECT 2714.530 482.840 2714.850 482.900 ;
        RECT 2714.070 448.500 2714.390 448.760 ;
        RECT 2714.160 448.360 2714.300 448.500 ;
        RECT 2714.530 448.360 2714.850 448.420 ;
        RECT 2714.160 448.220 2714.850 448.360 ;
        RECT 2714.530 448.160 2714.850 448.220 ;
        RECT 2714.070 434.760 2714.390 434.820 ;
        RECT 2716.370 434.760 2716.690 434.820 ;
        RECT 2714.070 434.620 2716.690 434.760 ;
        RECT 2714.070 434.560 2714.390 434.620 ;
        RECT 2716.370 434.560 2716.690 434.620 ;
        RECT 2714.530 338.200 2714.850 338.260 ;
        RECT 2715.450 338.200 2715.770 338.260 ;
        RECT 2714.530 338.060 2715.770 338.200 ;
        RECT 2714.530 338.000 2714.850 338.060 ;
        RECT 2715.450 338.000 2715.770 338.060 ;
        RECT 2715.450 303.860 2715.770 303.920 ;
        RECT 2714.160 303.720 2715.770 303.860 ;
        RECT 2714.160 303.580 2714.300 303.720 ;
        RECT 2715.450 303.660 2715.770 303.720 ;
        RECT 2714.070 303.320 2714.390 303.580 ;
        RECT 2714.070 255.240 2714.390 255.300 ;
        RECT 2714.990 255.240 2715.310 255.300 ;
        RECT 2714.070 255.100 2715.310 255.240 ;
        RECT 2714.070 255.040 2714.390 255.100 ;
        RECT 2714.990 255.040 2715.310 255.100 ;
        RECT 2714.990 241.300 2715.310 241.360 ;
        RECT 2716.370 241.300 2716.690 241.360 ;
        RECT 2714.990 241.160 2716.690 241.300 ;
        RECT 2714.990 241.100 2715.310 241.160 ;
        RECT 2716.370 241.100 2716.690 241.160 ;
        RECT 2715.450 193.360 2715.770 193.420 ;
        RECT 2716.370 193.360 2716.690 193.420 ;
        RECT 2715.450 193.220 2716.690 193.360 ;
        RECT 2715.450 193.160 2715.770 193.220 ;
        RECT 2716.370 193.160 2716.690 193.220 ;
        RECT 2715.450 151.540 2715.770 151.600 ;
        RECT 2900.830 151.540 2901.150 151.600 ;
        RECT 2715.450 151.400 2901.150 151.540 ;
        RECT 2715.450 151.340 2715.770 151.400 ;
        RECT 2900.830 151.340 2901.150 151.400 ;
      LAYER via ;
        RECT 2710.880 1173.040 2711.140 1173.300 ;
        RECT 2714.100 1173.040 2714.360 1173.300 ;
        RECT 2713.180 1158.760 2713.440 1159.020 ;
        RECT 2714.100 1158.760 2714.360 1159.020 ;
        RECT 2713.180 1110.820 2713.440 1111.080 ;
        RECT 2714.560 1110.820 2714.820 1111.080 ;
        RECT 2714.560 1076.820 2714.820 1077.080 ;
        RECT 2714.100 1076.140 2714.360 1076.400 ;
        RECT 2713.640 1062.200 2713.900 1062.460 ;
        RECT 2714.100 1062.200 2714.360 1062.460 ;
        RECT 2713.640 1014.260 2713.900 1014.520 ;
        RECT 2714.560 1014.260 2714.820 1014.520 ;
        RECT 2714.560 980.260 2714.820 980.520 ;
        RECT 2714.100 979.580 2714.360 979.840 ;
        RECT 2714.100 869.420 2714.360 869.680 ;
        RECT 2715.020 869.420 2715.280 869.680 ;
        RECT 2714.100 814.000 2714.360 814.260 ;
        RECT 2715.020 814.000 2715.280 814.260 ;
        RECT 2714.100 766.060 2714.360 766.320 ;
        RECT 2715.020 766.060 2715.280 766.320 ;
        RECT 2715.020 717.440 2715.280 717.700 ;
        RECT 2715.940 717.440 2716.200 717.700 ;
        RECT 2715.020 669.500 2715.280 669.760 ;
        RECT 2715.940 669.500 2716.200 669.760 ;
        RECT 2715.020 620.540 2715.280 620.800 ;
        RECT 2716.860 620.540 2717.120 620.800 ;
        RECT 2715.020 496.780 2715.280 497.040 ;
        RECT 2715.940 496.780 2716.200 497.040 ;
        RECT 2714.100 482.840 2714.360 483.100 ;
        RECT 2714.560 482.840 2714.820 483.100 ;
        RECT 2714.100 448.500 2714.360 448.760 ;
        RECT 2714.560 448.160 2714.820 448.420 ;
        RECT 2714.100 434.560 2714.360 434.820 ;
        RECT 2716.400 434.560 2716.660 434.820 ;
        RECT 2714.560 338.000 2714.820 338.260 ;
        RECT 2715.480 338.000 2715.740 338.260 ;
        RECT 2715.480 303.660 2715.740 303.920 ;
        RECT 2714.100 303.320 2714.360 303.580 ;
        RECT 2714.100 255.040 2714.360 255.300 ;
        RECT 2715.020 255.040 2715.280 255.300 ;
        RECT 2715.020 241.100 2715.280 241.360 ;
        RECT 2716.400 241.100 2716.660 241.360 ;
        RECT 2715.480 193.160 2715.740 193.420 ;
        RECT 2716.400 193.160 2716.660 193.420 ;
        RECT 2715.480 151.340 2715.740 151.600 ;
        RECT 2900.860 151.340 2901.120 151.600 ;
      LAYER met2 ;
        RECT 2714.550 1225.515 2714.830 1225.885 ;
        RECT 2714.620 1207.525 2714.760 1225.515 ;
        RECT 2710.870 1207.155 2711.150 1207.525 ;
        RECT 2714.550 1207.155 2714.830 1207.525 ;
        RECT 2710.940 1173.330 2711.080 1207.155 ;
        RECT 2710.880 1173.010 2711.140 1173.330 ;
        RECT 2714.100 1173.010 2714.360 1173.330 ;
        RECT 2714.160 1159.050 2714.300 1173.010 ;
        RECT 2713.180 1158.730 2713.440 1159.050 ;
        RECT 2714.100 1158.730 2714.360 1159.050 ;
        RECT 2713.240 1111.110 2713.380 1158.730 ;
        RECT 2713.180 1110.790 2713.440 1111.110 ;
        RECT 2714.560 1110.790 2714.820 1111.110 ;
        RECT 2714.620 1077.110 2714.760 1110.790 ;
        RECT 2714.560 1076.790 2714.820 1077.110 ;
        RECT 2714.100 1076.110 2714.360 1076.430 ;
        RECT 2714.160 1062.490 2714.300 1076.110 ;
        RECT 2713.640 1062.170 2713.900 1062.490 ;
        RECT 2714.100 1062.170 2714.360 1062.490 ;
        RECT 2713.700 1014.550 2713.840 1062.170 ;
        RECT 2713.640 1014.230 2713.900 1014.550 ;
        RECT 2714.560 1014.230 2714.820 1014.550 ;
        RECT 2714.620 980.550 2714.760 1014.230 ;
        RECT 2714.560 980.230 2714.820 980.550 ;
        RECT 2714.100 979.550 2714.360 979.870 ;
        RECT 2714.160 931.330 2714.300 979.550 ;
        RECT 2714.160 931.190 2714.760 931.330 ;
        RECT 2714.620 893.930 2714.760 931.190 ;
        RECT 2714.160 893.790 2714.760 893.930 ;
        RECT 2714.160 869.710 2714.300 893.790 ;
        RECT 2714.100 869.390 2714.360 869.710 ;
        RECT 2715.020 869.565 2715.280 869.710 ;
        RECT 2715.010 869.195 2715.290 869.565 ;
        RECT 2715.010 820.915 2715.290 821.285 ;
        RECT 2715.080 814.290 2715.220 820.915 ;
        RECT 2714.100 813.970 2714.360 814.290 ;
        RECT 2715.020 813.970 2715.280 814.290 ;
        RECT 2714.160 766.350 2714.300 813.970 ;
        RECT 2714.100 766.030 2714.360 766.350 ;
        RECT 2715.020 766.030 2715.280 766.350 ;
        RECT 2715.080 717.730 2715.220 766.030 ;
        RECT 2715.020 717.410 2715.280 717.730 ;
        RECT 2715.940 717.410 2716.200 717.730 ;
        RECT 2716.000 669.790 2716.140 717.410 ;
        RECT 2715.020 669.470 2715.280 669.790 ;
        RECT 2715.940 669.470 2716.200 669.790 ;
        RECT 2715.080 620.830 2715.220 669.470 ;
        RECT 2715.020 620.510 2715.280 620.830 ;
        RECT 2716.860 620.510 2717.120 620.830 ;
        RECT 2716.920 531.605 2717.060 620.510 ;
        RECT 2715.930 531.235 2716.210 531.605 ;
        RECT 2716.850 531.235 2717.130 531.605 ;
        RECT 2715.080 497.070 2715.220 497.225 ;
        RECT 2716.000 497.070 2716.140 531.235 ;
        RECT 2715.020 496.810 2715.280 497.070 ;
        RECT 2714.620 496.750 2715.280 496.810 ;
        RECT 2715.940 496.750 2716.200 497.070 ;
        RECT 2714.620 496.670 2715.220 496.750 ;
        RECT 2714.620 483.130 2714.760 496.670 ;
        RECT 2714.100 482.810 2714.360 483.130 ;
        RECT 2714.560 482.810 2714.820 483.130 ;
        RECT 2714.160 448.790 2714.300 482.810 ;
        RECT 2714.100 448.470 2714.360 448.790 ;
        RECT 2714.560 448.130 2714.820 448.450 ;
        RECT 2714.620 434.930 2714.760 448.130 ;
        RECT 2714.160 434.850 2714.760 434.930 ;
        RECT 2714.100 434.790 2714.760 434.850 ;
        RECT 2714.100 434.530 2714.360 434.790 ;
        RECT 2716.400 434.530 2716.660 434.850 ;
        RECT 2716.460 386.650 2716.600 434.530 ;
        RECT 2716.000 386.510 2716.600 386.650 ;
        RECT 2716.000 386.085 2716.140 386.510 ;
        RECT 2714.550 385.715 2714.830 386.085 ;
        RECT 2715.930 385.715 2716.210 386.085 ;
        RECT 2714.620 338.290 2714.760 385.715 ;
        RECT 2714.560 337.970 2714.820 338.290 ;
        RECT 2715.480 337.970 2715.740 338.290 ;
        RECT 2715.540 303.950 2715.680 337.970 ;
        RECT 2715.480 303.630 2715.740 303.950 ;
        RECT 2714.100 303.290 2714.360 303.610 ;
        RECT 2714.160 255.330 2714.300 303.290 ;
        RECT 2714.100 255.010 2714.360 255.330 ;
        RECT 2715.020 255.010 2715.280 255.330 ;
        RECT 2715.080 241.390 2715.220 255.010 ;
        RECT 2715.020 241.070 2715.280 241.390 ;
        RECT 2716.400 241.070 2716.660 241.390 ;
        RECT 2716.460 193.450 2716.600 241.070 ;
        RECT 2715.480 193.130 2715.740 193.450 ;
        RECT 2716.400 193.130 2716.660 193.450 ;
        RECT 2715.540 151.630 2715.680 193.130 ;
        RECT 2715.480 151.310 2715.740 151.630 ;
        RECT 2900.860 151.310 2901.120 151.630 ;
        RECT 2900.920 146.725 2901.060 151.310 ;
        RECT 2900.850 146.355 2901.130 146.725 ;
      LAYER via2 ;
        RECT 2714.550 1225.560 2714.830 1225.840 ;
        RECT 2710.870 1207.200 2711.150 1207.480 ;
        RECT 2714.550 1207.200 2714.830 1207.480 ;
        RECT 2715.010 869.240 2715.290 869.520 ;
        RECT 2715.010 820.960 2715.290 821.240 ;
        RECT 2715.930 531.280 2716.210 531.560 ;
        RECT 2716.850 531.280 2717.130 531.560 ;
        RECT 2714.550 385.760 2714.830 386.040 ;
        RECT 2715.930 385.760 2716.210 386.040 ;
        RECT 2900.850 146.400 2901.130 146.680 ;
      LAYER met3 ;
        RECT 2714.525 1225.850 2714.855 1225.865 ;
        RECT 2699.740 1225.800 2714.855 1225.850 ;
        RECT 2696.000 1225.550 2714.855 1225.800 ;
        RECT 2696.000 1225.200 2700.000 1225.550 ;
        RECT 2714.525 1225.535 2714.855 1225.550 ;
        RECT 2710.845 1207.490 2711.175 1207.505 ;
        RECT 2714.525 1207.490 2714.855 1207.505 ;
        RECT 2710.845 1207.190 2714.855 1207.490 ;
        RECT 2710.845 1207.175 2711.175 1207.190 ;
        RECT 2714.525 1207.175 2714.855 1207.190 ;
        RECT 2714.985 869.540 2715.315 869.545 ;
        RECT 2714.985 869.530 2715.570 869.540 ;
        RECT 2714.985 869.230 2715.770 869.530 ;
        RECT 2714.985 869.220 2715.570 869.230 ;
        RECT 2714.985 869.215 2715.315 869.220 ;
        RECT 2714.985 821.260 2715.315 821.265 ;
        RECT 2714.985 821.250 2715.570 821.260 ;
        RECT 2714.985 820.950 2715.770 821.250 ;
        RECT 2714.985 820.940 2715.570 820.950 ;
        RECT 2714.985 820.935 2715.315 820.940 ;
        RECT 2715.905 531.570 2716.235 531.585 ;
        RECT 2716.825 531.570 2717.155 531.585 ;
        RECT 2715.905 531.270 2717.155 531.570 ;
        RECT 2715.905 531.255 2716.235 531.270 ;
        RECT 2716.825 531.255 2717.155 531.270 ;
        RECT 2714.525 386.050 2714.855 386.065 ;
        RECT 2715.905 386.050 2716.235 386.065 ;
        RECT 2714.525 385.750 2716.235 386.050 ;
        RECT 2714.525 385.735 2714.855 385.750 ;
        RECT 2715.905 385.735 2716.235 385.750 ;
        RECT 2900.825 146.690 2901.155 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2900.825 146.390 2924.800 146.690 ;
        RECT 2900.825 146.375 2901.155 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
      LAYER via3 ;
        RECT 2715.220 869.220 2715.540 869.540 ;
        RECT 2715.220 820.940 2715.540 821.260 ;
      LAYER met4 ;
        RECT 2715.215 869.215 2715.545 869.545 ;
        RECT 2715.230 821.265 2715.530 869.215 ;
        RECT 2715.215 820.935 2715.545 821.265 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2859.890 2491.080 2860.210 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 2859.890 2490.940 2901.150 2491.080 ;
        RECT 2859.890 2490.880 2860.210 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 2713.150 1545.540 2713.470 1545.600 ;
        RECT 2859.890 1545.540 2860.210 1545.600 ;
        RECT 2713.150 1545.400 2860.210 1545.540 ;
        RECT 2713.150 1545.340 2713.470 1545.400 ;
        RECT 2859.890 1545.340 2860.210 1545.400 ;
      LAYER via ;
        RECT 2859.920 2490.880 2860.180 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 2713.180 1545.340 2713.440 1545.600 ;
        RECT 2859.920 1545.340 2860.180 1545.600 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 2859.920 2490.850 2860.180 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 2859.980 1545.630 2860.120 2490.850 ;
        RECT 2713.180 1545.310 2713.440 1545.630 ;
        RECT 2859.920 1545.310 2860.180 1545.630 ;
        RECT 2713.240 1542.085 2713.380 1545.310 ;
        RECT 2713.170 1541.715 2713.450 1542.085 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
        RECT 2713.170 1541.760 2713.450 1542.040 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
        RECT 2713.145 1542.050 2713.475 1542.065 ;
        RECT 2699.740 1542.000 2713.475 1542.050 ;
        RECT 2696.000 1541.750 2713.475 1542.000 ;
        RECT 2696.000 1541.400 2700.000 1541.750 ;
        RECT 2713.145 1541.735 2713.475 1541.750 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2866.790 2725.680 2867.110 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 2866.790 2725.540 2901.150 2725.680 ;
        RECT 2866.790 2725.480 2867.110 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 2713.150 1573.080 2713.470 1573.140 ;
        RECT 2866.790 1573.080 2867.110 1573.140 ;
        RECT 2713.150 1572.940 2867.110 1573.080 ;
        RECT 2713.150 1572.880 2713.470 1572.940 ;
        RECT 2866.790 1572.880 2867.110 1572.940 ;
      LAYER via ;
        RECT 2866.820 2725.480 2867.080 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 2713.180 1572.880 2713.440 1573.140 ;
        RECT 2866.820 1572.880 2867.080 1573.140 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 2866.820 2725.450 2867.080 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 2713.170 1572.995 2713.450 1573.365 ;
        RECT 2866.880 1573.170 2867.020 2725.450 ;
        RECT 2713.180 1572.850 2713.440 1572.995 ;
        RECT 2866.820 1572.850 2867.080 1573.170 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
        RECT 2713.170 1573.040 2713.450 1573.320 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
        RECT 2713.145 1573.330 2713.475 1573.345 ;
        RECT 2699.740 1573.280 2713.475 1573.330 ;
        RECT 2696.000 1573.030 2713.475 1573.280 ;
        RECT 2696.000 1572.680 2700.000 1573.030 ;
        RECT 2713.145 1573.015 2713.475 1573.030 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2873.690 2960.280 2874.010 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 2873.690 2960.140 2901.150 2960.280 ;
        RECT 2873.690 2960.080 2874.010 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
        RECT 2713.150 1607.760 2713.470 1607.820 ;
        RECT 2873.690 1607.760 2874.010 1607.820 ;
        RECT 2713.150 1607.620 2874.010 1607.760 ;
        RECT 2713.150 1607.560 2713.470 1607.620 ;
        RECT 2873.690 1607.560 2874.010 1607.620 ;
      LAYER via ;
        RECT 2873.720 2960.080 2873.980 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
        RECT 2713.180 1607.560 2713.440 1607.820 ;
        RECT 2873.720 1607.560 2873.980 1607.820 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 2873.720 2960.050 2873.980 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 2873.780 1607.850 2873.920 2960.050 ;
        RECT 2713.180 1607.530 2713.440 1607.850 ;
        RECT 2873.720 1607.530 2873.980 1607.850 ;
        RECT 2713.240 1605.325 2713.380 1607.530 ;
        RECT 2713.170 1604.955 2713.450 1605.325 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
        RECT 2713.170 1605.000 2713.450 1605.280 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
        RECT 2713.145 1605.290 2713.475 1605.305 ;
        RECT 2699.740 1605.240 2713.475 1605.290 ;
        RECT 2696.000 1604.990 2713.475 1605.240 ;
        RECT 2696.000 1604.640 2700.000 1604.990 ;
        RECT 2713.145 1604.975 2713.475 1604.990 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2825.390 3194.880 2825.710 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 2825.390 3194.740 2901.150 3194.880 ;
        RECT 2825.390 3194.680 2825.710 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
        RECT 2713.150 1642.100 2713.470 1642.160 ;
        RECT 2825.390 1642.100 2825.710 1642.160 ;
        RECT 2713.150 1641.960 2825.710 1642.100 ;
        RECT 2713.150 1641.900 2713.470 1641.960 ;
        RECT 2825.390 1641.900 2825.710 1641.960 ;
      LAYER via ;
        RECT 2825.420 3194.680 2825.680 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
        RECT 2713.180 1641.900 2713.440 1642.160 ;
        RECT 2825.420 1641.900 2825.680 1642.160 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 2825.420 3194.650 2825.680 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 2825.480 1642.190 2825.620 3194.650 ;
        RECT 2713.180 1641.870 2713.440 1642.190 ;
        RECT 2825.420 1641.870 2825.680 1642.190 ;
        RECT 2713.240 1636.605 2713.380 1641.870 ;
        RECT 2713.170 1636.235 2713.450 1636.605 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
        RECT 2713.170 1636.280 2713.450 1636.560 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
        RECT 2713.145 1636.570 2713.475 1636.585 ;
        RECT 2699.740 1636.520 2713.475 1636.570 ;
        RECT 2696.000 1636.270 2713.475 1636.520 ;
        RECT 2696.000 1635.920 2700.000 1636.270 ;
        RECT 2713.145 1636.255 2713.475 1636.270 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2770.190 3429.480 2770.510 3429.540 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2770.190 3429.340 2901.150 3429.480 ;
        RECT 2770.190 3429.280 2770.510 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
        RECT 2713.150 1669.640 2713.470 1669.700 ;
        RECT 2770.190 1669.640 2770.510 1669.700 ;
        RECT 2713.150 1669.500 2770.510 1669.640 ;
        RECT 2713.150 1669.440 2713.470 1669.500 ;
        RECT 2770.190 1669.440 2770.510 1669.500 ;
      LAYER via ;
        RECT 2770.220 3429.280 2770.480 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
        RECT 2713.180 1669.440 2713.440 1669.700 ;
        RECT 2770.220 1669.440 2770.480 1669.700 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 2770.220 3429.250 2770.480 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 2770.280 1669.730 2770.420 3429.250 ;
        RECT 2713.180 1669.410 2713.440 1669.730 ;
        RECT 2770.220 1669.410 2770.480 1669.730 ;
        RECT 2713.240 1668.565 2713.380 1669.410 ;
        RECT 2713.170 1668.195 2713.450 1668.565 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
        RECT 2713.170 1668.240 2713.450 1668.520 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
        RECT 2713.145 1668.530 2713.475 1668.545 ;
        RECT 2699.740 1668.480 2713.475 1668.530 ;
        RECT 2696.000 1668.230 2713.475 1668.480 ;
        RECT 2696.000 1667.880 2700.000 1668.230 ;
        RECT 2713.145 1668.215 2713.475 1668.230 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2716.370 3380.860 2716.690 3380.920 ;
        RECT 2717.750 3380.860 2718.070 3380.920 ;
        RECT 2716.370 3380.720 2718.070 3380.860 ;
        RECT 2716.370 3380.660 2716.690 3380.720 ;
        RECT 2717.750 3380.660 2718.070 3380.720 ;
        RECT 2717.290 3236.360 2717.610 3236.420 ;
        RECT 2717.750 3236.360 2718.070 3236.420 ;
        RECT 2717.290 3236.220 2718.070 3236.360 ;
        RECT 2717.290 3236.160 2717.610 3236.220 ;
        RECT 2717.750 3236.160 2718.070 3236.220 ;
        RECT 2717.290 3202.020 2717.610 3202.080 ;
        RECT 2717.750 3202.020 2718.070 3202.080 ;
        RECT 2717.290 3201.880 2718.070 3202.020 ;
        RECT 2717.290 3201.820 2717.610 3201.880 ;
        RECT 2717.750 3201.820 2718.070 3201.880 ;
        RECT 2716.830 3153.400 2717.150 3153.460 ;
        RECT 2717.750 3153.400 2718.070 3153.460 ;
        RECT 2716.830 3153.260 2718.070 3153.400 ;
        RECT 2716.830 3153.200 2717.150 3153.260 ;
        RECT 2717.750 3153.200 2718.070 3153.260 ;
        RECT 2716.830 3056.840 2717.150 3056.900 ;
        RECT 2717.750 3056.840 2718.070 3056.900 ;
        RECT 2716.830 3056.700 2718.070 3056.840 ;
        RECT 2716.830 3056.640 2717.150 3056.700 ;
        RECT 2717.750 3056.640 2718.070 3056.700 ;
        RECT 2716.830 2960.280 2717.150 2960.340 ;
        RECT 2717.750 2960.280 2718.070 2960.340 ;
        RECT 2716.830 2960.140 2718.070 2960.280 ;
        RECT 2716.830 2960.080 2717.150 2960.140 ;
        RECT 2717.750 2960.080 2718.070 2960.140 ;
        RECT 2716.830 2863.720 2717.150 2863.780 ;
        RECT 2717.750 2863.720 2718.070 2863.780 ;
        RECT 2716.830 2863.580 2718.070 2863.720 ;
        RECT 2716.830 2863.520 2717.150 2863.580 ;
        RECT 2717.750 2863.520 2718.070 2863.580 ;
        RECT 2716.830 2767.160 2717.150 2767.220 ;
        RECT 2717.750 2767.160 2718.070 2767.220 ;
        RECT 2716.830 2767.020 2718.070 2767.160 ;
        RECT 2716.830 2766.960 2717.150 2767.020 ;
        RECT 2717.750 2766.960 2718.070 2767.020 ;
        RECT 2716.830 2670.600 2717.150 2670.660 ;
        RECT 2717.750 2670.600 2718.070 2670.660 ;
        RECT 2716.830 2670.460 2718.070 2670.600 ;
        RECT 2716.830 2670.400 2717.150 2670.460 ;
        RECT 2717.750 2670.400 2718.070 2670.460 ;
        RECT 2716.830 2574.040 2717.150 2574.100 ;
        RECT 2717.750 2574.040 2718.070 2574.100 ;
        RECT 2716.830 2573.900 2718.070 2574.040 ;
        RECT 2716.830 2573.840 2717.150 2573.900 ;
        RECT 2717.750 2573.840 2718.070 2573.900 ;
        RECT 2716.370 2511.820 2716.690 2511.880 ;
        RECT 2717.750 2511.820 2718.070 2511.880 ;
        RECT 2716.370 2511.680 2718.070 2511.820 ;
        RECT 2716.370 2511.620 2716.690 2511.680 ;
        RECT 2717.750 2511.620 2718.070 2511.680 ;
        RECT 2716.370 2463.200 2716.690 2463.260 ;
        RECT 2717.750 2463.200 2718.070 2463.260 ;
        RECT 2716.370 2463.060 2718.070 2463.200 ;
        RECT 2716.370 2463.000 2716.690 2463.060 ;
        RECT 2717.750 2463.000 2718.070 2463.060 ;
        RECT 2716.830 2380.580 2717.150 2380.640 ;
        RECT 2718.210 2380.580 2718.530 2380.640 ;
        RECT 2716.830 2380.440 2718.530 2380.580 ;
        RECT 2716.830 2380.380 2717.150 2380.440 ;
        RECT 2718.210 2380.380 2718.530 2380.440 ;
        RECT 2716.830 2304.760 2717.150 2304.820 ;
        RECT 2718.210 2304.760 2718.530 2304.820 ;
        RECT 2716.830 2304.620 2718.530 2304.760 ;
        RECT 2716.830 2304.560 2717.150 2304.620 ;
        RECT 2718.210 2304.560 2718.530 2304.620 ;
        RECT 2711.770 2259.880 2712.090 2259.940 ;
        RECT 2716.830 2259.880 2717.150 2259.940 ;
        RECT 2711.770 2259.740 2717.150 2259.880 ;
        RECT 2711.770 2259.680 2712.090 2259.740 ;
        RECT 2716.830 2259.680 2717.150 2259.740 ;
        RECT 2711.770 2226.560 2712.090 2226.620 ;
        RECT 2718.670 2226.560 2718.990 2226.620 ;
        RECT 2711.770 2226.420 2718.990 2226.560 ;
        RECT 2711.770 2226.360 2712.090 2226.420 ;
        RECT 2718.670 2226.360 2718.990 2226.420 ;
        RECT 2716.830 2208.200 2717.150 2208.260 ;
        RECT 2718.670 2208.200 2718.990 2208.260 ;
        RECT 2716.830 2208.060 2718.990 2208.200 ;
        RECT 2716.830 2208.000 2717.150 2208.060 ;
        RECT 2718.670 2208.000 2718.990 2208.060 ;
        RECT 2716.830 2186.920 2717.150 2187.180 ;
        RECT 2716.370 2183.380 2716.690 2183.440 ;
        RECT 2716.920 2183.380 2717.060 2186.920 ;
        RECT 2716.370 2183.240 2717.060 2183.380 ;
        RECT 2716.370 2183.180 2716.690 2183.240 ;
        RECT 2716.370 2138.980 2716.690 2139.240 ;
        RECT 2716.460 2138.840 2716.600 2138.980 ;
        RECT 2716.830 2138.840 2717.150 2138.900 ;
        RECT 2716.460 2138.700 2717.150 2138.840 ;
        RECT 2716.830 2138.640 2717.150 2138.700 ;
        RECT 2716.830 2090.700 2717.150 2090.960 ;
        RECT 2716.920 2090.220 2717.060 2090.700 ;
        RECT 2717.290 2090.220 2717.610 2090.280 ;
        RECT 2716.920 2090.080 2717.610 2090.220 ;
        RECT 2717.290 2090.020 2717.610 2090.080 ;
        RECT 2717.290 2022.360 2717.610 2022.620 ;
        RECT 2717.380 2021.940 2717.520 2022.360 ;
        RECT 2717.290 2021.680 2717.610 2021.940 ;
        RECT 2715.910 1931.780 2716.230 1931.840 ;
        RECT 2717.290 1931.780 2717.610 1931.840 ;
        RECT 2715.910 1931.640 2717.610 1931.780 ;
        RECT 2715.910 1931.580 2716.230 1931.640 ;
        RECT 2717.290 1931.580 2717.610 1931.640 ;
        RECT 2715.910 1883.840 2716.230 1883.900 ;
        RECT 2716.830 1883.840 2717.150 1883.900 ;
        RECT 2715.910 1883.700 2717.150 1883.840 ;
        RECT 2715.910 1883.640 2716.230 1883.700 ;
        RECT 2716.830 1883.640 2717.150 1883.700 ;
        RECT 2715.910 1835.220 2716.230 1835.280 ;
        RECT 2717.290 1835.220 2717.610 1835.280 ;
        RECT 2715.910 1835.080 2717.610 1835.220 ;
        RECT 2715.910 1835.020 2716.230 1835.080 ;
        RECT 2717.290 1835.020 2717.610 1835.080 ;
        RECT 2715.910 1787.280 2716.230 1787.340 ;
        RECT 2716.830 1787.280 2717.150 1787.340 ;
        RECT 2715.910 1787.140 2717.150 1787.280 ;
        RECT 2715.910 1787.080 2716.230 1787.140 ;
        RECT 2716.830 1787.080 2717.150 1787.140 ;
      LAYER via ;
        RECT 2716.400 3380.660 2716.660 3380.920 ;
        RECT 2717.780 3380.660 2718.040 3380.920 ;
        RECT 2717.320 3236.160 2717.580 3236.420 ;
        RECT 2717.780 3236.160 2718.040 3236.420 ;
        RECT 2717.320 3201.820 2717.580 3202.080 ;
        RECT 2717.780 3201.820 2718.040 3202.080 ;
        RECT 2716.860 3153.200 2717.120 3153.460 ;
        RECT 2717.780 3153.200 2718.040 3153.460 ;
        RECT 2716.860 3056.640 2717.120 3056.900 ;
        RECT 2717.780 3056.640 2718.040 3056.900 ;
        RECT 2716.860 2960.080 2717.120 2960.340 ;
        RECT 2717.780 2960.080 2718.040 2960.340 ;
        RECT 2716.860 2863.520 2717.120 2863.780 ;
        RECT 2717.780 2863.520 2718.040 2863.780 ;
        RECT 2716.860 2766.960 2717.120 2767.220 ;
        RECT 2717.780 2766.960 2718.040 2767.220 ;
        RECT 2716.860 2670.400 2717.120 2670.660 ;
        RECT 2717.780 2670.400 2718.040 2670.660 ;
        RECT 2716.860 2573.840 2717.120 2574.100 ;
        RECT 2717.780 2573.840 2718.040 2574.100 ;
        RECT 2716.400 2511.620 2716.660 2511.880 ;
        RECT 2717.780 2511.620 2718.040 2511.880 ;
        RECT 2716.400 2463.000 2716.660 2463.260 ;
        RECT 2717.780 2463.000 2718.040 2463.260 ;
        RECT 2716.860 2380.380 2717.120 2380.640 ;
        RECT 2718.240 2380.380 2718.500 2380.640 ;
        RECT 2716.860 2304.560 2717.120 2304.820 ;
        RECT 2718.240 2304.560 2718.500 2304.820 ;
        RECT 2711.800 2259.680 2712.060 2259.940 ;
        RECT 2716.860 2259.680 2717.120 2259.940 ;
        RECT 2711.800 2226.360 2712.060 2226.620 ;
        RECT 2718.700 2226.360 2718.960 2226.620 ;
        RECT 2716.860 2208.000 2717.120 2208.260 ;
        RECT 2718.700 2208.000 2718.960 2208.260 ;
        RECT 2716.860 2186.920 2717.120 2187.180 ;
        RECT 2716.400 2183.180 2716.660 2183.440 ;
        RECT 2716.400 2138.980 2716.660 2139.240 ;
        RECT 2716.860 2138.640 2717.120 2138.900 ;
        RECT 2716.860 2090.700 2717.120 2090.960 ;
        RECT 2717.320 2090.020 2717.580 2090.280 ;
        RECT 2717.320 2022.360 2717.580 2022.620 ;
        RECT 2717.320 2021.680 2717.580 2021.940 ;
        RECT 2715.940 1931.580 2716.200 1931.840 ;
        RECT 2717.320 1931.580 2717.580 1931.840 ;
        RECT 2715.940 1883.640 2716.200 1883.900 ;
        RECT 2716.860 1883.640 2717.120 1883.900 ;
        RECT 2715.940 1835.020 2716.200 1835.280 ;
        RECT 2717.320 1835.020 2717.580 1835.280 ;
        RECT 2715.940 1787.080 2716.200 1787.340 ;
        RECT 2716.860 1787.080 2717.120 1787.340 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3443.250 2717.520 3517.600 ;
        RECT 2717.380 3443.110 2717.980 3443.250 ;
        RECT 2717.840 3380.950 2717.980 3443.110 ;
        RECT 2716.400 3380.630 2716.660 3380.950 ;
        RECT 2717.780 3380.630 2718.040 3380.950 ;
        RECT 2716.460 3346.010 2716.600 3380.630 ;
        RECT 2716.460 3345.870 2717.520 3346.010 ;
        RECT 2717.380 3298.410 2717.520 3345.870 ;
        RECT 2717.380 3298.270 2717.980 3298.410 ;
        RECT 2717.840 3236.450 2717.980 3298.270 ;
        RECT 2717.320 3236.130 2717.580 3236.450 ;
        RECT 2717.780 3236.130 2718.040 3236.450 ;
        RECT 2717.380 3202.110 2717.520 3236.130 ;
        RECT 2717.320 3201.790 2717.580 3202.110 ;
        RECT 2717.780 3201.790 2718.040 3202.110 ;
        RECT 2717.840 3153.490 2717.980 3201.790 ;
        RECT 2716.860 3153.170 2717.120 3153.490 ;
        RECT 2717.780 3153.170 2718.040 3153.490 ;
        RECT 2716.920 3152.890 2717.060 3153.170 ;
        RECT 2716.920 3152.750 2717.520 3152.890 ;
        RECT 2717.380 3105.290 2717.520 3152.750 ;
        RECT 2717.380 3105.150 2717.980 3105.290 ;
        RECT 2717.840 3056.930 2717.980 3105.150 ;
        RECT 2716.860 3056.610 2717.120 3056.930 ;
        RECT 2717.780 3056.610 2718.040 3056.930 ;
        RECT 2716.920 3056.330 2717.060 3056.610 ;
        RECT 2716.920 3056.190 2717.520 3056.330 ;
        RECT 2717.380 3008.730 2717.520 3056.190 ;
        RECT 2717.380 3008.590 2717.980 3008.730 ;
        RECT 2717.840 2960.370 2717.980 3008.590 ;
        RECT 2716.860 2960.050 2717.120 2960.370 ;
        RECT 2717.780 2960.050 2718.040 2960.370 ;
        RECT 2716.920 2959.770 2717.060 2960.050 ;
        RECT 2716.920 2959.630 2717.520 2959.770 ;
        RECT 2717.380 2912.170 2717.520 2959.630 ;
        RECT 2717.380 2912.030 2717.980 2912.170 ;
        RECT 2717.840 2863.810 2717.980 2912.030 ;
        RECT 2716.860 2863.490 2717.120 2863.810 ;
        RECT 2717.780 2863.490 2718.040 2863.810 ;
        RECT 2716.920 2863.210 2717.060 2863.490 ;
        RECT 2716.920 2863.070 2717.520 2863.210 ;
        RECT 2717.380 2815.610 2717.520 2863.070 ;
        RECT 2717.380 2815.470 2717.980 2815.610 ;
        RECT 2717.840 2767.250 2717.980 2815.470 ;
        RECT 2716.860 2766.930 2717.120 2767.250 ;
        RECT 2717.780 2766.930 2718.040 2767.250 ;
        RECT 2716.920 2766.650 2717.060 2766.930 ;
        RECT 2716.920 2766.510 2717.520 2766.650 ;
        RECT 2717.380 2719.050 2717.520 2766.510 ;
        RECT 2717.380 2718.910 2717.980 2719.050 ;
        RECT 2717.840 2670.690 2717.980 2718.910 ;
        RECT 2716.860 2670.370 2717.120 2670.690 ;
        RECT 2717.780 2670.370 2718.040 2670.690 ;
        RECT 2716.920 2670.090 2717.060 2670.370 ;
        RECT 2716.920 2669.950 2717.520 2670.090 ;
        RECT 2717.380 2622.490 2717.520 2669.950 ;
        RECT 2717.380 2622.350 2717.980 2622.490 ;
        RECT 2717.840 2574.130 2717.980 2622.350 ;
        RECT 2716.860 2573.810 2717.120 2574.130 ;
        RECT 2717.780 2573.810 2718.040 2574.130 ;
        RECT 2716.920 2573.530 2717.060 2573.810 ;
        RECT 2716.920 2573.390 2717.520 2573.530 ;
        RECT 2717.380 2560.045 2717.520 2573.390 ;
        RECT 2716.390 2559.675 2716.670 2560.045 ;
        RECT 2717.310 2559.675 2717.590 2560.045 ;
        RECT 2716.460 2511.910 2716.600 2559.675 ;
        RECT 2716.400 2511.590 2716.660 2511.910 ;
        RECT 2717.780 2511.590 2718.040 2511.910 ;
        RECT 2717.840 2463.290 2717.980 2511.590 ;
        RECT 2716.400 2462.970 2716.660 2463.290 ;
        RECT 2717.780 2462.970 2718.040 2463.290 ;
        RECT 2716.460 2415.205 2716.600 2462.970 ;
        RECT 2716.390 2414.835 2716.670 2415.205 ;
        RECT 2717.310 2414.835 2717.590 2415.205 ;
        RECT 2717.380 2404.890 2717.520 2414.835 ;
        RECT 2716.920 2404.750 2717.520 2404.890 ;
        RECT 2716.920 2380.670 2717.060 2404.750 ;
        RECT 2716.860 2380.350 2717.120 2380.670 ;
        RECT 2718.240 2380.350 2718.500 2380.670 ;
        RECT 2718.300 2304.850 2718.440 2380.350 ;
        RECT 2716.860 2304.530 2717.120 2304.850 ;
        RECT 2718.240 2304.530 2718.500 2304.850 ;
        RECT 2716.920 2259.970 2717.060 2304.530 ;
        RECT 2711.800 2259.650 2712.060 2259.970 ;
        RECT 2716.860 2259.650 2717.120 2259.970 ;
        RECT 2711.860 2226.650 2712.000 2259.650 ;
        RECT 2711.800 2226.330 2712.060 2226.650 ;
        RECT 2718.700 2226.330 2718.960 2226.650 ;
        RECT 2718.760 2208.290 2718.900 2226.330 ;
        RECT 2716.860 2207.970 2717.120 2208.290 ;
        RECT 2718.700 2207.970 2718.960 2208.290 ;
        RECT 2716.920 2187.210 2717.060 2207.970 ;
        RECT 2716.860 2186.890 2717.120 2187.210 ;
        RECT 2716.400 2183.150 2716.660 2183.470 ;
        RECT 2716.460 2139.270 2716.600 2183.150 ;
        RECT 2716.400 2138.950 2716.660 2139.270 ;
        RECT 2716.860 2138.610 2717.120 2138.930 ;
        RECT 2716.920 2090.990 2717.060 2138.610 ;
        RECT 2716.860 2090.670 2717.120 2090.990 ;
        RECT 2717.320 2089.990 2717.580 2090.310 ;
        RECT 2717.380 2022.650 2717.520 2089.990 ;
        RECT 2717.320 2022.330 2717.580 2022.650 ;
        RECT 2717.320 2021.650 2717.580 2021.970 ;
        RECT 2717.380 1997.685 2717.520 2021.650 ;
        RECT 2717.310 1997.315 2717.590 1997.685 ;
        RECT 2717.310 1944.955 2717.590 1945.325 ;
        RECT 2717.380 1931.870 2717.520 1944.955 ;
        RECT 2715.940 1931.550 2716.200 1931.870 ;
        RECT 2717.320 1931.550 2717.580 1931.870 ;
        RECT 2716.000 1883.930 2716.140 1931.550 ;
        RECT 2715.940 1883.610 2716.200 1883.930 ;
        RECT 2716.860 1883.610 2717.120 1883.930 ;
        RECT 2716.920 1883.445 2717.060 1883.610 ;
        RECT 2716.850 1883.075 2717.130 1883.445 ;
        RECT 2717.310 1848.395 2717.590 1848.765 ;
        RECT 2717.380 1835.310 2717.520 1848.395 ;
        RECT 2715.940 1834.990 2716.200 1835.310 ;
        RECT 2717.320 1834.990 2717.580 1835.310 ;
        RECT 2716.000 1787.370 2716.140 1834.990 ;
        RECT 2715.940 1787.050 2716.200 1787.370 ;
        RECT 2716.860 1787.050 2717.120 1787.370 ;
        RECT 2716.920 1786.885 2717.060 1787.050 ;
        RECT 2716.850 1786.515 2717.130 1786.885 ;
        RECT 2717.310 1751.835 2717.590 1752.205 ;
        RECT 2717.380 1699.845 2717.520 1751.835 ;
        RECT 2717.310 1699.475 2717.590 1699.845 ;
      LAYER via2 ;
        RECT 2716.390 2559.720 2716.670 2560.000 ;
        RECT 2717.310 2559.720 2717.590 2560.000 ;
        RECT 2716.390 2414.880 2716.670 2415.160 ;
        RECT 2717.310 2414.880 2717.590 2415.160 ;
        RECT 2717.310 1997.360 2717.590 1997.640 ;
        RECT 2717.310 1945.000 2717.590 1945.280 ;
        RECT 2716.850 1883.120 2717.130 1883.400 ;
        RECT 2717.310 1848.440 2717.590 1848.720 ;
        RECT 2716.850 1786.560 2717.130 1786.840 ;
        RECT 2717.310 1751.880 2717.590 1752.160 ;
        RECT 2717.310 1699.520 2717.590 1699.800 ;
      LAYER met3 ;
        RECT 2716.365 2560.010 2716.695 2560.025 ;
        RECT 2717.285 2560.010 2717.615 2560.025 ;
        RECT 2716.365 2559.710 2717.615 2560.010 ;
        RECT 2716.365 2559.695 2716.695 2559.710 ;
        RECT 2717.285 2559.695 2717.615 2559.710 ;
        RECT 2716.365 2415.170 2716.695 2415.185 ;
        RECT 2717.285 2415.170 2717.615 2415.185 ;
        RECT 2716.365 2414.870 2717.615 2415.170 ;
        RECT 2716.365 2414.855 2716.695 2414.870 ;
        RECT 2717.285 2414.855 2717.615 2414.870 ;
        RECT 2717.285 1997.660 2717.615 1997.665 ;
        RECT 2717.030 1997.650 2717.615 1997.660 ;
        RECT 2716.830 1997.350 2717.615 1997.650 ;
        RECT 2717.030 1997.340 2717.615 1997.350 ;
        RECT 2717.285 1997.335 2717.615 1997.340 ;
        RECT 2717.285 1945.300 2717.615 1945.305 ;
        RECT 2717.030 1945.290 2717.615 1945.300 ;
        RECT 2716.830 1944.990 2717.615 1945.290 ;
        RECT 2717.030 1944.980 2717.615 1944.990 ;
        RECT 2717.285 1944.975 2717.615 1944.980 ;
        RECT 2716.825 1883.420 2717.155 1883.425 ;
        RECT 2716.825 1883.410 2717.410 1883.420 ;
        RECT 2716.825 1883.110 2717.610 1883.410 ;
        RECT 2716.825 1883.100 2717.410 1883.110 ;
        RECT 2716.825 1883.095 2717.155 1883.100 ;
        RECT 2717.285 1848.740 2717.615 1848.745 ;
        RECT 2717.030 1848.730 2717.615 1848.740 ;
        RECT 2716.830 1848.430 2717.615 1848.730 ;
        RECT 2717.030 1848.420 2717.615 1848.430 ;
        RECT 2717.285 1848.415 2717.615 1848.420 ;
        RECT 2716.825 1786.860 2717.155 1786.865 ;
        RECT 2716.825 1786.850 2717.410 1786.860 ;
        RECT 2716.825 1786.550 2717.610 1786.850 ;
        RECT 2716.825 1786.540 2717.410 1786.550 ;
        RECT 2716.825 1786.535 2717.155 1786.540 ;
        RECT 2717.285 1752.180 2717.615 1752.185 ;
        RECT 2717.030 1752.170 2717.615 1752.180 ;
        RECT 2716.830 1751.870 2717.615 1752.170 ;
        RECT 2717.030 1751.860 2717.615 1751.870 ;
        RECT 2717.285 1751.855 2717.615 1751.860 ;
        RECT 2717.285 1699.810 2717.615 1699.825 ;
        RECT 2699.740 1699.760 2717.615 1699.810 ;
        RECT 2696.000 1699.510 2717.615 1699.760 ;
        RECT 2696.000 1699.160 2700.000 1699.510 ;
        RECT 2717.285 1699.495 2717.615 1699.510 ;
      LAYER via3 ;
        RECT 2717.060 1997.340 2717.380 1997.660 ;
        RECT 2717.060 1944.980 2717.380 1945.300 ;
        RECT 2717.060 1883.100 2717.380 1883.420 ;
        RECT 2717.060 1848.420 2717.380 1848.740 ;
        RECT 2717.060 1786.540 2717.380 1786.860 ;
        RECT 2717.060 1751.860 2717.380 1752.180 ;
      LAYER met4 ;
        RECT 2717.055 1997.335 2717.385 1997.665 ;
        RECT 2717.070 1945.305 2717.370 1997.335 ;
        RECT 2717.055 1944.975 2717.385 1945.305 ;
        RECT 2717.055 1883.095 2717.385 1883.425 ;
        RECT 2717.070 1848.745 2717.370 1883.095 ;
        RECT 2717.055 1848.415 2717.385 1848.745 ;
        RECT 2717.055 1786.535 2717.385 1786.865 ;
        RECT 2717.070 1752.185 2717.370 1786.535 ;
        RECT 2717.055 1751.855 2717.385 1752.185 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2392.530 3504.620 2392.850 3504.680 ;
        RECT 2697.970 3504.620 2698.290 3504.680 ;
        RECT 2392.530 3504.480 2698.290 3504.620 ;
        RECT 2392.530 3504.420 2392.850 3504.480 ;
        RECT 2697.970 3504.420 2698.290 3504.480 ;
      LAYER via ;
        RECT 2392.560 3504.420 2392.820 3504.680 ;
        RECT 2698.000 3504.420 2698.260 3504.680 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3504.710 2392.760 3517.600 ;
        RECT 2392.560 3504.390 2392.820 3504.710 ;
        RECT 2698.000 3504.390 2698.260 3504.710 ;
        RECT 2698.060 1732.485 2698.200 3504.390 ;
        RECT 2697.990 1732.115 2698.270 1732.485 ;
      LAYER via2 ;
        RECT 2697.990 1732.160 2698.270 1732.440 ;
      LAYER met3 ;
        RECT 2697.965 1732.450 2698.295 1732.465 ;
        RECT 2697.750 1732.135 2698.295 1732.450 ;
        RECT 2697.750 1731.720 2698.050 1732.135 ;
        RECT 2696.000 1731.120 2700.000 1731.720 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2068.230 3504.280 2068.550 3504.340 ;
        RECT 2698.430 3504.280 2698.750 3504.340 ;
        RECT 2068.230 3504.140 2698.750 3504.280 ;
        RECT 2068.230 3504.080 2068.550 3504.140 ;
        RECT 2698.430 3504.080 2698.750 3504.140 ;
      LAYER via ;
        RECT 2068.260 3504.080 2068.520 3504.340 ;
        RECT 2698.460 3504.080 2698.720 3504.340 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3504.370 2068.460 3517.600 ;
        RECT 2068.260 3504.050 2068.520 3504.370 ;
        RECT 2698.460 3504.050 2698.720 3504.370 ;
        RECT 2698.520 1765.805 2698.660 3504.050 ;
        RECT 2698.450 1765.435 2698.730 1765.805 ;
      LAYER via2 ;
        RECT 2698.450 1765.480 2698.730 1765.760 ;
      LAYER met3 ;
        RECT 2698.425 1765.770 2698.755 1765.785 ;
        RECT 2698.425 1765.455 2698.970 1765.770 ;
        RECT 2698.670 1763.000 2698.970 1765.455 ;
        RECT 2696.000 1762.400 2700.000 1763.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1743.930 3503.940 1744.250 3504.000 ;
        RECT 2698.890 3503.940 2699.210 3504.000 ;
        RECT 1743.930 3503.800 2699.210 3503.940 ;
        RECT 1743.930 3503.740 1744.250 3503.800 ;
        RECT 2698.890 3503.740 2699.210 3503.800 ;
      LAYER via ;
        RECT 1743.960 3503.740 1744.220 3504.000 ;
        RECT 2698.920 3503.740 2699.180 3504.000 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3504.030 1744.160 3517.600 ;
        RECT 1743.960 3503.710 1744.220 3504.030 ;
        RECT 2698.920 3503.710 2699.180 3504.030 ;
        RECT 2698.980 1797.765 2699.120 3503.710 ;
        RECT 2698.910 1797.395 2699.190 1797.765 ;
      LAYER via2 ;
        RECT 2698.910 1797.440 2699.190 1797.720 ;
      LAYER met3 ;
        RECT 2698.885 1797.730 2699.215 1797.745 ;
        RECT 2698.670 1797.415 2699.215 1797.730 ;
        RECT 2698.670 1794.960 2698.970 1797.415 ;
        RECT 2696.000 1794.360 2700.000 1794.960 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3503.260 1419.490 3503.320 ;
        RECT 2696.130 3503.260 2696.450 3503.320 ;
        RECT 1419.170 3503.120 2696.450 3503.260 ;
        RECT 1419.170 3503.060 1419.490 3503.120 ;
        RECT 2696.130 3503.060 2696.450 3503.120 ;
        RECT 2696.130 1828.420 2696.450 1828.480 ;
        RECT 2697.510 1828.420 2697.830 1828.480 ;
        RECT 2696.130 1828.280 2697.830 1828.420 ;
        RECT 2696.130 1828.220 2696.450 1828.280 ;
        RECT 2697.510 1828.220 2697.830 1828.280 ;
      LAYER via ;
        RECT 1419.200 3503.060 1419.460 3503.320 ;
        RECT 2696.160 3503.060 2696.420 3503.320 ;
        RECT 2696.160 1828.220 2696.420 1828.480 ;
        RECT 2697.540 1828.220 2697.800 1828.480 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3503.350 1419.400 3517.600 ;
        RECT 1419.200 3503.030 1419.460 3503.350 ;
        RECT 2696.160 3503.030 2696.420 3503.350 ;
        RECT 2696.220 1828.510 2696.360 3503.030 ;
        RECT 2696.160 1828.190 2696.420 1828.510 ;
        RECT 2697.540 1828.365 2697.800 1828.510 ;
        RECT 2697.530 1827.995 2697.810 1828.365 ;
      LAYER via2 ;
        RECT 2697.530 1828.040 2697.810 1828.320 ;
      LAYER met3 ;
        RECT 2697.505 1828.330 2697.835 1828.345 ;
        RECT 2697.100 1828.030 2698.050 1828.330 ;
        RECT 2697.505 1828.015 2698.050 1828.030 ;
        RECT 2697.750 1826.240 2698.050 1828.015 ;
        RECT 2696.000 1825.640 2700.000 1826.240 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2715.450 545.400 2715.770 545.660 ;
        RECT 2715.540 544.980 2715.680 545.400 ;
        RECT 2715.450 544.720 2715.770 544.980 ;
        RECT 2900.830 386.140 2901.150 386.200 ;
        RECT 2715.540 386.000 2901.150 386.140 ;
        RECT 2715.540 385.860 2715.680 386.000 ;
        RECT 2900.830 385.940 2901.150 386.000 ;
        RECT 2715.450 385.600 2715.770 385.860 ;
      LAYER via ;
        RECT 2715.480 545.400 2715.740 545.660 ;
        RECT 2715.480 544.720 2715.740 544.980 ;
        RECT 2900.860 385.940 2901.120 386.200 ;
        RECT 2715.480 385.600 2715.740 385.860 ;
      LAYER met2 ;
        RECT 2715.470 1257.475 2715.750 1257.845 ;
        RECT 2715.540 545.690 2715.680 1257.475 ;
        RECT 2715.480 545.370 2715.740 545.690 ;
        RECT 2715.480 544.690 2715.740 545.010 ;
        RECT 2715.540 385.890 2715.680 544.690 ;
        RECT 2900.860 385.910 2901.120 386.230 ;
        RECT 2715.480 385.570 2715.740 385.890 ;
        RECT 2900.920 381.325 2901.060 385.910 ;
        RECT 2900.850 380.955 2901.130 381.325 ;
      LAYER via2 ;
        RECT 2715.470 1257.520 2715.750 1257.800 ;
        RECT 2900.850 381.000 2901.130 381.280 ;
      LAYER met3 ;
        RECT 2715.445 1257.810 2715.775 1257.825 ;
        RECT 2699.740 1257.760 2715.775 1257.810 ;
        RECT 2696.000 1257.510 2715.775 1257.760 ;
        RECT 2696.000 1257.160 2700.000 1257.510 ;
        RECT 2715.445 1257.495 2715.775 1257.510 ;
        RECT 2900.825 381.290 2901.155 381.305 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2900.825 380.990 2924.800 381.290 ;
        RECT 2900.825 380.975 2901.155 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3502.920 1095.190 3502.980 ;
        RECT 2699.810 3502.920 2700.130 3502.980 ;
        RECT 1094.870 3502.780 2700.130 3502.920 ;
        RECT 1094.870 3502.720 1095.190 3502.780 ;
        RECT 2699.810 3502.720 2700.130 3502.780 ;
      LAYER via ;
        RECT 1094.900 3502.720 1095.160 3502.980 ;
        RECT 2699.840 3502.720 2700.100 3502.980 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3503.010 1095.100 3517.600 ;
        RECT 1094.900 3502.690 1095.160 3503.010 ;
        RECT 2699.840 3502.690 2700.100 3503.010 ;
        RECT 2699.900 1860.325 2700.040 3502.690 ;
        RECT 2699.830 1859.955 2700.110 1860.325 ;
      LAYER via2 ;
        RECT 2699.830 1860.000 2700.110 1860.280 ;
      LAYER met3 ;
        RECT 2699.805 1860.290 2700.135 1860.305 ;
        RECT 2699.590 1859.975 2700.135 1860.290 ;
        RECT 2699.590 1857.520 2699.890 1859.975 ;
        RECT 2696.000 1856.920 2700.000 1857.520 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3502.240 770.890 3502.300 ;
        RECT 2700.270 3502.240 2700.590 3502.300 ;
        RECT 770.570 3502.100 2700.590 3502.240 ;
        RECT 770.570 3502.040 770.890 3502.100 ;
        RECT 2700.270 3502.040 2700.590 3502.100 ;
      LAYER via ;
        RECT 770.600 3502.040 770.860 3502.300 ;
        RECT 2700.300 3502.040 2700.560 3502.300 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3502.330 770.800 3517.600 ;
        RECT 770.600 3502.010 770.860 3502.330 ;
        RECT 2700.300 3502.010 2700.560 3502.330 ;
        RECT 2700.360 1890.245 2700.500 3502.010 ;
        RECT 2700.290 1889.875 2700.570 1890.245 ;
      LAYER via2 ;
        RECT 2700.290 1889.920 2700.570 1890.200 ;
      LAYER met3 ;
        RECT 2700.265 1890.210 2700.595 1890.225 ;
        RECT 2699.590 1889.910 2700.595 1890.210 ;
        RECT 2699.590 1889.480 2699.890 1889.910 ;
        RECT 2700.265 1889.895 2700.595 1889.910 ;
        RECT 2696.000 1888.880 2700.000 1889.480 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3503.205 446.040 3517.600 ;
        RECT 445.830 3502.835 446.110 3503.205 ;
      LAYER via2 ;
        RECT 445.830 3502.880 446.110 3503.160 ;
      LAYER met3 ;
        RECT 445.805 3503.170 446.135 3503.185 ;
        RECT 2692.190 3503.170 2692.570 3503.180 ;
        RECT 445.805 3502.870 2692.570 3503.170 ;
        RECT 445.805 3502.855 446.135 3502.870 ;
        RECT 2692.190 3502.860 2692.570 3502.870 ;
        RECT 2696.790 1922.540 2697.170 1922.860 ;
        RECT 2696.830 1920.760 2697.130 1922.540 ;
        RECT 2696.000 1920.160 2700.000 1920.760 ;
      LAYER via3 ;
        RECT 2692.220 3502.860 2692.540 3503.180 ;
        RECT 2696.820 1922.540 2697.140 1922.860 ;
      LAYER met4 ;
        RECT 2692.215 3502.855 2692.545 3503.185 ;
        RECT 2692.230 1997.650 2692.530 3502.855 ;
        RECT 2692.230 1997.350 2693.450 1997.650 ;
        RECT 2693.150 1994.250 2693.450 1997.350 ;
        RECT 2692.230 1993.950 2693.450 1994.250 ;
        RECT 2692.230 1922.850 2692.530 1993.950 ;
        RECT 2696.815 1922.850 2697.145 1922.865 ;
        RECT 2692.230 1922.550 2697.145 1922.850 ;
        RECT 2696.815 1922.535 2697.145 1922.550 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3502.525 121.740 3517.600 ;
        RECT 121.530 3502.155 121.810 3502.525 ;
      LAYER via2 ;
        RECT 121.530 3502.200 121.810 3502.480 ;
      LAYER met3 ;
        RECT 121.505 3502.490 121.835 3502.505 ;
        RECT 2700.470 3502.490 2700.850 3502.500 ;
        RECT 121.505 3502.190 2700.850 3502.490 ;
        RECT 121.505 3502.175 121.835 3502.190 ;
        RECT 2700.470 3502.180 2700.850 3502.190 ;
        RECT 2700.470 1952.770 2700.850 1952.780 ;
        RECT 2699.740 1952.720 2700.850 1952.770 ;
        RECT 2696.000 1952.470 2700.850 1952.720 ;
        RECT 2696.000 1952.120 2700.000 1952.470 ;
        RECT 2700.470 1952.460 2700.850 1952.470 ;
      LAYER via3 ;
        RECT 2700.500 3502.180 2700.820 3502.500 ;
        RECT 2700.500 1952.460 2700.820 1952.780 ;
      LAYER met4 ;
        RECT 2700.495 3502.175 2700.825 3502.505 ;
        RECT 2700.510 1952.785 2700.810 3502.175 ;
        RECT 2700.495 1952.455 2700.825 1952.785 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 2706.250 3339.720 2706.570 3339.780 ;
        RECT 17.090 3339.580 2706.570 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 2706.250 3339.520 2706.570 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 2706.280 3339.520 2706.540 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 2706.280 3339.490 2706.540 3339.810 ;
        RECT 2706.340 1984.085 2706.480 3339.490 ;
        RECT 2706.270 1983.715 2706.550 1984.085 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
        RECT 2706.270 1983.760 2706.550 1984.040 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
        RECT 2706.245 1984.050 2706.575 1984.065 ;
        RECT 2699.740 1984.000 2706.575 1984.050 ;
        RECT 2696.000 1983.750 2706.575 1984.000 ;
        RECT 2696.000 1983.400 2700.000 1983.750 ;
        RECT 2706.245 1983.735 2706.575 1983.750 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3051.740 17.410 3051.800 ;
        RECT 2708.550 3051.740 2708.870 3051.800 ;
        RECT 17.090 3051.600 2708.870 3051.740 ;
        RECT 17.090 3051.540 17.410 3051.600 ;
        RECT 2708.550 3051.540 2708.870 3051.600 ;
      LAYER via ;
        RECT 17.120 3051.540 17.380 3051.800 ;
        RECT 2708.580 3051.540 2708.840 3051.800 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3051.830 17.320 3051.995 ;
        RECT 17.120 3051.510 17.380 3051.830 ;
        RECT 2708.580 3051.510 2708.840 3051.830 ;
        RECT 2708.640 2016.045 2708.780 3051.510 ;
        RECT 2708.570 2015.675 2708.850 2016.045 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
        RECT 2708.570 2015.720 2708.850 2016.000 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
        RECT 2708.545 2016.010 2708.875 2016.025 ;
        RECT 2699.740 2015.960 2708.875 2016.010 ;
        RECT 2696.000 2015.710 2708.875 2015.960 ;
        RECT 2696.000 2015.360 2700.000 2015.710 ;
        RECT 2708.545 2015.695 2708.875 2015.710 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.010 2390.780 18.330 2390.840 ;
        RECT 2714.990 2390.780 2715.310 2390.840 ;
        RECT 18.010 2390.640 2715.310 2390.780 ;
        RECT 18.010 2390.580 18.330 2390.640 ;
        RECT 2714.990 2390.580 2715.310 2390.640 ;
      LAYER via ;
        RECT 18.040 2390.580 18.300 2390.840 ;
        RECT 2715.020 2390.580 2715.280 2390.840 ;
      LAYER met2 ;
        RECT 18.030 2765.035 18.310 2765.405 ;
        RECT 18.100 2390.870 18.240 2765.035 ;
        RECT 18.040 2390.550 18.300 2390.870 ;
        RECT 2715.020 2390.550 2715.280 2390.870 ;
        RECT 2715.080 2047.325 2715.220 2390.550 ;
        RECT 2715.010 2046.955 2715.290 2047.325 ;
      LAYER via2 ;
        RECT 18.030 2765.080 18.310 2765.360 ;
        RECT 2715.010 2047.000 2715.290 2047.280 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 18.005 2765.370 18.335 2765.385 ;
        RECT -4.800 2765.070 18.335 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 18.005 2765.055 18.335 2765.070 ;
        RECT 2714.985 2047.290 2715.315 2047.305 ;
        RECT 2699.740 2047.240 2715.315 2047.290 ;
        RECT 2696.000 2046.990 2715.315 2047.240 ;
        RECT 2696.000 2046.640 2700.000 2046.990 ;
        RECT 2714.985 2046.975 2715.315 2046.990 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2477.480 16.950 2477.540 ;
        RECT 2704.870 2477.480 2705.190 2477.540 ;
        RECT 16.630 2477.340 2705.190 2477.480 ;
        RECT 16.630 2477.280 16.950 2477.340 ;
        RECT 2704.870 2477.280 2705.190 2477.340 ;
      LAYER via ;
        RECT 16.660 2477.280 16.920 2477.540 ;
        RECT 2704.900 2477.280 2705.160 2477.540 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.660 2477.250 16.920 2477.395 ;
        RECT 2704.900 2477.250 2705.160 2477.570 ;
        RECT 2704.960 2079.285 2705.100 2477.250 ;
        RECT 2704.890 2078.915 2705.170 2079.285 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
        RECT 2704.890 2078.960 2705.170 2079.240 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
        RECT 2704.865 2079.250 2705.195 2079.265 ;
        RECT 2699.740 2079.200 2705.195 2079.250 ;
        RECT 2696.000 2078.950 2705.195 2079.200 ;
        RECT 2696.000 2078.600 2700.000 2078.950 ;
        RECT 2704.865 2078.935 2705.195 2078.950 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.570 2394.520 1299.890 2394.580 ;
        RECT 2715.910 2394.520 2716.230 2394.580 ;
        RECT 1299.570 2394.380 2716.230 2394.520 ;
        RECT 1299.570 2394.320 1299.890 2394.380 ;
        RECT 2715.910 2394.320 2716.230 2394.380 ;
        RECT 15.710 2194.260 16.030 2194.320 ;
        RECT 1299.570 2194.260 1299.890 2194.320 ;
        RECT 15.710 2194.120 1299.890 2194.260 ;
        RECT 15.710 2194.060 16.030 2194.120 ;
        RECT 1299.570 2194.060 1299.890 2194.120 ;
      LAYER via ;
        RECT 1299.600 2394.320 1299.860 2394.580 ;
        RECT 2715.940 2394.320 2716.200 2394.580 ;
        RECT 15.740 2194.060 16.000 2194.320 ;
        RECT 1299.600 2194.060 1299.860 2194.320 ;
      LAYER met2 ;
        RECT 1299.600 2394.290 1299.860 2394.610 ;
        RECT 2715.940 2394.290 2716.200 2394.610 ;
        RECT 1299.660 2194.350 1299.800 2394.290 ;
        RECT 15.740 2194.030 16.000 2194.350 ;
        RECT 1299.600 2194.030 1299.860 2194.350 ;
        RECT 15.800 2190.125 15.940 2194.030 ;
        RECT 15.730 2189.755 16.010 2190.125 ;
        RECT 2716.000 2110.565 2716.140 2394.290 ;
        RECT 2715.930 2110.195 2716.210 2110.565 ;
      LAYER via2 ;
        RECT 15.730 2189.800 16.010 2190.080 ;
        RECT 2715.930 2110.240 2716.210 2110.520 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 15.705 2190.090 16.035 2190.105 ;
        RECT -4.800 2189.790 16.035 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 15.705 2189.775 16.035 2189.790 ;
        RECT 2715.905 2110.530 2716.235 2110.545 ;
        RECT 2699.740 2110.480 2716.235 2110.530 ;
        RECT 2696.000 2110.230 2716.235 2110.480 ;
        RECT 2696.000 2109.880 2700.000 2110.230 ;
        RECT 2715.905 2110.215 2716.235 2110.230 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.250 2395.880 1303.570 2395.940 ;
        RECT 2704.410 2395.880 2704.730 2395.940 ;
        RECT 1303.250 2395.740 2704.730 2395.880 ;
        RECT 1303.250 2395.680 1303.570 2395.740 ;
        RECT 2704.410 2395.680 2704.730 2395.740 ;
        RECT 16.170 1904.240 16.490 1904.300 ;
        RECT 1303.250 1904.240 1303.570 1904.300 ;
        RECT 16.170 1904.100 1303.570 1904.240 ;
        RECT 16.170 1904.040 16.490 1904.100 ;
        RECT 1303.250 1904.040 1303.570 1904.100 ;
      LAYER via ;
        RECT 1303.280 2395.680 1303.540 2395.940 ;
        RECT 2704.440 2395.680 2704.700 2395.940 ;
        RECT 16.200 1904.040 16.460 1904.300 ;
        RECT 1303.280 1904.040 1303.540 1904.300 ;
      LAYER met2 ;
        RECT 1303.280 2395.650 1303.540 2395.970 ;
        RECT 2704.440 2395.650 2704.700 2395.970 ;
        RECT 1303.340 1904.330 1303.480 2395.650 ;
        RECT 2704.500 2141.845 2704.640 2395.650 ;
        RECT 2704.430 2141.475 2704.710 2141.845 ;
        RECT 16.200 1904.010 16.460 1904.330 ;
        RECT 1303.280 1904.010 1303.540 1904.330 ;
        RECT 16.260 1903.165 16.400 1904.010 ;
        RECT 16.190 1902.795 16.470 1903.165 ;
      LAYER via2 ;
        RECT 2704.430 2141.520 2704.710 2141.800 ;
        RECT 16.190 1902.840 16.470 1903.120 ;
      LAYER met3 ;
        RECT 2704.405 2141.810 2704.735 2141.825 ;
        RECT 2699.740 2141.760 2704.735 2141.810 ;
        RECT 2696.000 2141.510 2704.735 2141.760 ;
        RECT 2696.000 2141.160 2700.000 2141.510 ;
        RECT 2704.405 2141.495 2704.735 2141.510 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 16.165 1903.130 16.495 1903.145 ;
        RECT -4.800 1902.830 16.495 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 16.165 1902.815 16.495 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1283.740 2713.470 1283.800 ;
        RECT 2790.890 1283.740 2791.210 1283.800 ;
        RECT 2713.150 1283.600 2791.210 1283.740 ;
        RECT 2713.150 1283.540 2713.470 1283.600 ;
        RECT 2790.890 1283.540 2791.210 1283.600 ;
        RECT 2790.890 620.740 2791.210 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 2790.890 620.600 2901.150 620.740 ;
        RECT 2790.890 620.540 2791.210 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 2713.180 1283.540 2713.440 1283.800 ;
        RECT 2790.920 1283.540 2791.180 1283.800 ;
        RECT 2790.920 620.540 2791.180 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 2713.170 1288.755 2713.450 1289.125 ;
        RECT 2713.240 1283.830 2713.380 1288.755 ;
        RECT 2713.180 1283.510 2713.440 1283.830 ;
        RECT 2790.920 1283.510 2791.180 1283.830 ;
        RECT 2790.980 620.830 2791.120 1283.510 ;
        RECT 2790.920 620.510 2791.180 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 2713.170 1288.800 2713.450 1289.080 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 2713.145 1289.090 2713.475 1289.105 ;
        RECT 2699.740 1289.040 2713.475 1289.090 ;
        RECT 2696.000 1288.790 2713.475 1289.040 ;
        RECT 2696.000 1288.440 2700.000 1288.790 ;
        RECT 2713.145 1288.775 2713.475 1288.790 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1301.870 2395.200 1302.190 2395.260 ;
        RECT 2717.290 2395.200 2717.610 2395.260 ;
        RECT 1301.870 2395.060 2717.610 2395.200 ;
        RECT 1301.870 2395.000 1302.190 2395.060 ;
        RECT 2717.290 2395.000 2717.610 2395.060 ;
        RECT 16.170 1621.360 16.490 1621.420 ;
        RECT 1301.870 1621.360 1302.190 1621.420 ;
        RECT 16.170 1621.220 1302.190 1621.360 ;
        RECT 16.170 1621.160 16.490 1621.220 ;
        RECT 1301.870 1621.160 1302.190 1621.220 ;
      LAYER via ;
        RECT 1301.900 2395.000 1302.160 2395.260 ;
        RECT 2717.320 2395.000 2717.580 2395.260 ;
        RECT 16.200 1621.160 16.460 1621.420 ;
        RECT 1301.900 1621.160 1302.160 1621.420 ;
      LAYER met2 ;
        RECT 1301.900 2394.970 1302.160 2395.290 ;
        RECT 2717.320 2394.970 2717.580 2395.290 ;
        RECT 1301.960 1621.450 1302.100 2394.970 ;
        RECT 2717.380 2173.805 2717.520 2394.970 ;
        RECT 2717.310 2173.435 2717.590 2173.805 ;
        RECT 16.200 1621.130 16.460 1621.450 ;
        RECT 1301.900 1621.130 1302.160 1621.450 ;
        RECT 16.260 1615.525 16.400 1621.130 ;
        RECT 16.190 1615.155 16.470 1615.525 ;
      LAYER via2 ;
        RECT 2717.310 2173.480 2717.590 2173.760 ;
        RECT 16.190 1615.200 16.470 1615.480 ;
      LAYER met3 ;
        RECT 2717.285 2173.770 2717.615 2173.785 ;
        RECT 2699.740 2173.720 2717.615 2173.770 ;
        RECT 2696.000 2173.470 2717.615 2173.720 ;
        RECT 2696.000 2173.120 2700.000 2173.470 ;
        RECT 2717.285 2173.455 2717.615 2173.470 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.165 1615.490 16.495 1615.505 ;
        RECT -4.800 1615.190 16.495 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.165 1615.175 16.495 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1300.490 2394.860 1300.810 2394.920 ;
        RECT 2712.230 2394.860 2712.550 2394.920 ;
        RECT 1300.490 2394.720 2712.550 2394.860 ;
        RECT 1300.490 2394.660 1300.810 2394.720 ;
        RECT 2712.230 2394.660 2712.550 2394.720 ;
        RECT 17.090 1400.700 17.410 1400.760 ;
        RECT 1300.490 1400.700 1300.810 1400.760 ;
        RECT 17.090 1400.560 1300.810 1400.700 ;
        RECT 17.090 1400.500 17.410 1400.560 ;
        RECT 1300.490 1400.500 1300.810 1400.560 ;
      LAYER via ;
        RECT 1300.520 2394.660 1300.780 2394.920 ;
        RECT 2712.260 2394.660 2712.520 2394.920 ;
        RECT 17.120 1400.500 17.380 1400.760 ;
        RECT 1300.520 1400.500 1300.780 1400.760 ;
      LAYER met2 ;
        RECT 1300.520 2394.630 1300.780 2394.950 ;
        RECT 2712.260 2394.630 2712.520 2394.950 ;
        RECT 1300.580 1400.790 1300.720 2394.630 ;
        RECT 2712.320 2205.085 2712.460 2394.630 ;
        RECT 2712.250 2204.715 2712.530 2205.085 ;
        RECT 17.120 1400.645 17.380 1400.790 ;
        RECT 17.110 1400.275 17.390 1400.645 ;
        RECT 1300.520 1400.470 1300.780 1400.790 ;
      LAYER via2 ;
        RECT 2712.250 2204.760 2712.530 2205.040 ;
        RECT 17.110 1400.320 17.390 1400.600 ;
      LAYER met3 ;
        RECT 2712.225 2205.050 2712.555 2205.065 ;
        RECT 2699.740 2205.000 2712.555 2205.050 ;
        RECT 2696.000 2204.750 2712.555 2205.000 ;
        RECT 2696.000 2204.400 2700.000 2204.750 ;
        RECT 2712.225 2204.735 2712.555 2204.750 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 17.085 1400.610 17.415 1400.625 ;
        RECT -4.800 1400.310 17.415 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 17.085 1400.295 17.415 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 1186.840 17.410 1186.900 ;
        RECT 2702.110 1186.840 2702.430 1186.900 ;
        RECT 17.090 1186.700 2702.430 1186.840 ;
        RECT 17.090 1186.640 17.410 1186.700 ;
        RECT 2702.110 1186.640 2702.430 1186.700 ;
      LAYER via ;
        RECT 17.120 1186.640 17.380 1186.900 ;
        RECT 2702.140 1186.640 2702.400 1186.900 ;
      LAYER met2 ;
        RECT 2702.130 2236.675 2702.410 2237.045 ;
        RECT 2702.200 1186.930 2702.340 2236.675 ;
        RECT 17.120 1186.610 17.380 1186.930 ;
        RECT 2702.140 1186.610 2702.400 1186.930 ;
        RECT 17.180 1185.085 17.320 1186.610 ;
        RECT 17.110 1184.715 17.390 1185.085 ;
      LAYER via2 ;
        RECT 2702.130 2236.720 2702.410 2237.000 ;
        RECT 17.110 1184.760 17.390 1185.040 ;
      LAYER met3 ;
        RECT 2702.105 2237.010 2702.435 2237.025 ;
        RECT 2699.740 2236.960 2702.435 2237.010 ;
        RECT 2696.000 2236.710 2702.435 2236.960 ;
        RECT 2696.000 2236.360 2700.000 2236.710 ;
        RECT 2702.105 2236.695 2702.435 2236.710 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 17.085 1185.050 17.415 1185.065 ;
        RECT -4.800 1184.750 17.415 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 17.085 1184.735 17.415 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 1004.260 20.630 1004.320 ;
        RECT 2718.210 1004.260 2718.530 1004.320 ;
        RECT 20.310 1004.120 2718.530 1004.260 ;
        RECT 20.310 1004.060 20.630 1004.120 ;
        RECT 2718.210 1004.060 2718.530 1004.120 ;
      LAYER via ;
        RECT 20.340 1004.060 20.600 1004.320 ;
        RECT 2718.240 1004.060 2718.500 1004.320 ;
      LAYER met2 ;
        RECT 2718.230 2267.955 2718.510 2268.325 ;
        RECT 2718.300 1004.350 2718.440 2267.955 ;
        RECT 20.340 1004.030 20.600 1004.350 ;
        RECT 2718.240 1004.030 2718.500 1004.350 ;
        RECT 20.400 969.525 20.540 1004.030 ;
        RECT 20.330 969.155 20.610 969.525 ;
      LAYER via2 ;
        RECT 2718.230 2268.000 2718.510 2268.280 ;
        RECT 20.330 969.200 20.610 969.480 ;
      LAYER met3 ;
        RECT 2718.205 2268.290 2718.535 2268.305 ;
        RECT 2699.740 2268.240 2718.535 2268.290 ;
        RECT 2696.000 2267.990 2718.535 2268.240 ;
        RECT 2696.000 2267.640 2700.000 2267.990 ;
        RECT 2718.205 2267.975 2718.535 2267.990 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 20.305 969.490 20.635 969.505 ;
        RECT -4.800 969.190 20.635 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 20.305 969.175 20.635 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 18.950 1003.835 19.230 1004.205 ;
        RECT 19.020 753.965 19.160 1003.835 ;
        RECT 18.950 753.595 19.230 753.965 ;
      LAYER via2 ;
        RECT 18.950 1003.880 19.230 1004.160 ;
        RECT 18.950 753.640 19.230 753.920 ;
      LAYER met3 ;
        RECT 2715.190 2300.250 2715.570 2300.260 ;
        RECT 2699.740 2300.200 2715.570 2300.250 ;
        RECT 2696.000 2299.950 2715.570 2300.200 ;
        RECT 2696.000 2299.600 2700.000 2299.950 ;
        RECT 2715.190 2299.940 2715.570 2299.950 ;
        RECT 18.925 1004.170 19.255 1004.185 ;
        RECT 2715.190 1004.170 2715.570 1004.180 ;
        RECT 18.925 1003.870 2715.570 1004.170 ;
        RECT 18.925 1003.855 19.255 1003.870 ;
        RECT 2715.190 1003.860 2715.570 1003.870 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 18.925 753.930 19.255 753.945 ;
        RECT -4.800 753.630 19.255 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 18.925 753.615 19.255 753.630 ;
      LAYER via3 ;
        RECT 2715.220 2299.940 2715.540 2300.260 ;
        RECT 2715.220 1003.860 2715.540 1004.180 ;
      LAYER met4 ;
        RECT 2715.215 2299.935 2715.545 2300.265 ;
        RECT 2715.230 1004.185 2715.530 2299.935 ;
        RECT 2715.215 1003.855 2715.545 1004.185 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 544.920 16.490 544.980 ;
        RECT 2711.310 544.920 2711.630 544.980 ;
        RECT 16.170 544.780 2711.630 544.920 ;
        RECT 16.170 544.720 16.490 544.780 ;
        RECT 2711.310 544.720 2711.630 544.780 ;
      LAYER via ;
        RECT 16.200 544.720 16.460 544.980 ;
        RECT 2711.340 544.720 2711.600 544.980 ;
      LAYER met2 ;
        RECT 2711.330 2331.195 2711.610 2331.565 ;
        RECT 2711.400 545.010 2711.540 2331.195 ;
        RECT 16.200 544.690 16.460 545.010 ;
        RECT 2711.340 544.690 2711.600 545.010 ;
        RECT 16.260 538.405 16.400 544.690 ;
        RECT 16.190 538.035 16.470 538.405 ;
      LAYER via2 ;
        RECT 2711.330 2331.240 2711.610 2331.520 ;
        RECT 16.190 538.080 16.470 538.360 ;
      LAYER met3 ;
        RECT 2711.305 2331.530 2711.635 2331.545 ;
        RECT 2699.740 2331.480 2711.635 2331.530 ;
        RECT 2696.000 2331.230 2711.635 2331.480 ;
        RECT 2696.000 2330.880 2700.000 2331.230 ;
        RECT 2711.305 2331.215 2711.635 2331.230 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 16.165 538.370 16.495 538.385 ;
        RECT -4.800 538.070 16.495 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 16.165 538.055 16.495 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2707.830 2363.490 2708.210 2363.500 ;
        RECT 2699.740 2363.440 2708.210 2363.490 ;
        RECT 2696.000 2363.190 2708.210 2363.440 ;
        RECT 2696.000 2362.840 2700.000 2363.190 ;
        RECT 2707.830 2363.180 2708.210 2363.190 ;
        RECT 2707.830 324.170 2708.210 324.180 ;
        RECT 3.070 323.870 2708.210 324.170 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 3.070 322.810 3.370 323.870 ;
        RECT 2707.830 323.860 2708.210 323.870 ;
        RECT -4.800 322.510 3.370 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
      LAYER via3 ;
        RECT 2707.860 2363.180 2708.180 2363.500 ;
        RECT 2707.860 323.860 2708.180 324.180 ;
      LAYER met4 ;
        RECT 2707.855 2363.175 2708.185 2363.505 ;
        RECT 2707.870 324.185 2708.170 2363.175 ;
        RECT 2707.855 323.855 2708.185 324.185 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2712.430 2394.770 2712.810 2394.780 ;
        RECT 2699.740 2394.720 2712.810 2394.770 ;
        RECT 2696.000 2394.470 2712.810 2394.720 ;
        RECT 2696.000 2394.120 2700.000 2394.470 ;
        RECT 2712.430 2394.460 2712.810 2394.470 ;
        RECT 2712.430 109.970 2712.810 109.980 ;
        RECT 3.070 109.670 2712.810 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 2712.430 109.660 2712.810 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 2712.460 2394.460 2712.780 2394.780 ;
        RECT 2712.460 109.660 2712.780 109.980 ;
      LAYER met4 ;
        RECT 2712.455 2394.455 2712.785 2394.785 ;
        RECT 2712.470 109.985 2712.770 2394.455 ;
        RECT 2712.455 109.655 2712.785 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2721.890 855.340 2722.210 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2721.890 855.200 2901.150 855.340 ;
        RECT 2721.890 855.140 2722.210 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2721.920 855.140 2722.180 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 2721.910 1320.715 2722.190 1321.085 ;
        RECT 2721.980 855.430 2722.120 1320.715 ;
        RECT 2721.920 855.110 2722.180 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 2721.910 1320.760 2722.190 1321.040 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 2721.885 1321.050 2722.215 1321.065 ;
        RECT 2699.740 1321.000 2722.215 1321.050 ;
        RECT 2696.000 1320.750 2722.215 1321.000 ;
        RECT 2696.000 1320.400 2700.000 1320.750 ;
        RECT 2721.885 1320.735 2722.215 1320.750 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2717.290 1089.940 2717.610 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 2717.290 1089.800 2901.150 1089.940 ;
        RECT 2717.290 1089.740 2717.610 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 2717.320 1089.740 2717.580 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 2717.310 1351.995 2717.590 1352.365 ;
        RECT 2717.380 1090.030 2717.520 1351.995 ;
        RECT 2717.320 1089.710 2717.580 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 2717.310 1352.040 2717.590 1352.320 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 2717.285 1352.330 2717.615 1352.345 ;
        RECT 2699.740 1352.280 2717.615 1352.330 ;
        RECT 2696.000 1352.030 2717.615 1352.280 ;
        RECT 2696.000 1351.680 2700.000 1352.030 ;
        RECT 2717.285 1352.015 2717.615 1352.030 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2715.450 1324.540 2715.770 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 2715.450 1324.400 2901.150 1324.540 ;
        RECT 2715.450 1324.340 2715.770 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 2715.480 1324.340 2715.740 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 2715.470 1383.955 2715.750 1384.325 ;
        RECT 2715.540 1324.630 2715.680 1383.955 ;
        RECT 2715.480 1324.310 2715.740 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 2715.470 1384.000 2715.750 1384.280 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 2715.445 1384.290 2715.775 1384.305 ;
        RECT 2699.740 1384.240 2715.775 1384.290 ;
        RECT 2696.000 1383.990 2715.775 1384.240 ;
        RECT 2696.000 1383.640 2700.000 1383.990 ;
        RECT 2715.445 1383.975 2715.775 1383.990 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1421.440 2713.470 1421.500 ;
        RECT 2903.130 1421.440 2903.450 1421.500 ;
        RECT 2713.150 1421.300 2903.450 1421.440 ;
        RECT 2713.150 1421.240 2713.470 1421.300 ;
        RECT 2903.130 1421.240 2903.450 1421.300 ;
      LAYER via ;
        RECT 2713.180 1421.240 2713.440 1421.500 ;
        RECT 2903.160 1421.240 2903.420 1421.500 ;
      LAYER met2 ;
        RECT 2903.150 1553.955 2903.430 1554.325 ;
        RECT 2903.220 1421.530 2903.360 1553.955 ;
        RECT 2713.180 1421.210 2713.440 1421.530 ;
        RECT 2903.160 1421.210 2903.420 1421.530 ;
        RECT 2713.240 1415.605 2713.380 1421.210 ;
        RECT 2713.170 1415.235 2713.450 1415.605 ;
      LAYER via2 ;
        RECT 2903.150 1554.000 2903.430 1554.280 ;
        RECT 2713.170 1415.280 2713.450 1415.560 ;
      LAYER met3 ;
        RECT 2903.125 1554.290 2903.455 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2903.125 1553.990 2924.800 1554.290 ;
        RECT 2903.125 1553.975 2903.455 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 2713.145 1415.570 2713.475 1415.585 ;
        RECT 2699.740 1415.520 2713.475 1415.570 ;
        RECT 2696.000 1415.270 2713.475 1415.520 ;
        RECT 2696.000 1414.920 2700.000 1415.270 ;
        RECT 2713.145 1415.255 2713.475 1415.270 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2713.150 1448.980 2713.470 1449.040 ;
        RECT 2901.750 1448.980 2902.070 1449.040 ;
        RECT 2713.150 1448.840 2902.070 1448.980 ;
        RECT 2713.150 1448.780 2713.470 1448.840 ;
        RECT 2901.750 1448.780 2902.070 1448.840 ;
      LAYER via ;
        RECT 2713.180 1448.780 2713.440 1449.040 ;
        RECT 2901.780 1448.780 2902.040 1449.040 ;
      LAYER met2 ;
        RECT 2901.770 1789.235 2902.050 1789.605 ;
        RECT 2901.840 1449.070 2901.980 1789.235 ;
        RECT 2713.180 1448.750 2713.440 1449.070 ;
        RECT 2901.780 1448.750 2902.040 1449.070 ;
        RECT 2713.240 1447.565 2713.380 1448.750 ;
        RECT 2713.170 1447.195 2713.450 1447.565 ;
      LAYER via2 ;
        RECT 2901.770 1789.280 2902.050 1789.560 ;
        RECT 2713.170 1447.240 2713.450 1447.520 ;
      LAYER met3 ;
        RECT 2901.745 1789.570 2902.075 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2901.745 1789.270 2924.800 1789.570 ;
        RECT 2901.745 1789.255 2902.075 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
        RECT 2713.145 1447.530 2713.475 1447.545 ;
        RECT 2699.740 1447.480 2713.475 1447.530 ;
        RECT 2696.000 1447.230 2713.475 1447.480 ;
        RECT 2696.000 1446.880 2700.000 1447.230 ;
        RECT 2713.145 1447.215 2713.475 1447.230 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2749.950 2021.880 2750.270 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 2749.950 2021.740 2901.150 2021.880 ;
        RECT 2749.950 2021.680 2750.270 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
        RECT 2713.150 1483.320 2713.470 1483.380 ;
        RECT 2749.950 1483.320 2750.270 1483.380 ;
        RECT 2713.150 1483.180 2750.270 1483.320 ;
        RECT 2713.150 1483.120 2713.470 1483.180 ;
        RECT 2749.950 1483.120 2750.270 1483.180 ;
      LAYER via ;
        RECT 2749.980 2021.680 2750.240 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
        RECT 2713.180 1483.120 2713.440 1483.380 ;
        RECT 2749.980 1483.120 2750.240 1483.380 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 2749.980 2021.650 2750.240 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 2750.040 1483.410 2750.180 2021.650 ;
        RECT 2713.180 1483.090 2713.440 1483.410 ;
        RECT 2749.980 1483.090 2750.240 1483.410 ;
        RECT 2713.240 1478.845 2713.380 1483.090 ;
        RECT 2713.170 1478.475 2713.450 1478.845 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
        RECT 2713.170 1478.520 2713.450 1478.800 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
        RECT 2713.145 1478.810 2713.475 1478.825 ;
        RECT 2699.740 1478.760 2713.475 1478.810 ;
        RECT 2696.000 1478.510 2713.475 1478.760 ;
        RECT 2696.000 1478.160 2700.000 1478.510 ;
        RECT 2713.145 1478.495 2713.475 1478.510 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2818.950 2256.480 2819.270 2256.540 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 2818.950 2256.340 2901.150 2256.480 ;
        RECT 2818.950 2256.280 2819.270 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
        RECT 2713.150 1510.860 2713.470 1510.920 ;
        RECT 2818.950 1510.860 2819.270 1510.920 ;
        RECT 2713.150 1510.720 2819.270 1510.860 ;
        RECT 2713.150 1510.660 2713.470 1510.720 ;
        RECT 2818.950 1510.660 2819.270 1510.720 ;
      LAYER via ;
        RECT 2818.980 2256.280 2819.240 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
        RECT 2713.180 1510.660 2713.440 1510.920 ;
        RECT 2818.980 1510.660 2819.240 1510.920 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 2818.980 2256.250 2819.240 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 2819.040 1510.950 2819.180 2256.250 ;
        RECT 2713.180 1510.630 2713.440 1510.950 ;
        RECT 2818.980 1510.630 2819.240 1510.950 ;
        RECT 2713.240 1510.125 2713.380 1510.630 ;
        RECT 2713.170 1509.755 2713.450 1510.125 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
        RECT 2713.170 1509.800 2713.450 1510.080 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
        RECT 2713.145 1510.090 2713.475 1510.105 ;
        RECT 2699.740 1510.040 2713.475 1510.090 ;
        RECT 2696.000 1509.790 2713.475 1510.040 ;
        RECT 2696.000 1509.440 2700.000 1509.790 ;
        RECT 2713.145 1509.775 2713.475 1509.790 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 634.410 2325.500 634.730 2325.560 ;
        RECT 1283.470 2325.500 1283.790 2325.560 ;
        RECT 634.410 2325.360 1283.790 2325.500 ;
        RECT 634.410 2325.300 634.730 2325.360 ;
        RECT 1283.470 2325.300 1283.790 2325.360 ;
      LAYER via ;
        RECT 634.440 2325.300 634.700 2325.560 ;
        RECT 1283.500 2325.300 1283.760 2325.560 ;
      LAYER met2 ;
        RECT 1283.490 2330.515 1283.770 2330.885 ;
        RECT 1283.560 2325.590 1283.700 2330.515 ;
        RECT 634.440 2325.270 634.700 2325.590 ;
        RECT 1283.500 2325.270 1283.760 2325.590 ;
        RECT 634.500 17.410 634.640 2325.270 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2330.560 1283.770 2330.840 ;
      LAYER met3 ;
        RECT 1283.465 2330.850 1283.795 2330.865 ;
        RECT 1283.465 2330.800 1300.420 2330.850 ;
        RECT 1283.465 2330.550 1304.000 2330.800 ;
        RECT 1283.465 2330.535 1283.795 2330.550 ;
        RECT 1300.000 2330.200 1304.000 2330.550 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 655.110 2360.180 655.430 2360.240 ;
        RECT 1283.470 2360.180 1283.790 2360.240 ;
        RECT 655.110 2360.040 1283.790 2360.180 ;
        RECT 655.110 2359.980 655.430 2360.040 ;
        RECT 1283.470 2359.980 1283.790 2360.040 ;
        RECT 650.970 17.920 651.290 17.980 ;
        RECT 655.110 17.920 655.430 17.980 ;
        RECT 650.970 17.780 655.430 17.920 ;
        RECT 650.970 17.720 651.290 17.780 ;
        RECT 655.110 17.720 655.430 17.780 ;
      LAYER via ;
        RECT 655.140 2359.980 655.400 2360.240 ;
        RECT 1283.500 2359.980 1283.760 2360.240 ;
        RECT 651.000 17.720 651.260 17.980 ;
        RECT 655.140 17.720 655.400 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2362.475 1283.770 2362.845 ;
        RECT 1283.560 2360.270 1283.700 2362.475 ;
        RECT 655.140 2359.950 655.400 2360.270 ;
        RECT 1283.500 2359.950 1283.760 2360.270 ;
        RECT 655.200 18.010 655.340 2359.950 ;
        RECT 651.000 17.690 651.260 18.010 ;
        RECT 655.140 17.690 655.400 18.010 ;
        RECT 651.060 2.400 651.200 17.690 ;
        RECT 650.850 -4.800 651.410 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2362.520 1283.770 2362.800 ;
      LAYER met3 ;
        RECT 1283.465 2362.810 1283.795 2362.825 ;
        RECT 1283.465 2362.760 1300.420 2362.810 ;
        RECT 1283.465 2362.510 1304.000 2362.760 ;
        RECT 1283.465 2362.495 1283.795 2362.510 ;
        RECT 1300.000 2362.160 1304.000 2362.510 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 641.310 2339.440 641.630 2339.500 ;
        RECT 1283.470 2339.440 1283.790 2339.500 ;
        RECT 641.310 2339.300 1283.790 2339.440 ;
        RECT 641.310 2339.240 641.630 2339.300 ;
        RECT 1283.470 2339.240 1283.790 2339.300 ;
        RECT 639.010 17.920 639.330 17.980 ;
        RECT 641.310 17.920 641.630 17.980 ;
        RECT 639.010 17.780 641.630 17.920 ;
        RECT 639.010 17.720 639.330 17.780 ;
        RECT 641.310 17.720 641.630 17.780 ;
      LAYER via ;
        RECT 641.340 2339.240 641.600 2339.500 ;
        RECT 1283.500 2339.240 1283.760 2339.500 ;
        RECT 639.040 17.720 639.300 17.980 ;
        RECT 641.340 17.720 641.600 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2341.395 1283.770 2341.765 ;
        RECT 1283.560 2339.530 1283.700 2341.395 ;
        RECT 641.340 2339.210 641.600 2339.530 ;
        RECT 1283.500 2339.210 1283.760 2339.530 ;
        RECT 641.400 18.010 641.540 2339.210 ;
        RECT 639.040 17.690 639.300 18.010 ;
        RECT 641.340 17.690 641.600 18.010 ;
        RECT 639.100 2.400 639.240 17.690 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2341.440 1283.770 2341.720 ;
      LAYER met3 ;
        RECT 1283.465 2341.730 1283.795 2341.745 ;
        RECT 1283.465 2341.680 1300.420 2341.730 ;
        RECT 1283.465 2341.430 1304.000 2341.680 ;
        RECT 1283.465 2341.415 1283.795 2341.430 ;
        RECT 1300.000 2341.080 1304.000 2341.430 ;
    END
  END la_data_out[0]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 662.010 2366.980 662.330 2367.040 ;
        RECT 1283.470 2366.980 1283.790 2367.040 ;
        RECT 662.010 2366.840 1283.790 2366.980 ;
        RECT 662.010 2366.780 662.330 2366.840 ;
        RECT 1283.470 2366.780 1283.790 2366.840 ;
        RECT 656.950 17.920 657.270 17.980 ;
        RECT 662.010 17.920 662.330 17.980 ;
        RECT 656.950 17.780 662.330 17.920 ;
        RECT 656.950 17.720 657.270 17.780 ;
        RECT 662.010 17.720 662.330 17.780 ;
      LAYER via ;
        RECT 662.040 2366.780 662.300 2367.040 ;
        RECT 1283.500 2366.780 1283.760 2367.040 ;
        RECT 656.980 17.720 657.240 17.980 ;
        RECT 662.040 17.720 662.300 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2373.355 1283.770 2373.725 ;
        RECT 1283.560 2367.070 1283.700 2373.355 ;
        RECT 662.040 2366.750 662.300 2367.070 ;
        RECT 1283.500 2366.750 1283.760 2367.070 ;
        RECT 662.100 18.010 662.240 2366.750 ;
        RECT 656.980 17.690 657.240 18.010 ;
        RECT 662.040 17.690 662.300 18.010 ;
        RECT 657.040 2.400 657.180 17.690 ;
        RECT 656.830 -4.800 657.390 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2373.400 1283.770 2373.680 ;
      LAYER met3 ;
        RECT 1283.465 2373.690 1283.795 2373.705 ;
        RECT 1283.465 2373.640 1300.420 2373.690 ;
        RECT 1283.465 2373.390 1304.000 2373.640 ;
        RECT 1283.465 2373.375 1283.795 2373.390 ;
        RECT 1300.000 2373.040 1304.000 2373.390 ;
    END
  END la_data_out[1]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 675.810 2394.520 676.130 2394.580 ;
        RECT 1283.470 2394.520 1283.790 2394.580 ;
        RECT 675.810 2394.380 1283.790 2394.520 ;
        RECT 675.810 2394.320 676.130 2394.380 ;
        RECT 1283.470 2394.320 1283.790 2394.380 ;
      LAYER via ;
        RECT 675.840 2394.320 676.100 2394.580 ;
        RECT 1283.500 2394.320 1283.760 2394.580 ;
      LAYER met2 ;
        RECT 675.840 2394.290 676.100 2394.610 ;
        RECT 1283.490 2394.435 1283.770 2394.805 ;
        RECT 1283.500 2394.290 1283.760 2394.435 ;
        RECT 675.900 3.130 676.040 2394.290 ;
        RECT 674.520 2.990 676.040 3.130 ;
        RECT 674.520 2.400 674.660 2.990 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2394.480 1283.770 2394.760 ;
      LAYER met3 ;
        RECT 1283.465 2394.770 1283.795 2394.785 ;
        RECT 1283.465 2394.720 1300.420 2394.770 ;
        RECT 1283.465 2394.470 1304.000 2394.720 ;
        RECT 1283.465 2394.455 1283.795 2394.470 ;
        RECT 1300.000 2394.120 1304.000 2394.470 ;
    END
  END la_data_out[2]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 2346.240 648.530 2346.300 ;
        RECT 1283.470 2346.240 1283.790 2346.300 ;
        RECT 648.210 2346.100 1283.790 2346.240 ;
        RECT 648.210 2346.040 648.530 2346.100 ;
        RECT 1283.470 2346.040 1283.790 2346.100 ;
        RECT 644.990 17.920 645.310 17.980 ;
        RECT 648.210 17.920 648.530 17.980 ;
        RECT 644.990 17.780 648.530 17.920 ;
        RECT 644.990 17.720 645.310 17.780 ;
        RECT 648.210 17.720 648.530 17.780 ;
      LAYER via ;
        RECT 648.240 2346.040 648.500 2346.300 ;
        RECT 1283.500 2346.040 1283.760 2346.300 ;
        RECT 645.020 17.720 645.280 17.980 ;
        RECT 648.240 17.720 648.500 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2351.595 1283.770 2351.965 ;
        RECT 1283.560 2346.330 1283.700 2351.595 ;
        RECT 648.240 2346.010 648.500 2346.330 ;
        RECT 1283.500 2346.010 1283.760 2346.330 ;
        RECT 648.300 18.010 648.440 2346.010 ;
        RECT 645.020 17.690 645.280 18.010 ;
        RECT 648.240 17.690 648.500 18.010 ;
        RECT 645.080 2.400 645.220 17.690 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2351.640 1283.770 2351.920 ;
      LAYER met3 ;
        RECT 1283.465 2351.930 1283.795 2351.945 ;
        RECT 1283.465 2351.880 1300.420 2351.930 ;
        RECT 1283.465 2351.630 1304.000 2351.880 ;
        RECT 1283.465 2351.615 1283.795 2351.630 ;
        RECT 1300.000 2351.280 1304.000 2351.630 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 2380.580 669.230 2380.640 ;
        RECT 1283.470 2380.580 1283.790 2380.640 ;
        RECT 668.910 2380.440 1283.790 2380.580 ;
        RECT 668.910 2380.380 669.230 2380.440 ;
        RECT 1283.470 2380.380 1283.790 2380.440 ;
        RECT 662.930 17.920 663.250 17.980 ;
        RECT 668.910 17.920 669.230 17.980 ;
        RECT 662.930 17.780 669.230 17.920 ;
        RECT 662.930 17.720 663.250 17.780 ;
        RECT 668.910 17.720 669.230 17.780 ;
      LAYER via ;
        RECT 668.940 2380.380 669.200 2380.640 ;
        RECT 1283.500 2380.380 1283.760 2380.640 ;
        RECT 662.960 17.720 663.220 17.980 ;
        RECT 668.940 17.720 669.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2383.555 1283.770 2383.925 ;
        RECT 1283.560 2380.670 1283.700 2383.555 ;
        RECT 668.940 2380.350 669.200 2380.670 ;
        RECT 1283.500 2380.350 1283.760 2380.670 ;
        RECT 669.000 18.010 669.140 2380.350 ;
        RECT 662.960 17.690 663.220 18.010 ;
        RECT 668.940 17.690 669.200 18.010 ;
        RECT 663.020 2.400 663.160 17.690 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2383.600 1283.770 2383.880 ;
      LAYER met3 ;
        RECT 1283.465 2383.890 1283.795 2383.905 ;
        RECT 1283.465 2383.840 1300.420 2383.890 ;
        RECT 1283.465 2383.590 1304.000 2383.840 ;
        RECT 1283.465 2383.575 1283.795 2383.590 ;
        RECT 1300.000 2383.240 1304.000 2383.590 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1518.070 2591.040 1518.390 2591.100 ;
        RECT 2118.370 2591.040 2118.690 2591.100 ;
        RECT 1518.070 2590.900 2118.690 2591.040 ;
        RECT 1518.070 2590.840 1518.390 2590.900 ;
        RECT 2118.370 2590.840 2118.690 2590.900 ;
        RECT 1305.550 2588.320 1305.870 2588.380 ;
        RECT 1518.070 2588.320 1518.390 2588.380 ;
        RECT 1305.550 2588.180 1518.390 2588.320 ;
        RECT 1305.550 2588.120 1305.870 2588.180 ;
        RECT 1518.070 2588.120 1518.390 2588.180 ;
        RECT 1414.200 1204.720 1449.300 1204.860 ;
        RECT 1414.200 1203.500 1414.340 1204.720 ;
        RECT 1449.160 1203.560 1449.300 1204.720 ;
        RECT 1558.640 1204.380 1594.200 1204.520 ;
        RECT 1558.640 1204.180 1558.780 1204.380 ;
        RECT 1497.000 1204.040 1558.780 1204.180 ;
        RECT 1497.000 1203.560 1497.140 1204.040 ;
        RECT 1594.060 1203.560 1594.200 1204.380 ;
        RECT 1641.900 1204.040 1656.300 1204.180 ;
        RECT 1641.900 1203.560 1642.040 1204.040 ;
        RECT 1656.160 1203.840 1656.300 1204.040 ;
        RECT 1656.160 1203.700 1657.220 1203.840 ;
        RECT 1400.400 1203.360 1414.340 1203.500 ;
        RECT 1352.010 1203.160 1352.330 1203.220 ;
        RECT 1366.270 1203.160 1366.590 1203.220 ;
        RECT 1352.010 1203.020 1366.590 1203.160 ;
        RECT 1352.010 1202.960 1352.330 1203.020 ;
        RECT 1366.270 1202.960 1366.590 1203.020 ;
        RECT 1366.730 1203.160 1367.050 1203.220 ;
        RECT 1400.400 1203.160 1400.540 1203.360 ;
        RECT 1449.070 1203.300 1449.390 1203.560 ;
        RECT 1496.910 1203.300 1497.230 1203.560 ;
        RECT 1593.970 1203.300 1594.290 1203.560 ;
        RECT 1641.810 1203.300 1642.130 1203.560 ;
        RECT 1657.080 1203.500 1657.220 1203.700 ;
        RECT 1738.960 1203.700 1787.400 1203.840 ;
        RECT 1738.960 1203.500 1739.100 1203.700 ;
        RECT 1787.260 1203.560 1787.400 1203.700 ;
        RECT 1657.080 1203.360 1739.100 1203.500 ;
        RECT 1787.170 1203.300 1787.490 1203.560 ;
        RECT 1835.010 1203.500 1835.330 1203.560 ;
        RECT 1840.070 1203.500 1840.390 1203.560 ;
        RECT 1835.010 1203.360 1840.390 1203.500 ;
        RECT 1835.010 1203.300 1835.330 1203.360 ;
        RECT 1840.070 1203.300 1840.390 1203.360 ;
        RECT 1366.730 1203.020 1400.540 1203.160 ;
        RECT 1366.730 1202.960 1367.050 1203.020 ;
        RECT 1289.910 1202.820 1290.230 1202.880 ;
        RECT 1304.170 1202.820 1304.490 1202.880 ;
        RECT 1289.910 1202.680 1304.490 1202.820 ;
        RECT 1289.910 1202.620 1290.230 1202.680 ;
        RECT 1304.170 1202.620 1304.490 1202.680 ;
        RECT 1449.070 1202.820 1449.390 1202.880 ;
        RECT 1496.910 1202.820 1497.230 1202.880 ;
        RECT 1449.070 1202.680 1497.230 1202.820 ;
        RECT 1449.070 1202.620 1449.390 1202.680 ;
        RECT 1496.910 1202.620 1497.230 1202.680 ;
        RECT 1593.970 1202.820 1594.290 1202.880 ;
        RECT 1641.810 1202.820 1642.130 1202.880 ;
        RECT 1593.970 1202.680 1642.130 1202.820 ;
        RECT 1593.970 1202.620 1594.290 1202.680 ;
        RECT 1641.810 1202.620 1642.130 1202.680 ;
        RECT 1304.170 1202.140 1304.490 1202.200 ;
        RECT 1305.550 1202.140 1305.870 1202.200 ;
        RECT 1352.010 1202.140 1352.330 1202.200 ;
        RECT 1304.170 1202.000 1352.330 1202.140 ;
        RECT 1304.170 1201.940 1304.490 1202.000 ;
        RECT 1305.550 1201.940 1305.870 1202.000 ;
        RECT 1352.010 1201.940 1352.330 1202.000 ;
        RECT 6.510 1200.780 6.830 1200.840 ;
        RECT 1289.910 1200.780 1290.230 1200.840 ;
        RECT 6.510 1200.640 1290.230 1200.780 ;
        RECT 6.510 1200.580 6.830 1200.640 ;
        RECT 1289.910 1200.580 1290.230 1200.640 ;
        RECT 1840.070 1200.440 1840.390 1200.500 ;
        RECT 1866.290 1200.440 1866.610 1200.500 ;
        RECT 1840.070 1200.300 1866.610 1200.440 ;
        RECT 1840.070 1200.240 1840.390 1200.300 ;
        RECT 1866.290 1200.240 1866.610 1200.300 ;
        RECT 2.830 17.580 3.150 17.640 ;
        RECT 6.510 17.580 6.830 17.640 ;
        RECT 2.830 17.440 6.830 17.580 ;
        RECT 2.830 17.380 3.150 17.440 ;
        RECT 6.510 17.380 6.830 17.440 ;
      LAYER via ;
        RECT 1518.100 2590.840 1518.360 2591.100 ;
        RECT 2118.400 2590.840 2118.660 2591.100 ;
        RECT 1305.580 2588.120 1305.840 2588.380 ;
        RECT 1518.100 2588.120 1518.360 2588.380 ;
        RECT 1352.040 1202.960 1352.300 1203.220 ;
        RECT 1366.300 1202.960 1366.560 1203.220 ;
        RECT 1366.760 1202.960 1367.020 1203.220 ;
        RECT 1449.100 1203.300 1449.360 1203.560 ;
        RECT 1496.940 1203.300 1497.200 1203.560 ;
        RECT 1594.000 1203.300 1594.260 1203.560 ;
        RECT 1641.840 1203.300 1642.100 1203.560 ;
        RECT 1787.200 1203.300 1787.460 1203.560 ;
        RECT 1835.040 1203.300 1835.300 1203.560 ;
        RECT 1840.100 1203.300 1840.360 1203.560 ;
        RECT 1289.940 1202.620 1290.200 1202.880 ;
        RECT 1304.200 1202.620 1304.460 1202.880 ;
        RECT 1449.100 1202.620 1449.360 1202.880 ;
        RECT 1496.940 1202.620 1497.200 1202.880 ;
        RECT 1594.000 1202.620 1594.260 1202.880 ;
        RECT 1641.840 1202.620 1642.100 1202.880 ;
        RECT 1304.200 1201.940 1304.460 1202.200 ;
        RECT 1305.580 1201.940 1305.840 1202.200 ;
        RECT 1352.040 1201.940 1352.300 1202.200 ;
        RECT 6.540 1200.580 6.800 1200.840 ;
        RECT 1289.940 1200.580 1290.200 1200.840 ;
        RECT 1840.100 1200.240 1840.360 1200.500 ;
        RECT 1866.320 1200.240 1866.580 1200.500 ;
        RECT 2.860 17.380 3.120 17.640 ;
        RECT 6.540 17.380 6.800 17.640 ;
      LAYER met2 ;
        RECT 1518.090 2590.955 1518.370 2591.325 ;
        RECT 2118.390 2590.955 2118.670 2591.325 ;
        RECT 1518.100 2590.810 1518.360 2590.955 ;
        RECT 2118.400 2590.810 2118.660 2590.955 ;
        RECT 1518.160 2588.410 1518.300 2590.810 ;
        RECT 1305.580 2588.090 1305.840 2588.410 ;
        RECT 1518.100 2588.090 1518.360 2588.410 ;
        RECT 1289.930 1205.115 1290.210 1205.485 ;
        RECT 1290.000 1202.910 1290.140 1205.115 ;
        RECT 1289.940 1202.590 1290.200 1202.910 ;
        RECT 1304.200 1202.590 1304.460 1202.910 ;
        RECT 1290.000 1200.870 1290.140 1202.590 ;
        RECT 1304.260 1202.230 1304.400 1202.590 ;
        RECT 1305.640 1202.230 1305.780 2588.090 ;
        RECT 1366.360 1203.250 1366.960 1203.330 ;
        RECT 1449.100 1203.270 1449.360 1203.590 ;
        RECT 1496.940 1203.270 1497.200 1203.590 ;
        RECT 1594.000 1203.270 1594.260 1203.590 ;
        RECT 1641.840 1203.270 1642.100 1203.590 ;
        RECT 1787.200 1203.445 1787.460 1203.590 ;
        RECT 1352.040 1202.930 1352.300 1203.250 ;
        RECT 1366.300 1203.190 1367.020 1203.250 ;
        RECT 1366.300 1202.930 1366.560 1203.190 ;
        RECT 1366.760 1202.930 1367.020 1203.190 ;
        RECT 1352.100 1202.230 1352.240 1202.930 ;
        RECT 1449.160 1202.910 1449.300 1203.270 ;
        RECT 1497.000 1202.910 1497.140 1203.270 ;
        RECT 1594.060 1202.910 1594.200 1203.270 ;
        RECT 1641.900 1202.910 1642.040 1203.270 ;
        RECT 1787.190 1203.075 1787.470 1203.445 ;
        RECT 1834.570 1203.330 1834.850 1203.445 ;
        RECT 1835.040 1203.330 1835.300 1203.590 ;
        RECT 1834.570 1203.270 1835.300 1203.330 ;
        RECT 1840.100 1203.270 1840.360 1203.590 ;
        RECT 1834.570 1203.190 1835.240 1203.270 ;
        RECT 1834.570 1203.075 1834.850 1203.190 ;
        RECT 1449.100 1202.590 1449.360 1202.910 ;
        RECT 1496.940 1202.590 1497.200 1202.910 ;
        RECT 1594.000 1202.590 1594.260 1202.910 ;
        RECT 1641.840 1202.590 1642.100 1202.910 ;
        RECT 1304.200 1201.910 1304.460 1202.230 ;
        RECT 1305.580 1201.910 1305.840 1202.230 ;
        RECT 1352.040 1201.910 1352.300 1202.230 ;
        RECT 6.540 1200.550 6.800 1200.870 ;
        RECT 1289.940 1200.550 1290.200 1200.870 ;
        RECT 6.600 17.670 6.740 1200.550 ;
        RECT 1840.160 1200.530 1840.300 1203.270 ;
        RECT 1840.100 1200.210 1840.360 1200.530 ;
        RECT 1866.320 1200.210 1866.580 1200.530 ;
        RECT 1866.380 1015.765 1866.520 1200.210 ;
        RECT 1866.310 1015.395 1866.590 1015.765 ;
        RECT 2.860 17.350 3.120 17.670 ;
        RECT 6.540 17.350 6.800 17.670 ;
        RECT 2.920 2.400 3.060 17.350 ;
        RECT 2.710 -4.800 3.270 2.400 ;
      LAYER via2 ;
        RECT 1518.090 2591.000 1518.370 2591.280 ;
        RECT 2118.390 2591.000 2118.670 2591.280 ;
        RECT 1289.930 1205.160 1290.210 1205.440 ;
        RECT 1787.190 1203.120 1787.470 1203.400 ;
        RECT 1834.570 1203.120 1834.850 1203.400 ;
        RECT 1866.310 1015.440 1866.590 1015.720 ;
      LAYER met3 ;
        RECT 1518.065 2591.300 1518.395 2591.305 ;
        RECT 1518.065 2591.290 1518.650 2591.300 ;
        RECT 2118.365 2591.290 2118.695 2591.305 ;
        RECT 2119.030 2591.290 2119.410 2591.300 ;
        RECT 1518.065 2590.990 1518.850 2591.290 ;
        RECT 2118.365 2590.990 2119.410 2591.290 ;
        RECT 1518.065 2590.980 1518.650 2590.990 ;
        RECT 1518.065 2590.975 1518.395 2590.980 ;
        RECT 2118.365 2590.975 2118.695 2590.990 ;
        RECT 2119.030 2590.980 2119.410 2590.990 ;
        RECT 1289.905 1205.450 1290.235 1205.465 ;
        RECT 1289.905 1205.400 1300.420 1205.450 ;
        RECT 1289.905 1205.150 1304.000 1205.400 ;
        RECT 1289.905 1205.135 1290.235 1205.150 ;
        RECT 1300.000 1204.800 1304.000 1205.150 ;
        RECT 1787.165 1203.410 1787.495 1203.425 ;
        RECT 1834.545 1203.410 1834.875 1203.425 ;
        RECT 1787.165 1203.110 1834.875 1203.410 ;
        RECT 1787.165 1203.095 1787.495 1203.110 ;
        RECT 1834.545 1203.095 1834.875 1203.110 ;
        RECT 1866.285 1015.730 1866.615 1015.745 ;
        RECT 1866.950 1015.730 1867.330 1015.740 ;
        RECT 2464.030 1015.730 2464.410 1015.740 ;
        RECT 1866.285 1015.430 2464.410 1015.730 ;
        RECT 1866.285 1015.415 1866.615 1015.430 ;
        RECT 1866.950 1015.420 1867.330 1015.430 ;
        RECT 2464.030 1015.420 2464.410 1015.430 ;
      LAYER via3 ;
        RECT 1518.300 2590.980 1518.620 2591.300 ;
        RECT 2119.060 2590.980 2119.380 2591.300 ;
        RECT 1866.980 1015.420 1867.300 1015.740 ;
        RECT 2464.060 1015.420 2464.380 1015.740 ;
      LAYER met4 ;
        RECT 1519.015 2601.150 1519.315 2604.600 ;
        RECT 1518.310 2600.850 1519.315 2601.150 ;
        RECT 1518.310 2591.305 1518.610 2600.850 ;
        RECT 1519.015 2600.000 1519.315 2600.850 ;
        RECT 2119.015 2601.150 2119.315 2604.600 ;
        RECT 2119.015 2600.000 2119.370 2601.150 ;
        RECT 2119.070 2591.305 2119.370 2600.000 ;
        RECT 1518.295 2590.975 1518.625 2591.305 ;
        RECT 2119.055 2590.975 2119.385 2591.305 ;
        RECT 1866.975 1015.415 1867.305 1015.745 ;
        RECT 2464.055 1015.415 2464.385 1015.745 ;
        RECT 1866.990 1006.235 1867.290 1015.415 ;
        RECT 1866.990 1004.550 1867.465 1006.235 ;
        RECT 2464.070 1004.850 2464.370 1015.415 ;
        RECT 2467.165 1004.850 2467.465 1006.235 ;
        RECT 2464.070 1004.550 2467.465 1004.850 ;
        RECT 1867.165 1001.635 1867.465 1004.550 ;
        RECT 2467.165 1001.635 2467.465 1004.550 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 13.410 1214.720 13.730 1214.780 ;
        RECT 1284.850 1214.720 1285.170 1214.780 ;
        RECT 13.410 1214.580 1285.170 1214.720 ;
        RECT 13.410 1214.520 13.730 1214.580 ;
        RECT 1284.850 1214.520 1285.170 1214.580 ;
        RECT 8.350 17.580 8.670 17.640 ;
        RECT 13.410 17.580 13.730 17.640 ;
        RECT 8.350 17.440 13.730 17.580 ;
        RECT 8.350 17.380 8.670 17.440 ;
        RECT 13.410 17.380 13.730 17.440 ;
      LAYER via ;
        RECT 13.440 1214.520 13.700 1214.780 ;
        RECT 1284.880 1214.520 1285.140 1214.780 ;
        RECT 8.380 17.380 8.640 17.640 ;
        RECT 13.440 17.380 13.700 17.640 ;
      LAYER met2 ;
        RECT 1284.870 1215.315 1285.150 1215.685 ;
        RECT 1284.940 1214.810 1285.080 1215.315 ;
        RECT 13.440 1214.490 13.700 1214.810 ;
        RECT 1284.880 1214.490 1285.140 1214.810 ;
        RECT 13.500 17.670 13.640 1214.490 ;
        RECT 8.380 17.350 8.640 17.670 ;
        RECT 13.440 17.350 13.700 17.670 ;
        RECT 8.440 2.400 8.580 17.350 ;
        RECT 8.230 -4.800 8.790 2.400 ;
      LAYER via2 ;
        RECT 1284.870 1215.360 1285.150 1215.640 ;
      LAYER met3 ;
        RECT 1284.845 1215.650 1285.175 1215.665 ;
        RECT 1284.845 1215.600 1300.420 1215.650 ;
        RECT 1284.845 1215.350 1304.000 1215.600 ;
        RECT 1284.845 1215.335 1285.175 1215.350 ;
        RECT 1300.000 1215.000 1304.000 1215.350 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.330 17.580 14.650 17.640 ;
        RECT 1287.150 17.580 1287.470 17.640 ;
        RECT 14.330 17.440 1287.470 17.580 ;
        RECT 14.330 17.380 14.650 17.440 ;
        RECT 1287.150 17.380 1287.470 17.440 ;
      LAYER via ;
        RECT 14.360 17.380 14.620 17.640 ;
        RECT 1287.180 17.380 1287.440 17.640 ;
      LAYER met2 ;
        RECT 1287.170 1226.195 1287.450 1226.565 ;
        RECT 1287.240 17.670 1287.380 1226.195 ;
        RECT 14.360 17.350 14.620 17.670 ;
        RECT 1287.180 17.350 1287.440 17.670 ;
        RECT 14.420 2.400 14.560 17.350 ;
        RECT 14.210 -4.800 14.770 2.400 ;
      LAYER via2 ;
        RECT 1287.170 1226.240 1287.450 1226.520 ;
      LAYER met3 ;
        RECT 1287.145 1226.530 1287.475 1226.545 ;
        RECT 1287.145 1226.480 1300.420 1226.530 ;
        RECT 1287.145 1226.230 1304.000 1226.480 ;
        RECT 1287.145 1226.215 1287.475 1226.230 ;
        RECT 1300.000 1225.880 1304.000 1226.230 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 41.010 1263.000 41.330 1263.060 ;
        RECT 1283.470 1263.000 1283.790 1263.060 ;
        RECT 41.010 1262.860 1283.790 1263.000 ;
        RECT 41.010 1262.800 41.330 1262.860 ;
        RECT 1283.470 1262.800 1283.790 1262.860 ;
        RECT 38.250 17.920 38.570 17.980 ;
        RECT 41.010 17.920 41.330 17.980 ;
        RECT 38.250 17.780 41.330 17.920 ;
        RECT 38.250 17.720 38.570 17.780 ;
        RECT 41.010 17.720 41.330 17.780 ;
      LAYER via ;
        RECT 41.040 1262.800 41.300 1263.060 ;
        RECT 1283.500 1262.800 1283.760 1263.060 ;
        RECT 38.280 17.720 38.540 17.980 ;
        RECT 41.040 17.720 41.300 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1268.355 1283.770 1268.725 ;
        RECT 1283.560 1263.090 1283.700 1268.355 ;
        RECT 41.040 1262.770 41.300 1263.090 ;
        RECT 1283.500 1262.770 1283.760 1263.090 ;
        RECT 41.100 18.010 41.240 1262.770 ;
        RECT 38.280 17.690 38.540 18.010 ;
        RECT 41.040 17.690 41.300 18.010 ;
        RECT 38.340 2.400 38.480 17.690 ;
        RECT 38.130 -4.800 38.690 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1268.400 1283.770 1268.680 ;
      LAYER met3 ;
        RECT 1283.465 1268.690 1283.795 1268.705 ;
        RECT 1283.465 1268.640 1300.420 1268.690 ;
        RECT 1283.465 1268.390 1304.000 1268.640 ;
        RECT 1283.465 1268.375 1283.795 1268.390 ;
        RECT 1300.000 1268.040 1304.000 1268.390 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 241.110 1628.500 241.430 1628.560 ;
        RECT 1283.470 1628.500 1283.790 1628.560 ;
        RECT 241.110 1628.360 1283.790 1628.500 ;
        RECT 241.110 1628.300 241.430 1628.360 ;
        RECT 1283.470 1628.300 1283.790 1628.360 ;
        RECT 241.110 468.560 241.430 468.820 ;
        RECT 241.200 467.800 241.340 468.560 ;
        RECT 241.110 467.540 241.430 467.800 ;
      LAYER via ;
        RECT 241.140 1628.300 241.400 1628.560 ;
        RECT 1283.500 1628.300 1283.760 1628.560 ;
        RECT 241.140 468.560 241.400 468.820 ;
        RECT 241.140 467.540 241.400 467.800 ;
      LAYER met2 ;
        RECT 1283.490 1629.435 1283.770 1629.805 ;
        RECT 1283.560 1628.590 1283.700 1629.435 ;
        RECT 241.140 1628.270 241.400 1628.590 ;
        RECT 1283.500 1628.270 1283.760 1628.590 ;
        RECT 241.200 468.850 241.340 1628.270 ;
        RECT 241.140 468.530 241.400 468.850 ;
        RECT 241.140 467.510 241.400 467.830 ;
        RECT 241.200 17.410 241.340 467.510 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1629.480 1283.770 1629.760 ;
      LAYER met3 ;
        RECT 1283.465 1629.770 1283.795 1629.785 ;
        RECT 1283.465 1629.720 1300.420 1629.770 ;
        RECT 1283.465 1629.470 1304.000 1629.720 ;
        RECT 1283.465 1629.455 1283.795 1629.470 ;
        RECT 1300.000 1629.120 1304.000 1629.470 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 261.810 1656.380 262.130 1656.440 ;
        RECT 1283.470 1656.380 1283.790 1656.440 ;
        RECT 261.810 1656.240 1283.790 1656.380 ;
        RECT 261.810 1656.180 262.130 1656.240 ;
        RECT 1283.470 1656.180 1283.790 1656.240 ;
        RECT 258.130 17.920 258.450 17.980 ;
        RECT 261.810 17.920 262.130 17.980 ;
        RECT 258.130 17.780 262.130 17.920 ;
        RECT 258.130 17.720 258.450 17.780 ;
        RECT 261.810 17.720 262.130 17.780 ;
      LAYER via ;
        RECT 261.840 1656.180 262.100 1656.440 ;
        RECT 1283.500 1656.180 1283.760 1656.440 ;
        RECT 258.160 17.720 258.420 17.980 ;
        RECT 261.840 17.720 262.100 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1661.395 1283.770 1661.765 ;
        RECT 1283.560 1656.470 1283.700 1661.395 ;
        RECT 261.840 1656.150 262.100 1656.470 ;
        RECT 1283.500 1656.150 1283.760 1656.470 ;
        RECT 261.900 18.010 262.040 1656.150 ;
        RECT 258.160 17.690 258.420 18.010 ;
        RECT 261.840 17.690 262.100 18.010 ;
        RECT 258.220 2.400 258.360 17.690 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1661.440 1283.770 1661.720 ;
      LAYER met3 ;
        RECT 1283.465 1661.730 1283.795 1661.745 ;
        RECT 1283.465 1661.680 1300.420 1661.730 ;
        RECT 1283.465 1661.430 1304.000 1661.680 ;
        RECT 1283.465 1661.415 1283.795 1661.430 ;
        RECT 1300.000 1661.080 1304.000 1661.430 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 1690.720 282.370 1690.780 ;
        RECT 1283.470 1690.720 1283.790 1690.780 ;
        RECT 282.050 1690.580 1283.790 1690.720 ;
        RECT 282.050 1690.520 282.370 1690.580 ;
        RECT 1283.470 1690.520 1283.790 1690.580 ;
        RECT 276.070 17.920 276.390 17.980 ;
        RECT 282.050 17.920 282.370 17.980 ;
        RECT 276.070 17.780 282.370 17.920 ;
        RECT 276.070 17.720 276.390 17.780 ;
        RECT 282.050 17.720 282.370 17.780 ;
      LAYER via ;
        RECT 282.080 1690.520 282.340 1690.780 ;
        RECT 1283.500 1690.520 1283.760 1690.780 ;
        RECT 276.100 17.720 276.360 17.980 ;
        RECT 282.080 17.720 282.340 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1693.355 1283.770 1693.725 ;
        RECT 1283.560 1690.810 1283.700 1693.355 ;
        RECT 282.080 1690.490 282.340 1690.810 ;
        RECT 1283.500 1690.490 1283.760 1690.810 ;
        RECT 282.140 18.010 282.280 1690.490 ;
        RECT 276.100 17.690 276.360 18.010 ;
        RECT 282.080 17.690 282.340 18.010 ;
        RECT 276.160 2.400 276.300 17.690 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1693.400 1283.770 1693.680 ;
      LAYER met3 ;
        RECT 1283.465 1693.690 1283.795 1693.705 ;
        RECT 1283.465 1693.640 1300.420 1693.690 ;
        RECT 1283.465 1693.390 1304.000 1693.640 ;
        RECT 1283.465 1693.375 1283.795 1693.390 ;
        RECT 1300.000 1693.040 1304.000 1693.390 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 296.310 1725.400 296.630 1725.460 ;
        RECT 1283.470 1725.400 1283.790 1725.460 ;
        RECT 296.310 1725.260 1283.790 1725.400 ;
        RECT 296.310 1725.200 296.630 1725.260 ;
        RECT 1283.470 1725.200 1283.790 1725.260 ;
        RECT 294.010 17.920 294.330 17.980 ;
        RECT 296.310 17.920 296.630 17.980 ;
        RECT 294.010 17.780 296.630 17.920 ;
        RECT 294.010 17.720 294.330 17.780 ;
        RECT 296.310 17.720 296.630 17.780 ;
      LAYER via ;
        RECT 296.340 1725.200 296.600 1725.460 ;
        RECT 1283.500 1725.200 1283.760 1725.460 ;
        RECT 294.040 17.720 294.300 17.980 ;
        RECT 296.340 17.720 296.600 17.980 ;
      LAYER met2 ;
        RECT 296.340 1725.170 296.600 1725.490 ;
        RECT 1283.490 1725.315 1283.770 1725.685 ;
        RECT 1283.500 1725.170 1283.760 1725.315 ;
        RECT 296.400 18.010 296.540 1725.170 ;
        RECT 294.040 17.690 294.300 18.010 ;
        RECT 296.340 17.690 296.600 18.010 ;
        RECT 294.100 2.400 294.240 17.690 ;
        RECT 293.890 -4.800 294.450 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1725.360 1283.770 1725.640 ;
      LAYER met3 ;
        RECT 1283.465 1725.650 1283.795 1725.665 ;
        RECT 1283.465 1725.600 1300.420 1725.650 ;
        RECT 1283.465 1725.350 1304.000 1725.600 ;
        RECT 1283.465 1725.335 1283.795 1725.350 ;
        RECT 1300.000 1725.000 1304.000 1725.350 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 317.010 1752.940 317.330 1753.000 ;
        RECT 1283.470 1752.940 1283.790 1753.000 ;
        RECT 317.010 1752.800 1283.790 1752.940 ;
        RECT 317.010 1752.740 317.330 1752.800 ;
        RECT 1283.470 1752.740 1283.790 1752.800 ;
        RECT 311.950 15.880 312.270 15.940 ;
        RECT 317.010 15.880 317.330 15.940 ;
        RECT 311.950 15.740 317.330 15.880 ;
        RECT 311.950 15.680 312.270 15.740 ;
        RECT 317.010 15.680 317.330 15.740 ;
      LAYER via ;
        RECT 317.040 1752.740 317.300 1753.000 ;
        RECT 1283.500 1752.740 1283.760 1753.000 ;
        RECT 311.980 15.680 312.240 15.940 ;
        RECT 317.040 15.680 317.300 15.940 ;
      LAYER met2 ;
        RECT 1283.490 1757.275 1283.770 1757.645 ;
        RECT 1283.560 1753.030 1283.700 1757.275 ;
        RECT 317.040 1752.710 317.300 1753.030 ;
        RECT 1283.500 1752.710 1283.760 1753.030 ;
        RECT 317.100 15.970 317.240 1752.710 ;
        RECT 311.980 15.650 312.240 15.970 ;
        RECT 317.040 15.650 317.300 15.970 ;
        RECT 312.040 2.400 312.180 15.650 ;
        RECT 311.830 -4.800 312.390 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1757.320 1283.770 1757.600 ;
      LAYER met3 ;
        RECT 1283.465 1757.610 1283.795 1757.625 ;
        RECT 1283.465 1757.560 1300.420 1757.610 ;
        RECT 1283.465 1757.310 1304.000 1757.560 ;
        RECT 1283.465 1757.295 1283.795 1757.310 ;
        RECT 1300.000 1756.960 1304.000 1757.310 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 330.810 1787.280 331.130 1787.340 ;
        RECT 1283.470 1787.280 1283.790 1787.340 ;
        RECT 330.810 1787.140 1283.790 1787.280 ;
        RECT 330.810 1787.080 331.130 1787.140 ;
        RECT 1283.470 1787.080 1283.790 1787.140 ;
      LAYER via ;
        RECT 330.840 1787.080 331.100 1787.340 ;
        RECT 1283.500 1787.080 1283.760 1787.340 ;
      LAYER met2 ;
        RECT 1283.490 1789.235 1283.770 1789.605 ;
        RECT 1283.560 1787.370 1283.700 1789.235 ;
        RECT 330.840 1787.050 331.100 1787.370 ;
        RECT 1283.500 1787.050 1283.760 1787.370 ;
        RECT 330.900 17.410 331.040 1787.050 ;
        RECT 329.980 17.270 331.040 17.410 ;
        RECT 329.980 2.400 330.120 17.270 ;
        RECT 329.770 -4.800 330.330 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1789.280 1283.770 1789.560 ;
      LAYER met3 ;
        RECT 1283.465 1789.570 1283.795 1789.585 ;
        RECT 1283.465 1789.520 1300.420 1789.570 ;
        RECT 1283.465 1789.270 1304.000 1789.520 ;
        RECT 1283.465 1789.255 1283.795 1789.270 ;
        RECT 1300.000 1788.920 1304.000 1789.270 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 351.510 1814.820 351.830 1814.880 ;
        RECT 1283.470 1814.820 1283.790 1814.880 ;
        RECT 351.510 1814.680 1283.790 1814.820 ;
        RECT 351.510 1814.620 351.830 1814.680 ;
        RECT 1283.470 1814.620 1283.790 1814.680 ;
        RECT 347.370 17.920 347.690 17.980 ;
        RECT 351.510 17.920 351.830 17.980 ;
        RECT 347.370 17.780 351.830 17.920 ;
        RECT 347.370 17.720 347.690 17.780 ;
        RECT 351.510 17.720 351.830 17.780 ;
      LAYER via ;
        RECT 351.540 1814.620 351.800 1814.880 ;
        RECT 1283.500 1814.620 1283.760 1814.880 ;
        RECT 347.400 17.720 347.660 17.980 ;
        RECT 351.540 17.720 351.800 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1820.515 1283.770 1820.885 ;
        RECT 1283.560 1814.910 1283.700 1820.515 ;
        RECT 351.540 1814.590 351.800 1814.910 ;
        RECT 1283.500 1814.590 1283.760 1814.910 ;
        RECT 351.600 18.010 351.740 1814.590 ;
        RECT 347.400 17.690 347.660 18.010 ;
        RECT 351.540 17.690 351.800 18.010 ;
        RECT 347.460 2.400 347.600 17.690 ;
        RECT 347.250 -4.800 347.810 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1820.560 1283.770 1820.840 ;
      LAYER met3 ;
        RECT 1283.465 1820.850 1283.795 1820.865 ;
        RECT 1283.465 1820.800 1300.420 1820.850 ;
        RECT 1283.465 1820.550 1304.000 1820.800 ;
        RECT 1283.465 1820.535 1283.795 1820.550 ;
        RECT 1300.000 1820.200 1304.000 1820.550 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 1849.500 365.630 1849.560 ;
        RECT 1283.470 1849.500 1283.790 1849.560 ;
        RECT 365.310 1849.360 1283.790 1849.500 ;
        RECT 365.310 1849.300 365.630 1849.360 ;
        RECT 1283.470 1849.300 1283.790 1849.360 ;
      LAYER via ;
        RECT 365.340 1849.300 365.600 1849.560 ;
        RECT 1283.500 1849.300 1283.760 1849.560 ;
      LAYER met2 ;
        RECT 1283.490 1852.475 1283.770 1852.845 ;
        RECT 1283.560 1849.590 1283.700 1852.475 ;
        RECT 365.340 1849.270 365.600 1849.590 ;
        RECT 1283.500 1849.270 1283.760 1849.590 ;
        RECT 365.400 2.400 365.540 1849.270 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1852.520 1283.770 1852.800 ;
      LAYER met3 ;
        RECT 1283.465 1852.810 1283.795 1852.825 ;
        RECT 1283.465 1852.760 1300.420 1852.810 ;
        RECT 1283.465 1852.510 1304.000 1852.760 ;
        RECT 1283.465 1852.495 1283.795 1852.510 ;
        RECT 1300.000 1852.160 1304.000 1852.510 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 386.010 1883.840 386.330 1883.900 ;
        RECT 1283.470 1883.840 1283.790 1883.900 ;
        RECT 386.010 1883.700 1283.790 1883.840 ;
        RECT 386.010 1883.640 386.330 1883.700 ;
        RECT 1283.470 1883.640 1283.790 1883.700 ;
        RECT 383.250 17.920 383.570 17.980 ;
        RECT 386.010 17.920 386.330 17.980 ;
        RECT 383.250 17.780 386.330 17.920 ;
        RECT 383.250 17.720 383.570 17.780 ;
        RECT 386.010 17.720 386.330 17.780 ;
      LAYER via ;
        RECT 386.040 1883.640 386.300 1883.900 ;
        RECT 1283.500 1883.640 1283.760 1883.900 ;
        RECT 383.280 17.720 383.540 17.980 ;
        RECT 386.040 17.720 386.300 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1884.435 1283.770 1884.805 ;
        RECT 1283.560 1883.930 1283.700 1884.435 ;
        RECT 386.040 1883.610 386.300 1883.930 ;
        RECT 1283.500 1883.610 1283.760 1883.930 ;
        RECT 386.100 18.010 386.240 1883.610 ;
        RECT 383.280 17.690 383.540 18.010 ;
        RECT 386.040 17.690 386.300 18.010 ;
        RECT 383.340 2.400 383.480 17.690 ;
        RECT 383.130 -4.800 383.690 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1884.480 1283.770 1884.760 ;
      LAYER met3 ;
        RECT 1283.465 1884.770 1283.795 1884.785 ;
        RECT 1283.465 1884.720 1300.420 1884.770 ;
        RECT 1283.465 1884.470 1304.000 1884.720 ;
        RECT 1283.465 1884.455 1283.795 1884.470 ;
        RECT 1300.000 1884.120 1304.000 1884.470 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 406.710 1911.380 407.030 1911.440 ;
        RECT 1283.470 1911.380 1283.790 1911.440 ;
        RECT 406.710 1911.240 1283.790 1911.380 ;
        RECT 406.710 1911.180 407.030 1911.240 ;
        RECT 1283.470 1911.180 1283.790 1911.240 ;
        RECT 401.190 17.920 401.510 17.980 ;
        RECT 406.710 17.920 407.030 17.980 ;
        RECT 401.190 17.780 407.030 17.920 ;
        RECT 401.190 17.720 401.510 17.780 ;
        RECT 406.710 17.720 407.030 17.780 ;
      LAYER via ;
        RECT 406.740 1911.180 407.000 1911.440 ;
        RECT 1283.500 1911.180 1283.760 1911.440 ;
        RECT 401.220 17.720 401.480 17.980 ;
        RECT 406.740 17.720 407.000 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1916.395 1283.770 1916.765 ;
        RECT 1283.560 1911.470 1283.700 1916.395 ;
        RECT 406.740 1911.150 407.000 1911.470 ;
        RECT 1283.500 1911.150 1283.760 1911.470 ;
        RECT 406.800 18.010 406.940 1911.150 ;
        RECT 401.220 17.690 401.480 18.010 ;
        RECT 406.740 17.690 407.000 18.010 ;
        RECT 401.280 2.400 401.420 17.690 ;
        RECT 401.070 -4.800 401.630 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1916.440 1283.770 1916.720 ;
      LAYER met3 ;
        RECT 1283.465 1916.730 1283.795 1916.745 ;
        RECT 1283.465 1916.680 1300.420 1916.730 ;
        RECT 1283.465 1916.430 1304.000 1916.680 ;
        RECT 1283.465 1916.415 1283.795 1916.430 ;
        RECT 1300.000 1916.080 1304.000 1916.430 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 1311.280 68.470 1311.340 ;
        RECT 1283.470 1311.280 1283.790 1311.340 ;
        RECT 68.150 1311.140 1283.790 1311.280 ;
        RECT 68.150 1311.080 68.470 1311.140 ;
        RECT 1283.470 1311.080 1283.790 1311.140 ;
        RECT 62.170 17.920 62.490 17.980 ;
        RECT 68.150 17.920 68.470 17.980 ;
        RECT 62.170 17.780 68.470 17.920 ;
        RECT 62.170 17.720 62.490 17.780 ;
        RECT 68.150 17.720 68.470 17.780 ;
      LAYER via ;
        RECT 68.180 1311.080 68.440 1311.340 ;
        RECT 1283.500 1311.080 1283.760 1311.340 ;
        RECT 62.200 17.720 62.460 17.980 ;
        RECT 68.180 17.720 68.440 17.980 ;
      LAYER met2 ;
        RECT 68.180 1311.050 68.440 1311.370 ;
        RECT 1283.490 1311.195 1283.770 1311.565 ;
        RECT 1283.500 1311.050 1283.760 1311.195 ;
        RECT 68.240 18.010 68.380 1311.050 ;
        RECT 62.200 17.690 62.460 18.010 ;
        RECT 68.180 17.690 68.440 18.010 ;
        RECT 62.260 2.400 62.400 17.690 ;
        RECT 62.050 -4.800 62.610 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1311.240 1283.770 1311.520 ;
      LAYER met3 ;
        RECT 1283.465 1311.530 1283.795 1311.545 ;
        RECT 1283.465 1311.480 1300.420 1311.530 ;
        RECT 1283.465 1311.230 1304.000 1311.480 ;
        RECT 1283.465 1311.215 1283.795 1311.230 ;
        RECT 1300.000 1310.880 1304.000 1311.230 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 420.510 1946.060 420.830 1946.120 ;
        RECT 1283.470 1946.060 1283.790 1946.120 ;
        RECT 420.510 1945.920 1283.790 1946.060 ;
        RECT 420.510 1945.860 420.830 1945.920 ;
        RECT 1283.470 1945.860 1283.790 1945.920 ;
      LAYER via ;
        RECT 420.540 1945.860 420.800 1946.120 ;
        RECT 1283.500 1945.860 1283.760 1946.120 ;
      LAYER met2 ;
        RECT 1283.490 1948.355 1283.770 1948.725 ;
        RECT 1283.560 1946.150 1283.700 1948.355 ;
        RECT 420.540 1945.830 420.800 1946.150 ;
        RECT 1283.500 1945.830 1283.760 1946.150 ;
        RECT 420.600 17.410 420.740 1945.830 ;
        RECT 419.220 17.270 420.740 17.410 ;
        RECT 419.220 2.400 419.360 17.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1948.400 1283.770 1948.680 ;
      LAYER met3 ;
        RECT 1283.465 1948.690 1283.795 1948.705 ;
        RECT 1283.465 1948.640 1300.420 1948.690 ;
        RECT 1283.465 1948.390 1304.000 1948.640 ;
        RECT 1283.465 1948.375 1283.795 1948.390 ;
        RECT 1300.000 1948.040 1304.000 1948.390 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 441.210 1980.400 441.530 1980.460 ;
        RECT 1283.470 1980.400 1283.790 1980.460 ;
        RECT 441.210 1980.260 1283.790 1980.400 ;
        RECT 441.210 1980.200 441.530 1980.260 ;
        RECT 1283.470 1980.200 1283.790 1980.260 ;
        RECT 436.610 17.920 436.930 17.980 ;
        RECT 441.210 17.920 441.530 17.980 ;
        RECT 436.610 17.780 441.530 17.920 ;
        RECT 436.610 17.720 436.930 17.780 ;
        RECT 441.210 17.720 441.530 17.780 ;
      LAYER via ;
        RECT 441.240 1980.200 441.500 1980.460 ;
        RECT 1283.500 1980.200 1283.760 1980.460 ;
        RECT 436.640 17.720 436.900 17.980 ;
        RECT 441.240 17.720 441.500 17.980 ;
      LAYER met2 ;
        RECT 441.240 1980.170 441.500 1980.490 ;
        RECT 1283.490 1980.315 1283.770 1980.685 ;
        RECT 1283.500 1980.170 1283.760 1980.315 ;
        RECT 441.300 18.010 441.440 1980.170 ;
        RECT 436.640 17.690 436.900 18.010 ;
        RECT 441.240 17.690 441.500 18.010 ;
        RECT 436.700 2.400 436.840 17.690 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1980.360 1283.770 1980.640 ;
      LAYER met3 ;
        RECT 1283.465 1980.650 1283.795 1980.665 ;
        RECT 1283.465 1980.600 1300.420 1980.650 ;
        RECT 1283.465 1980.350 1304.000 1980.600 ;
        RECT 1283.465 1980.335 1283.795 1980.350 ;
        RECT 1300.000 1980.000 1304.000 1980.350 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 455.010 2008.280 455.330 2008.340 ;
        RECT 1283.470 2008.280 1283.790 2008.340 ;
        RECT 455.010 2008.140 1283.790 2008.280 ;
        RECT 455.010 2008.080 455.330 2008.140 ;
        RECT 1283.470 2008.080 1283.790 2008.140 ;
      LAYER via ;
        RECT 455.040 2008.080 455.300 2008.340 ;
        RECT 1283.500 2008.080 1283.760 2008.340 ;
      LAYER met2 ;
        RECT 1283.490 2012.275 1283.770 2012.645 ;
        RECT 1283.560 2008.370 1283.700 2012.275 ;
        RECT 455.040 2008.050 455.300 2008.370 ;
        RECT 1283.500 2008.050 1283.760 2008.370 ;
        RECT 455.100 17.410 455.240 2008.050 ;
        RECT 454.640 17.270 455.240 17.410 ;
        RECT 454.640 2.400 454.780 17.270 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2012.320 1283.770 2012.600 ;
      LAYER met3 ;
        RECT 1283.465 2012.610 1283.795 2012.625 ;
        RECT 1283.465 2012.560 1300.420 2012.610 ;
        RECT 1283.465 2012.310 1304.000 2012.560 ;
        RECT 1283.465 2012.295 1283.795 2012.310 ;
        RECT 1300.000 2011.960 1304.000 2012.310 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 475.710 2042.620 476.030 2042.680 ;
        RECT 1283.470 2042.620 1283.790 2042.680 ;
        RECT 475.710 2042.480 1283.790 2042.620 ;
        RECT 475.710 2042.420 476.030 2042.480 ;
        RECT 1283.470 2042.420 1283.790 2042.480 ;
        RECT 472.490 17.920 472.810 17.980 ;
        RECT 475.710 17.920 476.030 17.980 ;
        RECT 472.490 17.780 476.030 17.920 ;
        RECT 472.490 17.720 472.810 17.780 ;
        RECT 475.710 17.720 476.030 17.780 ;
      LAYER via ;
        RECT 475.740 2042.420 476.000 2042.680 ;
        RECT 1283.500 2042.420 1283.760 2042.680 ;
        RECT 472.520 17.720 472.780 17.980 ;
        RECT 475.740 17.720 476.000 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2043.555 1283.770 2043.925 ;
        RECT 1283.560 2042.710 1283.700 2043.555 ;
        RECT 475.740 2042.390 476.000 2042.710 ;
        RECT 1283.500 2042.390 1283.760 2042.710 ;
        RECT 475.800 18.010 475.940 2042.390 ;
        RECT 472.520 17.690 472.780 18.010 ;
        RECT 475.740 17.690 476.000 18.010 ;
        RECT 472.580 2.400 472.720 17.690 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2043.600 1283.770 2043.880 ;
      LAYER met3 ;
        RECT 1283.465 2043.890 1283.795 2043.905 ;
        RECT 1283.465 2043.840 1300.420 2043.890 ;
        RECT 1283.465 2043.590 1304.000 2043.840 ;
        RECT 1283.465 2043.575 1283.795 2043.590 ;
        RECT 1300.000 2043.240 1304.000 2043.590 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 2070.160 496.270 2070.220 ;
        RECT 1283.470 2070.160 1283.790 2070.220 ;
        RECT 495.950 2070.020 1283.790 2070.160 ;
        RECT 495.950 2069.960 496.270 2070.020 ;
        RECT 1283.470 2069.960 1283.790 2070.020 ;
        RECT 490.430 17.920 490.750 17.980 ;
        RECT 495.950 17.920 496.270 17.980 ;
        RECT 490.430 17.780 496.270 17.920 ;
        RECT 490.430 17.720 490.750 17.780 ;
        RECT 495.950 17.720 496.270 17.780 ;
      LAYER via ;
        RECT 495.980 2069.960 496.240 2070.220 ;
        RECT 1283.500 2069.960 1283.760 2070.220 ;
        RECT 490.460 17.720 490.720 17.980 ;
        RECT 495.980 17.720 496.240 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2075.515 1283.770 2075.885 ;
        RECT 1283.560 2070.250 1283.700 2075.515 ;
        RECT 495.980 2069.930 496.240 2070.250 ;
        RECT 1283.500 2069.930 1283.760 2070.250 ;
        RECT 496.040 18.010 496.180 2069.930 ;
        RECT 490.460 17.690 490.720 18.010 ;
        RECT 495.980 17.690 496.240 18.010 ;
        RECT 490.520 2.400 490.660 17.690 ;
        RECT 490.310 -4.800 490.870 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2075.560 1283.770 2075.840 ;
      LAYER met3 ;
        RECT 1283.465 2075.850 1283.795 2075.865 ;
        RECT 1283.465 2075.800 1300.420 2075.850 ;
        RECT 1283.465 2075.550 1304.000 2075.800 ;
        RECT 1283.465 2075.535 1283.795 2075.550 ;
        RECT 1300.000 2075.200 1304.000 2075.550 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 510.210 2104.840 510.530 2104.900 ;
        RECT 1283.470 2104.840 1283.790 2104.900 ;
        RECT 510.210 2104.700 1283.790 2104.840 ;
        RECT 510.210 2104.640 510.530 2104.700 ;
        RECT 1283.470 2104.640 1283.790 2104.700 ;
        RECT 507.910 16.560 508.230 16.620 ;
        RECT 510.210 16.560 510.530 16.620 ;
        RECT 507.910 16.420 510.530 16.560 ;
        RECT 507.910 16.360 508.230 16.420 ;
        RECT 510.210 16.360 510.530 16.420 ;
      LAYER via ;
        RECT 510.240 2104.640 510.500 2104.900 ;
        RECT 1283.500 2104.640 1283.760 2104.900 ;
        RECT 507.940 16.360 508.200 16.620 ;
        RECT 510.240 16.360 510.500 16.620 ;
      LAYER met2 ;
        RECT 1283.490 2107.475 1283.770 2107.845 ;
        RECT 1283.560 2104.930 1283.700 2107.475 ;
        RECT 510.240 2104.610 510.500 2104.930 ;
        RECT 1283.500 2104.610 1283.760 2104.930 ;
        RECT 510.300 16.650 510.440 2104.610 ;
        RECT 507.940 16.330 508.200 16.650 ;
        RECT 510.240 16.330 510.500 16.650 ;
        RECT 508.000 2.400 508.140 16.330 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2107.520 1283.770 2107.800 ;
      LAYER met3 ;
        RECT 1283.465 2107.810 1283.795 2107.825 ;
        RECT 1283.465 2107.760 1300.420 2107.810 ;
        RECT 1283.465 2107.510 1304.000 2107.760 ;
        RECT 1283.465 2107.495 1283.795 2107.510 ;
        RECT 1300.000 2107.160 1304.000 2107.510 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 530.910 2139.180 531.230 2139.240 ;
        RECT 1283.470 2139.180 1283.790 2139.240 ;
        RECT 530.910 2139.040 1283.790 2139.180 ;
        RECT 530.910 2138.980 531.230 2139.040 ;
        RECT 1283.470 2138.980 1283.790 2139.040 ;
        RECT 525.850 17.920 526.170 17.980 ;
        RECT 530.910 17.920 531.230 17.980 ;
        RECT 525.850 17.780 531.230 17.920 ;
        RECT 525.850 17.720 526.170 17.780 ;
        RECT 530.910 17.720 531.230 17.780 ;
      LAYER via ;
        RECT 530.940 2138.980 531.200 2139.240 ;
        RECT 1283.500 2138.980 1283.760 2139.240 ;
        RECT 525.880 17.720 526.140 17.980 ;
        RECT 530.940 17.720 531.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2139.435 1283.770 2139.805 ;
        RECT 1283.560 2139.270 1283.700 2139.435 ;
        RECT 530.940 2138.950 531.200 2139.270 ;
        RECT 1283.500 2138.950 1283.760 2139.270 ;
        RECT 531.000 18.010 531.140 2138.950 ;
        RECT 525.880 17.690 526.140 18.010 ;
        RECT 530.940 17.690 531.200 18.010 ;
        RECT 525.940 2.400 526.080 17.690 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2139.480 1283.770 2139.760 ;
      LAYER met3 ;
        RECT 1283.465 2139.770 1283.795 2139.785 ;
        RECT 1283.465 2139.720 1300.420 2139.770 ;
        RECT 1283.465 2139.470 1304.000 2139.720 ;
        RECT 1283.465 2139.455 1283.795 2139.470 ;
        RECT 1300.000 2139.120 1304.000 2139.470 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 544.710 2166.720 545.030 2166.780 ;
        RECT 1283.470 2166.720 1283.790 2166.780 ;
        RECT 544.710 2166.580 1283.790 2166.720 ;
        RECT 544.710 2166.520 545.030 2166.580 ;
        RECT 1283.470 2166.520 1283.790 2166.580 ;
      LAYER via ;
        RECT 544.740 2166.520 545.000 2166.780 ;
        RECT 1283.500 2166.520 1283.760 2166.780 ;
      LAYER met2 ;
        RECT 1283.490 2171.395 1283.770 2171.765 ;
        RECT 1283.560 2166.810 1283.700 2171.395 ;
        RECT 544.740 2166.490 545.000 2166.810 ;
        RECT 1283.500 2166.490 1283.760 2166.810 ;
        RECT 544.800 17.410 544.940 2166.490 ;
        RECT 543.880 17.270 544.940 17.410 ;
        RECT 543.880 2.400 544.020 17.270 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2171.440 1283.770 2171.720 ;
      LAYER met3 ;
        RECT 1283.465 2171.730 1283.795 2171.745 ;
        RECT 1283.465 2171.680 1300.420 2171.730 ;
        RECT 1283.465 2171.430 1304.000 2171.680 ;
        RECT 1283.465 2171.415 1283.795 2171.430 ;
        RECT 1300.000 2171.080 1304.000 2171.430 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 2201.400 565.730 2201.460 ;
        RECT 1283.470 2201.400 1283.790 2201.460 ;
        RECT 565.410 2201.260 1283.790 2201.400 ;
        RECT 565.410 2201.200 565.730 2201.260 ;
        RECT 1283.470 2201.200 1283.790 2201.260 ;
        RECT 561.730 17.920 562.050 17.980 ;
        RECT 565.410 17.920 565.730 17.980 ;
        RECT 561.730 17.780 565.730 17.920 ;
        RECT 561.730 17.720 562.050 17.780 ;
        RECT 565.410 17.720 565.730 17.780 ;
      LAYER via ;
        RECT 565.440 2201.200 565.700 2201.460 ;
        RECT 1283.500 2201.200 1283.760 2201.460 ;
        RECT 561.760 17.720 562.020 17.980 ;
        RECT 565.440 17.720 565.700 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2203.355 1283.770 2203.725 ;
        RECT 1283.560 2201.490 1283.700 2203.355 ;
        RECT 565.440 2201.170 565.700 2201.490 ;
        RECT 1283.500 2201.170 1283.760 2201.490 ;
        RECT 565.500 18.010 565.640 2201.170 ;
        RECT 561.760 17.690 562.020 18.010 ;
        RECT 565.440 17.690 565.700 18.010 ;
        RECT 561.820 2.400 561.960 17.690 ;
        RECT 561.610 -4.800 562.170 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2203.400 1283.770 2203.680 ;
      LAYER met3 ;
        RECT 1283.465 2203.690 1283.795 2203.705 ;
        RECT 1283.465 2203.640 1300.420 2203.690 ;
        RECT 1283.465 2203.390 1304.000 2203.640 ;
        RECT 1283.465 2203.375 1283.795 2203.390 ;
        RECT 1300.000 2203.040 1304.000 2203.390 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 2228.940 585.970 2229.000 ;
        RECT 1283.470 2228.940 1283.790 2229.000 ;
        RECT 585.650 2228.800 1283.790 2228.940 ;
        RECT 585.650 2228.740 585.970 2228.800 ;
        RECT 1283.470 2228.740 1283.790 2228.800 ;
        RECT 579.670 17.920 579.990 17.980 ;
        RECT 585.650 17.920 585.970 17.980 ;
        RECT 579.670 17.780 585.970 17.920 ;
        RECT 579.670 17.720 579.990 17.780 ;
        RECT 585.650 17.720 585.970 17.780 ;
      LAYER via ;
        RECT 585.680 2228.740 585.940 2229.000 ;
        RECT 1283.500 2228.740 1283.760 2229.000 ;
        RECT 579.700 17.720 579.960 17.980 ;
        RECT 585.680 17.720 585.940 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2235.315 1283.770 2235.685 ;
        RECT 1283.560 2229.030 1283.700 2235.315 ;
        RECT 585.680 2228.710 585.940 2229.030 ;
        RECT 1283.500 2228.710 1283.760 2229.030 ;
        RECT 585.740 18.010 585.880 2228.710 ;
        RECT 579.700 17.690 579.960 18.010 ;
        RECT 585.680 17.690 585.940 18.010 ;
        RECT 579.760 2.400 579.900 17.690 ;
        RECT 579.550 -4.800 580.110 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2235.360 1283.770 2235.640 ;
      LAYER met3 ;
        RECT 1283.465 2235.650 1283.795 2235.665 ;
        RECT 1283.465 2235.600 1300.420 2235.650 ;
        RECT 1283.465 2235.350 1304.000 2235.600 ;
        RECT 1283.465 2235.335 1283.795 2235.350 ;
        RECT 1300.000 2235.000 1304.000 2235.350 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 89.310 1352.760 89.630 1352.820 ;
        RECT 1283.470 1352.760 1283.790 1352.820 ;
        RECT 89.310 1352.620 1283.790 1352.760 ;
        RECT 89.310 1352.560 89.630 1352.620 ;
        RECT 1283.470 1352.560 1283.790 1352.620 ;
        RECT 86.090 17.920 86.410 17.980 ;
        RECT 89.310 17.920 89.630 17.980 ;
        RECT 86.090 17.780 89.630 17.920 ;
        RECT 86.090 17.720 86.410 17.780 ;
        RECT 89.310 17.720 89.630 17.780 ;
      LAYER via ;
        RECT 89.340 1352.560 89.600 1352.820 ;
        RECT 1283.500 1352.560 1283.760 1352.820 ;
        RECT 86.120 17.720 86.380 17.980 ;
        RECT 89.340 17.720 89.600 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1353.355 1283.770 1353.725 ;
        RECT 1283.560 1352.850 1283.700 1353.355 ;
        RECT 89.340 1352.530 89.600 1352.850 ;
        RECT 1283.500 1352.530 1283.760 1352.850 ;
        RECT 89.400 18.010 89.540 1352.530 ;
        RECT 86.120 17.690 86.380 18.010 ;
        RECT 89.340 17.690 89.600 18.010 ;
        RECT 86.180 2.400 86.320 17.690 ;
        RECT 85.970 -4.800 86.530 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1353.400 1283.770 1353.680 ;
      LAYER met3 ;
        RECT 1283.465 1353.690 1283.795 1353.705 ;
        RECT 1283.465 1353.640 1300.420 1353.690 ;
        RECT 1283.465 1353.390 1304.000 1353.640 ;
        RECT 1283.465 1353.375 1283.795 1353.390 ;
        RECT 1300.000 1353.040 1304.000 1353.390 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 599.910 2263.280 600.230 2263.340 ;
        RECT 1283.470 2263.280 1283.790 2263.340 ;
        RECT 599.910 2263.140 1283.790 2263.280 ;
        RECT 599.910 2263.080 600.230 2263.140 ;
        RECT 1283.470 2263.080 1283.790 2263.140 ;
        RECT 597.150 17.920 597.470 17.980 ;
        RECT 599.910 17.920 600.230 17.980 ;
        RECT 597.150 17.780 600.230 17.920 ;
        RECT 597.150 17.720 597.470 17.780 ;
        RECT 599.910 17.720 600.230 17.780 ;
      LAYER via ;
        RECT 599.940 2263.080 600.200 2263.340 ;
        RECT 1283.500 2263.080 1283.760 2263.340 ;
        RECT 597.180 17.720 597.440 17.980 ;
        RECT 599.940 17.720 600.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2266.595 1283.770 2266.965 ;
        RECT 1283.560 2263.370 1283.700 2266.595 ;
        RECT 599.940 2263.050 600.200 2263.370 ;
        RECT 1283.500 2263.050 1283.760 2263.370 ;
        RECT 600.000 18.010 600.140 2263.050 ;
        RECT 597.180 17.690 597.440 18.010 ;
        RECT 599.940 17.690 600.200 18.010 ;
        RECT 597.240 2.400 597.380 17.690 ;
        RECT 597.030 -4.800 597.590 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2266.640 1283.770 2266.920 ;
      LAYER met3 ;
        RECT 1283.465 2266.930 1283.795 2266.945 ;
        RECT 1283.465 2266.880 1300.420 2266.930 ;
        RECT 1283.465 2266.630 1304.000 2266.880 ;
        RECT 1283.465 2266.615 1283.795 2266.630 ;
        RECT 1300.000 2266.280 1304.000 2266.630 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 2297.960 620.930 2298.020 ;
        RECT 1283.470 2297.960 1283.790 2298.020 ;
        RECT 620.610 2297.820 1283.790 2297.960 ;
        RECT 620.610 2297.760 620.930 2297.820 ;
        RECT 1283.470 2297.760 1283.790 2297.820 ;
        RECT 615.090 17.920 615.410 17.980 ;
        RECT 620.610 17.920 620.930 17.980 ;
        RECT 615.090 17.780 620.930 17.920 ;
        RECT 615.090 17.720 615.410 17.780 ;
        RECT 620.610 17.720 620.930 17.780 ;
      LAYER via ;
        RECT 620.640 2297.760 620.900 2298.020 ;
        RECT 1283.500 2297.760 1283.760 2298.020 ;
        RECT 615.120 17.720 615.380 17.980 ;
        RECT 620.640 17.720 620.900 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2298.555 1283.770 2298.925 ;
        RECT 1283.560 2298.050 1283.700 2298.555 ;
        RECT 620.640 2297.730 620.900 2298.050 ;
        RECT 1283.500 2297.730 1283.760 2298.050 ;
        RECT 620.700 18.010 620.840 2297.730 ;
        RECT 615.120 17.690 615.380 18.010 ;
        RECT 620.640 17.690 620.900 18.010 ;
        RECT 615.180 2.400 615.320 17.690 ;
        RECT 614.970 -4.800 615.530 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2298.600 1283.770 2298.880 ;
      LAYER met3 ;
        RECT 1283.465 2298.890 1283.795 2298.905 ;
        RECT 1283.465 2298.840 1300.420 2298.890 ;
        RECT 1283.465 2298.590 1304.000 2298.840 ;
        RECT 1283.465 2298.575 1283.795 2298.590 ;
        RECT 1300.000 2298.240 1304.000 2298.590 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 110.010 1393.900 110.330 1393.960 ;
        RECT 1283.470 1393.900 1283.790 1393.960 ;
        RECT 110.010 1393.760 1283.790 1393.900 ;
        RECT 110.010 1393.700 110.330 1393.760 ;
        RECT 1283.470 1393.700 1283.790 1393.760 ;
      LAYER via ;
        RECT 110.040 1393.700 110.300 1393.960 ;
        RECT 1283.500 1393.700 1283.760 1393.960 ;
      LAYER met2 ;
        RECT 1283.490 1396.195 1283.770 1396.565 ;
        RECT 1283.560 1393.990 1283.700 1396.195 ;
        RECT 110.040 1393.670 110.300 1393.990 ;
        RECT 1283.500 1393.670 1283.760 1393.990 ;
        RECT 110.100 17.410 110.240 1393.670 ;
        RECT 109.640 17.270 110.240 17.410 ;
        RECT 109.640 2.400 109.780 17.270 ;
        RECT 109.430 -4.800 109.990 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1396.240 1283.770 1396.520 ;
      LAYER met3 ;
        RECT 1283.465 1396.530 1283.795 1396.545 ;
        RECT 1283.465 1396.480 1300.420 1396.530 ;
        RECT 1283.465 1396.230 1304.000 1396.480 ;
        RECT 1283.465 1396.215 1283.795 1396.230 ;
        RECT 1300.000 1395.880 1304.000 1396.230 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 137.610 1435.380 137.930 1435.440 ;
        RECT 1283.470 1435.380 1283.790 1435.440 ;
        RECT 137.610 1435.240 1283.790 1435.380 ;
        RECT 137.610 1435.180 137.930 1435.240 ;
        RECT 1283.470 1435.180 1283.790 1435.240 ;
        RECT 133.470 17.920 133.790 17.980 ;
        RECT 137.610 17.920 137.930 17.980 ;
        RECT 133.470 17.780 137.930 17.920 ;
        RECT 133.470 17.720 133.790 17.780 ;
        RECT 137.610 17.720 137.930 17.780 ;
      LAYER via ;
        RECT 137.640 1435.180 137.900 1435.440 ;
        RECT 1283.500 1435.180 1283.760 1435.440 ;
        RECT 133.500 17.720 133.760 17.980 ;
        RECT 137.640 17.720 137.900 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1438.355 1283.770 1438.725 ;
        RECT 1283.560 1435.470 1283.700 1438.355 ;
        RECT 137.640 1435.150 137.900 1435.470 ;
        RECT 1283.500 1435.150 1283.760 1435.470 ;
        RECT 137.700 18.010 137.840 1435.150 ;
        RECT 133.500 17.690 133.760 18.010 ;
        RECT 137.640 17.690 137.900 18.010 ;
        RECT 133.560 2.400 133.700 17.690 ;
        RECT 133.350 -4.800 133.910 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1438.400 1283.770 1438.680 ;
      LAYER met3 ;
        RECT 1283.465 1438.690 1283.795 1438.705 ;
        RECT 1283.465 1438.640 1300.420 1438.690 ;
        RECT 1283.465 1438.390 1304.000 1438.640 ;
        RECT 1283.465 1438.375 1283.795 1438.390 ;
        RECT 1300.000 1438.040 1304.000 1438.390 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 1470.060 151.730 1470.120 ;
        RECT 1283.470 1470.060 1283.790 1470.120 ;
        RECT 151.410 1469.920 1283.790 1470.060 ;
        RECT 151.410 1469.860 151.730 1469.920 ;
        RECT 1283.470 1469.860 1283.790 1469.920 ;
      LAYER via ;
        RECT 151.440 1469.860 151.700 1470.120 ;
        RECT 1283.500 1469.860 1283.760 1470.120 ;
      LAYER met2 ;
        RECT 1283.490 1470.315 1283.770 1470.685 ;
        RECT 1283.560 1470.150 1283.700 1470.315 ;
        RECT 151.440 1469.830 151.700 1470.150 ;
        RECT 1283.500 1469.830 1283.760 1470.150 ;
        RECT 151.500 2.400 151.640 1469.830 ;
        RECT 151.290 -4.800 151.850 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1470.360 1283.770 1470.640 ;
      LAYER met3 ;
        RECT 1283.465 1470.650 1283.795 1470.665 ;
        RECT 1283.465 1470.600 1300.420 1470.650 ;
        RECT 1283.465 1470.350 1304.000 1470.600 ;
        RECT 1283.465 1470.335 1283.795 1470.350 ;
        RECT 1300.000 1470.000 1304.000 1470.350 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 1497.600 172.430 1497.660 ;
        RECT 1283.470 1497.600 1283.790 1497.660 ;
        RECT 172.110 1497.460 1283.790 1497.600 ;
        RECT 172.110 1497.400 172.430 1497.460 ;
        RECT 1283.470 1497.400 1283.790 1497.460 ;
        RECT 169.350 17.920 169.670 17.980 ;
        RECT 172.110 17.920 172.430 17.980 ;
        RECT 169.350 17.780 172.430 17.920 ;
        RECT 169.350 17.720 169.670 17.780 ;
        RECT 172.110 17.720 172.430 17.780 ;
      LAYER via ;
        RECT 172.140 1497.400 172.400 1497.660 ;
        RECT 1283.500 1497.400 1283.760 1497.660 ;
        RECT 169.380 17.720 169.640 17.980 ;
        RECT 172.140 17.720 172.400 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1502.275 1283.770 1502.645 ;
        RECT 1283.560 1497.690 1283.700 1502.275 ;
        RECT 172.140 1497.370 172.400 1497.690 ;
        RECT 1283.500 1497.370 1283.760 1497.690 ;
        RECT 172.200 18.010 172.340 1497.370 ;
        RECT 169.380 17.690 169.640 18.010 ;
        RECT 172.140 17.690 172.400 18.010 ;
        RECT 169.440 2.400 169.580 17.690 ;
        RECT 169.230 -4.800 169.790 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1502.320 1283.770 1502.600 ;
      LAYER met3 ;
        RECT 1283.465 1502.610 1283.795 1502.625 ;
        RECT 1283.465 1502.560 1300.420 1502.610 ;
        RECT 1283.465 1502.310 1304.000 1502.560 ;
        RECT 1283.465 1502.295 1283.795 1502.310 ;
        RECT 1300.000 1501.960 1304.000 1502.310 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.350 1531.940 192.670 1532.000 ;
        RECT 1283.470 1531.940 1283.790 1532.000 ;
        RECT 192.350 1531.800 1283.790 1531.940 ;
        RECT 192.350 1531.740 192.670 1531.800 ;
        RECT 1283.470 1531.740 1283.790 1531.800 ;
        RECT 186.830 17.920 187.150 17.980 ;
        RECT 192.350 17.920 192.670 17.980 ;
        RECT 186.830 17.780 192.670 17.920 ;
        RECT 186.830 17.720 187.150 17.780 ;
        RECT 192.350 17.720 192.670 17.780 ;
      LAYER via ;
        RECT 192.380 1531.740 192.640 1532.000 ;
        RECT 1283.500 1531.740 1283.760 1532.000 ;
        RECT 186.860 17.720 187.120 17.980 ;
        RECT 192.380 17.720 192.640 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1534.235 1283.770 1534.605 ;
        RECT 1283.560 1532.030 1283.700 1534.235 ;
        RECT 192.380 1531.710 192.640 1532.030 ;
        RECT 1283.500 1531.710 1283.760 1532.030 ;
        RECT 192.440 18.010 192.580 1531.710 ;
        RECT 186.860 17.690 187.120 18.010 ;
        RECT 192.380 17.690 192.640 18.010 ;
        RECT 186.920 2.400 187.060 17.690 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1534.280 1283.770 1534.560 ;
      LAYER met3 ;
        RECT 1283.465 1534.570 1283.795 1534.585 ;
        RECT 1283.465 1534.520 1300.420 1534.570 ;
        RECT 1283.465 1534.270 1304.000 1534.520 ;
        RECT 1283.465 1534.255 1283.795 1534.270 ;
        RECT 1300.000 1533.920 1304.000 1534.270 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 206.610 1566.620 206.930 1566.680 ;
        RECT 1283.470 1566.620 1283.790 1566.680 ;
        RECT 206.610 1566.480 1283.790 1566.620 ;
        RECT 206.610 1566.420 206.930 1566.480 ;
        RECT 1283.470 1566.420 1283.790 1566.480 ;
      LAYER via ;
        RECT 206.640 1566.420 206.900 1566.680 ;
        RECT 1283.500 1566.420 1283.760 1566.680 ;
      LAYER met2 ;
        RECT 206.640 1566.390 206.900 1566.710 ;
        RECT 1283.500 1566.565 1283.760 1566.710 ;
        RECT 206.700 17.410 206.840 1566.390 ;
        RECT 1283.490 1566.195 1283.770 1566.565 ;
        RECT 204.860 17.270 206.840 17.410 ;
        RECT 204.860 2.400 205.000 17.270 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1566.240 1283.770 1566.520 ;
      LAYER met3 ;
        RECT 1283.465 1566.530 1283.795 1566.545 ;
        RECT 1283.465 1566.480 1300.420 1566.530 ;
        RECT 1283.465 1566.230 1304.000 1566.480 ;
        RECT 1283.465 1566.215 1283.795 1566.230 ;
        RECT 1300.000 1565.880 1304.000 1566.230 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 227.310 1594.160 227.630 1594.220 ;
        RECT 1283.470 1594.160 1283.790 1594.220 ;
        RECT 227.310 1594.020 1283.790 1594.160 ;
        RECT 227.310 1593.960 227.630 1594.020 ;
        RECT 1283.470 1593.960 1283.790 1594.020 ;
        RECT 222.710 17.920 223.030 17.980 ;
        RECT 227.310 17.920 227.630 17.980 ;
        RECT 222.710 17.780 227.630 17.920 ;
        RECT 222.710 17.720 223.030 17.780 ;
        RECT 227.310 17.720 227.630 17.780 ;
      LAYER via ;
        RECT 227.340 1593.960 227.600 1594.220 ;
        RECT 1283.500 1593.960 1283.760 1594.220 ;
        RECT 222.740 17.720 223.000 17.980 ;
        RECT 227.340 17.720 227.600 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1597.475 1283.770 1597.845 ;
        RECT 1283.560 1594.250 1283.700 1597.475 ;
        RECT 227.340 1593.930 227.600 1594.250 ;
        RECT 1283.500 1593.930 1283.760 1594.250 ;
        RECT 227.400 18.010 227.540 1593.930 ;
        RECT 222.740 17.690 223.000 18.010 ;
        RECT 227.340 17.690 227.600 18.010 ;
        RECT 222.800 2.400 222.940 17.690 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1597.520 1283.770 1597.800 ;
      LAYER met3 ;
        RECT 1283.465 1597.810 1283.795 1597.825 ;
        RECT 1283.465 1597.760 1300.420 1597.810 ;
        RECT 1283.465 1597.510 1304.000 1597.760 ;
        RECT 1283.465 1597.495 1283.795 1597.510 ;
        RECT 1300.000 1597.160 1304.000 1597.510 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 17.240 20.630 17.300 ;
        RECT 1286.690 17.240 1287.010 17.300 ;
        RECT 20.310 17.100 1287.010 17.240 ;
        RECT 20.310 17.040 20.630 17.100 ;
        RECT 1286.690 17.040 1287.010 17.100 ;
      LAYER via ;
        RECT 20.340 17.040 20.600 17.300 ;
        RECT 1286.720 17.040 1286.980 17.300 ;
      LAYER met2 ;
        RECT 1286.710 1236.395 1286.990 1236.765 ;
        RECT 1286.780 17.330 1286.920 1236.395 ;
        RECT 20.340 17.010 20.600 17.330 ;
        RECT 1286.720 17.010 1286.980 17.330 ;
        RECT 20.400 2.400 20.540 17.010 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 1286.710 1236.440 1286.990 1236.720 ;
      LAYER met3 ;
        RECT 1286.685 1236.730 1287.015 1236.745 ;
        RECT 1286.685 1236.680 1300.420 1236.730 ;
        RECT 1286.685 1236.430 1304.000 1236.680 ;
        RECT 1286.685 1236.415 1287.015 1236.430 ;
        RECT 1300.000 1236.080 1304.000 1236.430 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 1276.600 48.230 1276.660 ;
        RECT 1283.470 1276.600 1283.790 1276.660 ;
        RECT 47.910 1276.460 1283.790 1276.600 ;
        RECT 47.910 1276.400 48.230 1276.460 ;
        RECT 1283.470 1276.400 1283.790 1276.460 ;
        RECT 47.910 467.200 48.230 467.460 ;
        RECT 48.000 466.780 48.140 467.200 ;
        RECT 47.910 466.520 48.230 466.780 ;
        RECT 44.230 17.920 44.550 17.980 ;
        RECT 47.910 17.920 48.230 17.980 ;
        RECT 44.230 17.780 48.230 17.920 ;
        RECT 44.230 17.720 44.550 17.780 ;
        RECT 47.910 17.720 48.230 17.780 ;
      LAYER via ;
        RECT 47.940 1276.400 48.200 1276.660 ;
        RECT 1283.500 1276.400 1283.760 1276.660 ;
        RECT 47.940 467.200 48.200 467.460 ;
        RECT 47.940 466.520 48.200 466.780 ;
        RECT 44.260 17.720 44.520 17.980 ;
        RECT 47.940 17.720 48.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1279.235 1283.770 1279.605 ;
        RECT 1283.560 1276.690 1283.700 1279.235 ;
        RECT 47.940 1276.370 48.200 1276.690 ;
        RECT 1283.500 1276.370 1283.760 1276.690 ;
        RECT 48.000 467.490 48.140 1276.370 ;
        RECT 47.940 467.170 48.200 467.490 ;
        RECT 47.940 466.490 48.200 466.810 ;
        RECT 48.000 18.010 48.140 466.490 ;
        RECT 44.260 17.690 44.520 18.010 ;
        RECT 47.940 17.690 48.200 18.010 ;
        RECT 44.320 2.400 44.460 17.690 ;
        RECT 44.110 -4.800 44.670 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1279.280 1283.770 1279.560 ;
      LAYER met3 ;
        RECT 1283.465 1279.570 1283.795 1279.585 ;
        RECT 1283.465 1279.520 1300.420 1279.570 ;
        RECT 1283.465 1279.270 1304.000 1279.520 ;
        RECT 1283.465 1279.255 1283.795 1279.270 ;
        RECT 1300.000 1278.920 1304.000 1279.270 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 1635.640 248.330 1635.700 ;
        RECT 1283.470 1635.640 1283.790 1635.700 ;
        RECT 248.010 1635.500 1283.790 1635.640 ;
        RECT 248.010 1635.440 248.330 1635.500 ;
        RECT 1283.470 1635.440 1283.790 1635.500 ;
      LAYER via ;
        RECT 248.040 1635.440 248.300 1635.700 ;
        RECT 1283.500 1635.440 1283.760 1635.700 ;
      LAYER met2 ;
        RECT 1283.490 1640.315 1283.770 1640.685 ;
        RECT 1283.560 1635.730 1283.700 1640.315 ;
        RECT 248.040 1635.410 248.300 1635.730 ;
        RECT 1283.500 1635.410 1283.760 1635.730 ;
        RECT 248.100 17.410 248.240 1635.410 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1640.360 1283.770 1640.640 ;
      LAYER met3 ;
        RECT 1283.465 1640.650 1283.795 1640.665 ;
        RECT 1283.465 1640.600 1300.420 1640.650 ;
        RECT 1283.465 1640.350 1304.000 1640.600 ;
        RECT 1283.465 1640.335 1283.795 1640.350 ;
        RECT 1300.000 1640.000 1304.000 1640.350 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 1669.980 269.030 1670.040 ;
        RECT 1283.470 1669.980 1283.790 1670.040 ;
        RECT 268.710 1669.840 1283.790 1669.980 ;
        RECT 268.710 1669.780 269.030 1669.840 ;
        RECT 1283.470 1669.780 1283.790 1669.840 ;
        RECT 264.110 17.920 264.430 17.980 ;
        RECT 268.710 17.920 269.030 17.980 ;
        RECT 264.110 17.780 269.030 17.920 ;
        RECT 264.110 17.720 264.430 17.780 ;
        RECT 268.710 17.720 269.030 17.780 ;
      LAYER via ;
        RECT 268.740 1669.780 269.000 1670.040 ;
        RECT 1283.500 1669.780 1283.760 1670.040 ;
        RECT 264.140 17.720 264.400 17.980 ;
        RECT 268.740 17.720 269.000 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1672.275 1283.770 1672.645 ;
        RECT 1283.560 1670.070 1283.700 1672.275 ;
        RECT 268.740 1669.750 269.000 1670.070 ;
        RECT 1283.500 1669.750 1283.760 1670.070 ;
        RECT 268.800 18.010 268.940 1669.750 ;
        RECT 264.140 17.690 264.400 18.010 ;
        RECT 268.740 17.690 269.000 18.010 ;
        RECT 264.200 2.400 264.340 17.690 ;
        RECT 263.990 -4.800 264.550 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1672.320 1283.770 1672.600 ;
      LAYER met3 ;
        RECT 1283.465 1672.610 1283.795 1672.625 ;
        RECT 1283.465 1672.560 1300.420 1672.610 ;
        RECT 1283.465 1672.310 1304.000 1672.560 ;
        RECT 1283.465 1672.295 1283.795 1672.310 ;
        RECT 1300.000 1671.960 1304.000 1672.310 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 1704.660 282.830 1704.720 ;
        RECT 1283.470 1704.660 1283.790 1704.720 ;
        RECT 282.510 1704.520 1283.790 1704.660 ;
        RECT 282.510 1704.460 282.830 1704.520 ;
        RECT 1283.470 1704.460 1283.790 1704.520 ;
      LAYER via ;
        RECT 282.540 1704.460 282.800 1704.720 ;
        RECT 1283.500 1704.460 1283.760 1704.720 ;
      LAYER met2 ;
        RECT 282.540 1704.430 282.800 1704.750 ;
        RECT 1283.500 1704.605 1283.760 1704.750 ;
        RECT 282.600 17.410 282.740 1704.430 ;
        RECT 1283.490 1704.235 1283.770 1704.605 ;
        RECT 282.140 17.270 282.740 17.410 ;
        RECT 282.140 2.400 282.280 17.270 ;
        RECT 281.930 -4.800 282.490 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1704.280 1283.770 1704.560 ;
      LAYER met3 ;
        RECT 1283.465 1704.570 1283.795 1704.585 ;
        RECT 1283.465 1704.520 1300.420 1704.570 ;
        RECT 1283.465 1704.270 1304.000 1704.520 ;
        RECT 1283.465 1704.255 1283.795 1704.270 ;
        RECT 1300.000 1703.920 1304.000 1704.270 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 1732.200 303.530 1732.260 ;
        RECT 1283.470 1732.200 1283.790 1732.260 ;
        RECT 303.210 1732.060 1283.790 1732.200 ;
        RECT 303.210 1732.000 303.530 1732.060 ;
        RECT 1283.470 1732.000 1283.790 1732.060 ;
        RECT 299.990 17.920 300.310 17.980 ;
        RECT 303.210 17.920 303.530 17.980 ;
        RECT 299.990 17.780 303.530 17.920 ;
        RECT 299.990 17.720 300.310 17.780 ;
        RECT 303.210 17.720 303.530 17.780 ;
      LAYER via ;
        RECT 303.240 1732.000 303.500 1732.260 ;
        RECT 1283.500 1732.000 1283.760 1732.260 ;
        RECT 300.020 17.720 300.280 17.980 ;
        RECT 303.240 17.720 303.500 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1735.515 1283.770 1735.885 ;
        RECT 1283.560 1732.290 1283.700 1735.515 ;
        RECT 303.240 1731.970 303.500 1732.290 ;
        RECT 1283.500 1731.970 1283.760 1732.290 ;
        RECT 303.300 18.010 303.440 1731.970 ;
        RECT 300.020 17.690 300.280 18.010 ;
        RECT 303.240 17.690 303.500 18.010 ;
        RECT 300.080 2.400 300.220 17.690 ;
        RECT 299.870 -4.800 300.430 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1735.560 1283.770 1735.840 ;
      LAYER met3 ;
        RECT 1283.465 1735.850 1283.795 1735.865 ;
        RECT 1283.465 1735.800 1300.420 1735.850 ;
        RECT 1283.465 1735.550 1304.000 1735.800 ;
        RECT 1283.465 1735.535 1283.795 1735.550 ;
        RECT 1300.000 1735.200 1304.000 1735.550 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.450 1766.540 323.770 1766.600 ;
        RECT 1283.470 1766.540 1283.790 1766.600 ;
        RECT 323.450 1766.400 1283.790 1766.540 ;
        RECT 323.450 1766.340 323.770 1766.400 ;
        RECT 1283.470 1766.340 1283.790 1766.400 ;
        RECT 317.930 17.920 318.250 17.980 ;
        RECT 323.450 17.920 323.770 17.980 ;
        RECT 317.930 17.780 323.770 17.920 ;
        RECT 317.930 17.720 318.250 17.780 ;
        RECT 323.450 17.720 323.770 17.780 ;
      LAYER via ;
        RECT 323.480 1766.340 323.740 1766.600 ;
        RECT 1283.500 1766.340 1283.760 1766.600 ;
        RECT 317.960 17.720 318.220 17.980 ;
        RECT 323.480 17.720 323.740 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1767.475 1283.770 1767.845 ;
        RECT 1283.560 1766.630 1283.700 1767.475 ;
        RECT 323.480 1766.310 323.740 1766.630 ;
        RECT 1283.500 1766.310 1283.760 1766.630 ;
        RECT 323.540 18.010 323.680 1766.310 ;
        RECT 317.960 17.690 318.220 18.010 ;
        RECT 323.480 17.690 323.740 18.010 ;
        RECT 318.020 2.400 318.160 17.690 ;
        RECT 317.810 -4.800 318.370 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1767.520 1283.770 1767.800 ;
      LAYER met3 ;
        RECT 1283.465 1767.810 1283.795 1767.825 ;
        RECT 1283.465 1767.760 1300.420 1767.810 ;
        RECT 1283.465 1767.510 1304.000 1767.760 ;
        RECT 1283.465 1767.495 1283.795 1767.510 ;
        RECT 1300.000 1767.160 1304.000 1767.510 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 337.710 1794.080 338.030 1794.140 ;
        RECT 1283.470 1794.080 1283.790 1794.140 ;
        RECT 337.710 1793.940 1283.790 1794.080 ;
        RECT 337.710 1793.880 338.030 1793.940 ;
        RECT 1283.470 1793.880 1283.790 1793.940 ;
      LAYER via ;
        RECT 337.740 1793.880 338.000 1794.140 ;
        RECT 1283.500 1793.880 1283.760 1794.140 ;
      LAYER met2 ;
        RECT 1283.490 1799.435 1283.770 1799.805 ;
        RECT 1283.560 1794.170 1283.700 1799.435 ;
        RECT 337.740 1793.850 338.000 1794.170 ;
        RECT 1283.500 1793.850 1283.760 1794.170 ;
        RECT 337.800 17.410 337.940 1793.850 ;
        RECT 335.960 17.270 337.940 17.410 ;
        RECT 335.960 2.400 336.100 17.270 ;
        RECT 335.750 -4.800 336.310 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1799.480 1283.770 1799.760 ;
      LAYER met3 ;
        RECT 1283.465 1799.770 1283.795 1799.785 ;
        RECT 1283.465 1799.720 1300.420 1799.770 ;
        RECT 1283.465 1799.470 1304.000 1799.720 ;
        RECT 1283.465 1799.455 1283.795 1799.470 ;
        RECT 1300.000 1799.120 1304.000 1799.470 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 1828.760 358.730 1828.820 ;
        RECT 1283.470 1828.760 1283.790 1828.820 ;
        RECT 358.410 1828.620 1283.790 1828.760 ;
        RECT 358.410 1828.560 358.730 1828.620 ;
        RECT 1283.470 1828.560 1283.790 1828.620 ;
        RECT 353.350 17.920 353.670 17.980 ;
        RECT 358.410 17.920 358.730 17.980 ;
        RECT 353.350 17.780 358.730 17.920 ;
        RECT 353.350 17.720 353.670 17.780 ;
        RECT 358.410 17.720 358.730 17.780 ;
      LAYER via ;
        RECT 358.440 1828.560 358.700 1828.820 ;
        RECT 1283.500 1828.560 1283.760 1828.820 ;
        RECT 353.380 17.720 353.640 17.980 ;
        RECT 358.440 17.720 358.700 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1831.395 1283.770 1831.765 ;
        RECT 1283.560 1828.850 1283.700 1831.395 ;
        RECT 358.440 1828.530 358.700 1828.850 ;
        RECT 1283.500 1828.530 1283.760 1828.850 ;
        RECT 358.500 18.010 358.640 1828.530 ;
        RECT 353.380 17.690 353.640 18.010 ;
        RECT 358.440 17.690 358.700 18.010 ;
        RECT 353.440 2.400 353.580 17.690 ;
        RECT 353.230 -4.800 353.790 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1831.440 1283.770 1831.720 ;
      LAYER met3 ;
        RECT 1283.465 1831.730 1283.795 1831.745 ;
        RECT 1283.465 1831.680 1300.420 1831.730 ;
        RECT 1283.465 1831.430 1304.000 1831.680 ;
        RECT 1283.465 1831.415 1283.795 1831.430 ;
        RECT 1300.000 1831.080 1304.000 1831.430 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 372.210 1863.100 372.530 1863.160 ;
        RECT 1283.470 1863.100 1283.790 1863.160 ;
        RECT 372.210 1862.960 1283.790 1863.100 ;
        RECT 372.210 1862.900 372.530 1862.960 ;
        RECT 1283.470 1862.900 1283.790 1862.960 ;
      LAYER via ;
        RECT 372.240 1862.900 372.500 1863.160 ;
        RECT 1283.500 1862.900 1283.760 1863.160 ;
      LAYER met2 ;
        RECT 1283.490 1863.355 1283.770 1863.725 ;
        RECT 1283.560 1863.190 1283.700 1863.355 ;
        RECT 372.240 1862.870 372.500 1863.190 ;
        RECT 1283.500 1862.870 1283.760 1863.190 ;
        RECT 372.300 17.410 372.440 1862.870 ;
        RECT 371.380 17.270 372.440 17.410 ;
        RECT 371.380 2.400 371.520 17.270 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1863.400 1283.770 1863.680 ;
      LAYER met3 ;
        RECT 1283.465 1863.690 1283.795 1863.705 ;
        RECT 1283.465 1863.640 1300.420 1863.690 ;
        RECT 1283.465 1863.390 1304.000 1863.640 ;
        RECT 1283.465 1863.375 1283.795 1863.390 ;
        RECT 1300.000 1863.040 1304.000 1863.390 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 1890.980 393.230 1891.040 ;
        RECT 1283.470 1890.980 1283.790 1891.040 ;
        RECT 392.910 1890.840 1283.790 1890.980 ;
        RECT 392.910 1890.780 393.230 1890.840 ;
        RECT 1283.470 1890.780 1283.790 1890.840 ;
        RECT 389.230 17.920 389.550 17.980 ;
        RECT 392.910 17.920 393.230 17.980 ;
        RECT 389.230 17.780 393.230 17.920 ;
        RECT 389.230 17.720 389.550 17.780 ;
        RECT 392.910 17.720 393.230 17.780 ;
      LAYER via ;
        RECT 392.940 1890.780 393.200 1891.040 ;
        RECT 1283.500 1890.780 1283.760 1891.040 ;
        RECT 389.260 17.720 389.520 17.980 ;
        RECT 392.940 17.720 393.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1895.315 1283.770 1895.685 ;
        RECT 1283.560 1891.070 1283.700 1895.315 ;
        RECT 392.940 1890.750 393.200 1891.070 ;
        RECT 1283.500 1890.750 1283.760 1891.070 ;
        RECT 393.000 18.010 393.140 1890.750 ;
        RECT 389.260 17.690 389.520 18.010 ;
        RECT 392.940 17.690 393.200 18.010 ;
        RECT 389.320 2.400 389.460 17.690 ;
        RECT 389.110 -4.800 389.670 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1895.360 1283.770 1895.640 ;
      LAYER met3 ;
        RECT 1283.465 1895.650 1283.795 1895.665 ;
        RECT 1283.465 1895.600 1300.420 1895.650 ;
        RECT 1283.465 1895.350 1304.000 1895.600 ;
        RECT 1283.465 1895.335 1283.795 1895.350 ;
        RECT 1300.000 1895.000 1304.000 1895.350 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.150 1925.320 413.470 1925.380 ;
        RECT 1283.470 1925.320 1283.790 1925.380 ;
        RECT 413.150 1925.180 1283.790 1925.320 ;
        RECT 413.150 1925.120 413.470 1925.180 ;
        RECT 1283.470 1925.120 1283.790 1925.180 ;
        RECT 407.170 17.920 407.490 17.980 ;
        RECT 413.150 17.920 413.470 17.980 ;
        RECT 407.170 17.780 413.470 17.920 ;
        RECT 407.170 17.720 407.490 17.780 ;
        RECT 413.150 17.720 413.470 17.780 ;
      LAYER via ;
        RECT 413.180 1925.120 413.440 1925.380 ;
        RECT 1283.500 1925.120 1283.760 1925.380 ;
        RECT 407.200 17.720 407.460 17.980 ;
        RECT 413.180 17.720 413.440 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1927.275 1283.770 1927.645 ;
        RECT 1283.560 1925.410 1283.700 1927.275 ;
        RECT 413.180 1925.090 413.440 1925.410 ;
        RECT 1283.500 1925.090 1283.760 1925.410 ;
        RECT 413.240 18.010 413.380 1925.090 ;
        RECT 407.200 17.690 407.460 18.010 ;
        RECT 413.180 17.690 413.440 18.010 ;
        RECT 407.260 2.400 407.400 17.690 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1927.320 1283.770 1927.600 ;
      LAYER met3 ;
        RECT 1283.465 1927.610 1283.795 1927.625 ;
        RECT 1283.465 1927.560 1300.420 1927.610 ;
        RECT 1283.465 1927.310 1304.000 1927.560 ;
        RECT 1283.465 1927.295 1283.795 1927.310 ;
        RECT 1300.000 1926.960 1304.000 1927.310 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.610 1318.080 68.930 1318.140 ;
        RECT 1283.470 1318.080 1283.790 1318.140 ;
        RECT 68.610 1317.940 1283.790 1318.080 ;
        RECT 68.610 1317.880 68.930 1317.940 ;
        RECT 1283.470 1317.880 1283.790 1317.940 ;
      LAYER via ;
        RECT 68.640 1317.880 68.900 1318.140 ;
        RECT 1283.500 1317.880 1283.760 1318.140 ;
      LAYER met2 ;
        RECT 1283.490 1321.395 1283.770 1321.765 ;
        RECT 1283.560 1318.170 1283.700 1321.395 ;
        RECT 68.640 1317.850 68.900 1318.170 ;
        RECT 1283.500 1317.850 1283.760 1318.170 ;
        RECT 68.700 17.410 68.840 1317.850 ;
        RECT 68.240 17.270 68.840 17.410 ;
        RECT 68.240 2.400 68.380 17.270 ;
        RECT 68.030 -4.800 68.590 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1321.440 1283.770 1321.720 ;
      LAYER met3 ;
        RECT 1283.465 1321.730 1283.795 1321.745 ;
        RECT 1283.465 1321.680 1300.420 1321.730 ;
        RECT 1283.465 1321.430 1304.000 1321.680 ;
        RECT 1283.465 1321.415 1283.795 1321.430 ;
        RECT 1300.000 1321.080 1304.000 1321.430 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 1952.860 427.730 1952.920 ;
        RECT 1283.470 1952.860 1283.790 1952.920 ;
        RECT 427.410 1952.720 1283.790 1952.860 ;
        RECT 427.410 1952.660 427.730 1952.720 ;
        RECT 1283.470 1952.660 1283.790 1952.720 ;
        RECT 424.650 17.920 424.970 17.980 ;
        RECT 427.410 17.920 427.730 17.980 ;
        RECT 424.650 17.780 427.730 17.920 ;
        RECT 424.650 17.720 424.970 17.780 ;
        RECT 427.410 17.720 427.730 17.780 ;
      LAYER via ;
        RECT 427.440 1952.660 427.700 1952.920 ;
        RECT 1283.500 1952.660 1283.760 1952.920 ;
        RECT 424.680 17.720 424.940 17.980 ;
        RECT 427.440 17.720 427.700 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1958.555 1283.770 1958.925 ;
        RECT 1283.560 1952.950 1283.700 1958.555 ;
        RECT 427.440 1952.630 427.700 1952.950 ;
        RECT 1283.500 1952.630 1283.760 1952.950 ;
        RECT 427.500 18.010 427.640 1952.630 ;
        RECT 424.680 17.690 424.940 18.010 ;
        RECT 427.440 17.690 427.700 18.010 ;
        RECT 424.740 2.400 424.880 17.690 ;
        RECT 424.530 -4.800 425.090 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1958.600 1283.770 1958.880 ;
      LAYER met3 ;
        RECT 1283.465 1958.890 1283.795 1958.905 ;
        RECT 1283.465 1958.840 1300.420 1958.890 ;
        RECT 1283.465 1958.590 1304.000 1958.840 ;
        RECT 1283.465 1958.575 1283.795 1958.590 ;
        RECT 1300.000 1958.240 1304.000 1958.590 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 448.110 1987.540 448.430 1987.600 ;
        RECT 1283.470 1987.540 1283.790 1987.600 ;
        RECT 448.110 1987.400 1283.790 1987.540 ;
        RECT 448.110 1987.340 448.430 1987.400 ;
        RECT 1283.470 1987.340 1283.790 1987.400 ;
        RECT 442.590 17.920 442.910 17.980 ;
        RECT 448.110 17.920 448.430 17.980 ;
        RECT 442.590 17.780 448.430 17.920 ;
        RECT 442.590 17.720 442.910 17.780 ;
        RECT 448.110 17.720 448.430 17.780 ;
      LAYER via ;
        RECT 448.140 1987.340 448.400 1987.600 ;
        RECT 1283.500 1987.340 1283.760 1987.600 ;
        RECT 442.620 17.720 442.880 17.980 ;
        RECT 448.140 17.720 448.400 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1990.515 1283.770 1990.885 ;
        RECT 1283.560 1987.630 1283.700 1990.515 ;
        RECT 448.140 1987.310 448.400 1987.630 ;
        RECT 1283.500 1987.310 1283.760 1987.630 ;
        RECT 448.200 18.010 448.340 1987.310 ;
        RECT 442.620 17.690 442.880 18.010 ;
        RECT 448.140 17.690 448.400 18.010 ;
        RECT 442.680 2.400 442.820 17.690 ;
        RECT 442.470 -4.800 443.030 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1990.560 1283.770 1990.840 ;
      LAYER met3 ;
        RECT 1283.465 1990.850 1283.795 1990.865 ;
        RECT 1283.465 1990.800 1300.420 1990.850 ;
        RECT 1283.465 1990.550 1304.000 1990.800 ;
        RECT 1283.465 1990.535 1283.795 1990.550 ;
        RECT 1300.000 1990.200 1304.000 1990.550 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 461.910 2021.880 462.230 2021.940 ;
        RECT 1283.470 2021.880 1283.790 2021.940 ;
        RECT 461.910 2021.740 1283.790 2021.880 ;
        RECT 461.910 2021.680 462.230 2021.740 ;
        RECT 1283.470 2021.680 1283.790 2021.740 ;
      LAYER via ;
        RECT 461.940 2021.680 462.200 2021.940 ;
        RECT 1283.500 2021.680 1283.760 2021.940 ;
      LAYER met2 ;
        RECT 1283.490 2022.475 1283.770 2022.845 ;
        RECT 1283.560 2021.970 1283.700 2022.475 ;
        RECT 461.940 2021.650 462.200 2021.970 ;
        RECT 1283.500 2021.650 1283.760 2021.970 ;
        RECT 462.000 17.410 462.140 2021.650 ;
        RECT 460.620 17.270 462.140 17.410 ;
        RECT 460.620 2.400 460.760 17.270 ;
        RECT 460.410 -4.800 460.970 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2022.520 1283.770 2022.800 ;
      LAYER met3 ;
        RECT 1283.465 2022.810 1283.795 2022.825 ;
        RECT 1283.465 2022.760 1300.420 2022.810 ;
        RECT 1283.465 2022.510 1304.000 2022.760 ;
        RECT 1283.465 2022.495 1283.795 2022.510 ;
        RECT 1300.000 2022.160 1304.000 2022.510 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 2049.420 482.930 2049.480 ;
        RECT 1283.470 2049.420 1283.790 2049.480 ;
        RECT 482.610 2049.280 1283.790 2049.420 ;
        RECT 482.610 2049.220 482.930 2049.280 ;
        RECT 1283.470 2049.220 1283.790 2049.280 ;
        RECT 478.470 17.920 478.790 17.980 ;
        RECT 482.610 17.920 482.930 17.980 ;
        RECT 478.470 17.780 482.930 17.920 ;
        RECT 478.470 17.720 478.790 17.780 ;
        RECT 482.610 17.720 482.930 17.780 ;
      LAYER via ;
        RECT 482.640 2049.220 482.900 2049.480 ;
        RECT 1283.500 2049.220 1283.760 2049.480 ;
        RECT 478.500 17.720 478.760 17.980 ;
        RECT 482.640 17.720 482.900 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2054.435 1283.770 2054.805 ;
        RECT 1283.560 2049.510 1283.700 2054.435 ;
        RECT 482.640 2049.190 482.900 2049.510 ;
        RECT 1283.500 2049.190 1283.760 2049.510 ;
        RECT 482.700 18.010 482.840 2049.190 ;
        RECT 478.500 17.690 478.760 18.010 ;
        RECT 482.640 17.690 482.900 18.010 ;
        RECT 478.560 2.400 478.700 17.690 ;
        RECT 478.350 -4.800 478.910 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2054.480 1283.770 2054.760 ;
      LAYER met3 ;
        RECT 1283.465 2054.770 1283.795 2054.785 ;
        RECT 1283.465 2054.720 1300.420 2054.770 ;
        RECT 1283.465 2054.470 1304.000 2054.720 ;
        RECT 1283.465 2054.455 1283.795 2054.470 ;
        RECT 1300.000 2054.120 1304.000 2054.470 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 2084.100 496.730 2084.160 ;
        RECT 1283.470 2084.100 1283.790 2084.160 ;
        RECT 496.410 2083.960 1283.790 2084.100 ;
        RECT 496.410 2083.900 496.730 2083.960 ;
        RECT 1283.470 2083.900 1283.790 2083.960 ;
      LAYER via ;
        RECT 496.440 2083.900 496.700 2084.160 ;
        RECT 1283.500 2083.900 1283.760 2084.160 ;
      LAYER met2 ;
        RECT 1283.490 2086.395 1283.770 2086.765 ;
        RECT 1283.560 2084.190 1283.700 2086.395 ;
        RECT 496.440 2083.870 496.700 2084.190 ;
        RECT 1283.500 2083.870 1283.760 2084.190 ;
        RECT 496.500 2.400 496.640 2083.870 ;
        RECT 496.290 -4.800 496.850 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2086.440 1283.770 2086.720 ;
      LAYER met3 ;
        RECT 1283.465 2086.730 1283.795 2086.745 ;
        RECT 1283.465 2086.680 1300.420 2086.730 ;
        RECT 1283.465 2086.430 1304.000 2086.680 ;
        RECT 1283.465 2086.415 1283.795 2086.430 ;
        RECT 1300.000 2086.080 1304.000 2086.430 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 2118.440 517.430 2118.500 ;
        RECT 1283.470 2118.440 1283.790 2118.500 ;
        RECT 517.110 2118.300 1283.790 2118.440 ;
        RECT 517.110 2118.240 517.430 2118.300 ;
        RECT 1283.470 2118.240 1283.790 2118.300 ;
        RECT 513.890 17.920 514.210 17.980 ;
        RECT 517.110 17.920 517.430 17.980 ;
        RECT 513.890 17.780 517.430 17.920 ;
        RECT 513.890 17.720 514.210 17.780 ;
        RECT 517.110 17.720 517.430 17.780 ;
      LAYER via ;
        RECT 517.140 2118.240 517.400 2118.500 ;
        RECT 1283.500 2118.240 1283.760 2118.500 ;
        RECT 513.920 17.720 514.180 17.980 ;
        RECT 517.140 17.720 517.400 17.980 ;
      LAYER met2 ;
        RECT 517.140 2118.210 517.400 2118.530 ;
        RECT 1283.490 2118.355 1283.770 2118.725 ;
        RECT 1283.500 2118.210 1283.760 2118.355 ;
        RECT 517.200 18.010 517.340 2118.210 ;
        RECT 513.920 17.690 514.180 18.010 ;
        RECT 517.140 17.690 517.400 18.010 ;
        RECT 513.980 2.400 514.120 17.690 ;
        RECT 513.770 -4.800 514.330 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2118.400 1283.770 2118.680 ;
      LAYER met3 ;
        RECT 1283.465 2118.690 1283.795 2118.705 ;
        RECT 1283.465 2118.640 1300.420 2118.690 ;
        RECT 1283.465 2118.390 1304.000 2118.640 ;
        RECT 1283.465 2118.375 1283.795 2118.390 ;
        RECT 1300.000 2118.040 1304.000 2118.390 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 2145.980 537.670 2146.040 ;
        RECT 1283.470 2145.980 1283.790 2146.040 ;
        RECT 537.350 2145.840 1283.790 2145.980 ;
        RECT 537.350 2145.780 537.670 2145.840 ;
        RECT 1283.470 2145.780 1283.790 2145.840 ;
        RECT 531.830 17.920 532.150 17.980 ;
        RECT 537.350 17.920 537.670 17.980 ;
        RECT 531.830 17.780 537.670 17.920 ;
        RECT 531.830 17.720 532.150 17.780 ;
        RECT 537.350 17.720 537.670 17.780 ;
      LAYER via ;
        RECT 537.380 2145.780 537.640 2146.040 ;
        RECT 1283.500 2145.780 1283.760 2146.040 ;
        RECT 531.860 17.720 532.120 17.980 ;
        RECT 537.380 17.720 537.640 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2150.315 1283.770 2150.685 ;
        RECT 1283.560 2146.070 1283.700 2150.315 ;
        RECT 537.380 2145.750 537.640 2146.070 ;
        RECT 1283.500 2145.750 1283.760 2146.070 ;
        RECT 537.440 18.010 537.580 2145.750 ;
        RECT 531.860 17.690 532.120 18.010 ;
        RECT 537.380 17.690 537.640 18.010 ;
        RECT 531.920 2.400 532.060 17.690 ;
        RECT 531.710 -4.800 532.270 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2150.360 1283.770 2150.640 ;
      LAYER met3 ;
        RECT 1283.465 2150.650 1283.795 2150.665 ;
        RECT 1283.465 2150.600 1300.420 2150.650 ;
        RECT 1283.465 2150.350 1304.000 2150.600 ;
        RECT 1283.465 2150.335 1283.795 2150.350 ;
        RECT 1300.000 2150.000 1304.000 2150.350 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 2180.660 551.930 2180.720 ;
        RECT 1283.470 2180.660 1283.790 2180.720 ;
        RECT 551.610 2180.520 1283.790 2180.660 ;
        RECT 551.610 2180.460 551.930 2180.520 ;
        RECT 1283.470 2180.460 1283.790 2180.520 ;
      LAYER via ;
        RECT 551.640 2180.460 551.900 2180.720 ;
        RECT 1283.500 2180.460 1283.760 2180.720 ;
      LAYER met2 ;
        RECT 1283.490 2181.595 1283.770 2181.965 ;
        RECT 1283.560 2180.750 1283.700 2181.595 ;
        RECT 551.640 2180.430 551.900 2180.750 ;
        RECT 1283.500 2180.430 1283.760 2180.750 ;
        RECT 551.700 17.410 551.840 2180.430 ;
        RECT 549.860 17.270 551.840 17.410 ;
        RECT 549.860 2.400 550.000 17.270 ;
        RECT 549.650 -4.800 550.210 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2181.640 1283.770 2181.920 ;
      LAYER met3 ;
        RECT 1283.465 2181.930 1283.795 2181.945 ;
        RECT 1283.465 2181.880 1300.420 2181.930 ;
        RECT 1283.465 2181.630 1304.000 2181.880 ;
        RECT 1283.465 2181.615 1283.795 2181.630 ;
        RECT 1300.000 2181.280 1304.000 2181.630 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 2208.200 572.630 2208.260 ;
        RECT 1283.470 2208.200 1283.790 2208.260 ;
        RECT 572.310 2208.060 1283.790 2208.200 ;
        RECT 572.310 2208.000 572.630 2208.060 ;
        RECT 1283.470 2208.000 1283.790 2208.060 ;
        RECT 567.710 17.920 568.030 17.980 ;
        RECT 572.310 17.920 572.630 17.980 ;
        RECT 567.710 17.780 572.630 17.920 ;
        RECT 567.710 17.720 568.030 17.780 ;
        RECT 572.310 17.720 572.630 17.780 ;
      LAYER via ;
        RECT 572.340 2208.000 572.600 2208.260 ;
        RECT 1283.500 2208.000 1283.760 2208.260 ;
        RECT 567.740 17.720 568.000 17.980 ;
        RECT 572.340 17.720 572.600 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2213.555 1283.770 2213.925 ;
        RECT 1283.560 2208.290 1283.700 2213.555 ;
        RECT 572.340 2207.970 572.600 2208.290 ;
        RECT 1283.500 2207.970 1283.760 2208.290 ;
        RECT 572.400 18.010 572.540 2207.970 ;
        RECT 567.740 17.690 568.000 18.010 ;
        RECT 572.340 17.690 572.600 18.010 ;
        RECT 567.800 2.400 567.940 17.690 ;
        RECT 567.590 -4.800 568.150 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2213.600 1283.770 2213.880 ;
      LAYER met3 ;
        RECT 1283.465 2213.890 1283.795 2213.905 ;
        RECT 1283.465 2213.840 1300.420 2213.890 ;
        RECT 1283.465 2213.590 1304.000 2213.840 ;
        RECT 1283.465 2213.575 1283.795 2213.590 ;
        RECT 1300.000 2213.240 1304.000 2213.590 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 2242.880 586.430 2242.940 ;
        RECT 1283.470 2242.880 1283.790 2242.940 ;
        RECT 586.110 2242.740 1283.790 2242.880 ;
        RECT 586.110 2242.680 586.430 2242.740 ;
        RECT 1283.470 2242.680 1283.790 2242.740 ;
      LAYER via ;
        RECT 586.140 2242.680 586.400 2242.940 ;
        RECT 1283.500 2242.680 1283.760 2242.940 ;
      LAYER met2 ;
        RECT 1283.490 2245.515 1283.770 2245.885 ;
        RECT 1283.560 2242.970 1283.700 2245.515 ;
        RECT 586.140 2242.650 586.400 2242.970 ;
        RECT 1283.500 2242.650 1283.760 2242.970 ;
        RECT 586.200 17.410 586.340 2242.650 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2245.560 1283.770 2245.840 ;
      LAYER met3 ;
        RECT 1283.465 2245.850 1283.795 2245.865 ;
        RECT 1283.465 2245.800 1300.420 2245.850 ;
        RECT 1283.465 2245.550 1304.000 2245.800 ;
        RECT 1283.465 2245.535 1283.795 2245.550 ;
        RECT 1300.000 2245.200 1304.000 2245.550 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 96.210 1359.560 96.530 1359.620 ;
        RECT 1283.470 1359.560 1283.790 1359.620 ;
        RECT 96.210 1359.420 1283.790 1359.560 ;
        RECT 96.210 1359.360 96.530 1359.420 ;
        RECT 1283.470 1359.360 1283.790 1359.420 ;
        RECT 91.610 17.920 91.930 17.980 ;
        RECT 96.210 17.920 96.530 17.980 ;
        RECT 91.610 17.780 96.530 17.920 ;
        RECT 91.610 17.720 91.930 17.780 ;
        RECT 96.210 17.720 96.530 17.780 ;
      LAYER via ;
        RECT 96.240 1359.360 96.500 1359.620 ;
        RECT 1283.500 1359.360 1283.760 1359.620 ;
        RECT 91.640 17.720 91.900 17.980 ;
        RECT 96.240 17.720 96.500 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1364.235 1283.770 1364.605 ;
        RECT 1283.560 1359.650 1283.700 1364.235 ;
        RECT 96.240 1359.330 96.500 1359.650 ;
        RECT 1283.500 1359.330 1283.760 1359.650 ;
        RECT 96.300 18.010 96.440 1359.330 ;
        RECT 91.640 17.690 91.900 18.010 ;
        RECT 96.240 17.690 96.500 18.010 ;
        RECT 91.700 2.400 91.840 17.690 ;
        RECT 91.490 -4.800 92.050 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1364.280 1283.770 1364.560 ;
      LAYER met3 ;
        RECT 1283.465 1364.570 1283.795 1364.585 ;
        RECT 1283.465 1364.520 1300.420 1364.570 ;
        RECT 1283.465 1364.270 1304.000 1364.520 ;
        RECT 1283.465 1364.255 1283.795 1364.270 ;
        RECT 1300.000 1363.920 1304.000 1364.270 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 2277.220 607.130 2277.280 ;
        RECT 1283.470 2277.220 1283.790 2277.280 ;
        RECT 606.810 2277.080 1283.790 2277.220 ;
        RECT 606.810 2277.020 607.130 2277.080 ;
        RECT 1283.470 2277.020 1283.790 2277.080 ;
        RECT 603.130 17.920 603.450 17.980 ;
        RECT 606.810 17.920 607.130 17.980 ;
        RECT 603.130 17.780 607.130 17.920 ;
        RECT 603.130 17.720 603.450 17.780 ;
        RECT 606.810 17.720 607.130 17.780 ;
      LAYER via ;
        RECT 606.840 2277.020 607.100 2277.280 ;
        RECT 1283.500 2277.020 1283.760 2277.280 ;
        RECT 603.160 17.720 603.420 17.980 ;
        RECT 606.840 17.720 607.100 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2277.475 1283.770 2277.845 ;
        RECT 1283.560 2277.310 1283.700 2277.475 ;
        RECT 606.840 2276.990 607.100 2277.310 ;
        RECT 1283.500 2276.990 1283.760 2277.310 ;
        RECT 606.900 18.010 607.040 2276.990 ;
        RECT 603.160 17.690 603.420 18.010 ;
        RECT 606.840 17.690 607.100 18.010 ;
        RECT 603.220 2.400 603.360 17.690 ;
        RECT 603.010 -4.800 603.570 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2277.520 1283.770 2277.800 ;
      LAYER met3 ;
        RECT 1283.465 2277.810 1283.795 2277.825 ;
        RECT 1283.465 2277.760 1300.420 2277.810 ;
        RECT 1283.465 2277.510 1304.000 2277.760 ;
        RECT 1283.465 2277.495 1283.795 2277.510 ;
        RECT 1300.000 2277.160 1304.000 2277.510 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 627.050 2304.760 627.370 2304.820 ;
        RECT 1283.470 2304.760 1283.790 2304.820 ;
        RECT 627.050 2304.620 1283.790 2304.760 ;
        RECT 627.050 2304.560 627.370 2304.620 ;
        RECT 1283.470 2304.560 1283.790 2304.620 ;
        RECT 621.070 17.920 621.390 17.980 ;
        RECT 627.050 17.920 627.370 17.980 ;
        RECT 621.070 17.780 627.370 17.920 ;
        RECT 621.070 17.720 621.390 17.780 ;
        RECT 627.050 17.720 627.370 17.780 ;
      LAYER via ;
        RECT 627.080 2304.560 627.340 2304.820 ;
        RECT 1283.500 2304.560 1283.760 2304.820 ;
        RECT 621.100 17.720 621.360 17.980 ;
        RECT 627.080 17.720 627.340 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2309.435 1283.770 2309.805 ;
        RECT 1283.560 2304.850 1283.700 2309.435 ;
        RECT 627.080 2304.530 627.340 2304.850 ;
        RECT 1283.500 2304.530 1283.760 2304.850 ;
        RECT 627.140 18.010 627.280 2304.530 ;
        RECT 621.100 17.690 621.360 18.010 ;
        RECT 627.080 17.690 627.340 18.010 ;
        RECT 621.160 2.400 621.300 17.690 ;
        RECT 620.950 -4.800 621.510 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2309.480 1283.770 2309.760 ;
      LAYER met3 ;
        RECT 1283.465 2309.770 1283.795 2309.785 ;
        RECT 1283.465 2309.720 1300.420 2309.770 ;
        RECT 1283.465 2309.470 1304.000 2309.720 ;
        RECT 1283.465 2309.455 1283.795 2309.470 ;
        RECT 1300.000 2309.120 1304.000 2309.470 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 1401.040 117.230 1401.100 ;
        RECT 1283.470 1401.040 1283.790 1401.100 ;
        RECT 116.910 1400.900 1283.790 1401.040 ;
        RECT 116.910 1400.840 117.230 1400.900 ;
        RECT 1283.470 1400.840 1283.790 1400.900 ;
      LAYER via ;
        RECT 116.940 1400.840 117.200 1401.100 ;
        RECT 1283.500 1400.840 1283.760 1401.100 ;
      LAYER met2 ;
        RECT 1283.490 1406.395 1283.770 1406.765 ;
        RECT 1283.560 1401.130 1283.700 1406.395 ;
        RECT 116.940 1400.810 117.200 1401.130 ;
        RECT 1283.500 1400.810 1283.760 1401.130 ;
        RECT 117.000 17.410 117.140 1400.810 ;
        RECT 115.620 17.270 117.140 17.410 ;
        RECT 115.620 2.400 115.760 17.270 ;
        RECT 115.410 -4.800 115.970 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1406.440 1283.770 1406.720 ;
      LAYER met3 ;
        RECT 1283.465 1406.730 1283.795 1406.745 ;
        RECT 1283.465 1406.680 1300.420 1406.730 ;
        RECT 1283.465 1406.430 1304.000 1406.680 ;
        RECT 1283.465 1406.415 1283.795 1406.430 ;
        RECT 1300.000 1406.080 1304.000 1406.430 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 144.510 1449.320 144.830 1449.380 ;
        RECT 1283.470 1449.320 1283.790 1449.380 ;
        RECT 144.510 1449.180 1283.790 1449.320 ;
        RECT 144.510 1449.120 144.830 1449.180 ;
        RECT 1283.470 1449.120 1283.790 1449.180 ;
        RECT 139.450 17.920 139.770 17.980 ;
        RECT 144.510 17.920 144.830 17.980 ;
        RECT 139.450 17.780 144.830 17.920 ;
        RECT 139.450 17.720 139.770 17.780 ;
        RECT 144.510 17.720 144.830 17.780 ;
      LAYER via ;
        RECT 144.540 1449.120 144.800 1449.380 ;
        RECT 1283.500 1449.120 1283.760 1449.380 ;
        RECT 139.480 17.720 139.740 17.980 ;
        RECT 144.540 17.720 144.800 17.980 ;
      LAYER met2 ;
        RECT 144.540 1449.090 144.800 1449.410 ;
        RECT 1283.490 1449.235 1283.770 1449.605 ;
        RECT 1283.500 1449.090 1283.760 1449.235 ;
        RECT 144.600 18.010 144.740 1449.090 ;
        RECT 139.480 17.690 139.740 18.010 ;
        RECT 144.540 17.690 144.800 18.010 ;
        RECT 139.540 2.400 139.680 17.690 ;
        RECT 139.330 -4.800 139.890 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1449.280 1283.770 1449.560 ;
      LAYER met3 ;
        RECT 1283.465 1449.570 1283.795 1449.585 ;
        RECT 1283.465 1449.520 1300.420 1449.570 ;
        RECT 1283.465 1449.270 1304.000 1449.520 ;
        RECT 1283.465 1449.255 1283.795 1449.270 ;
        RECT 1300.000 1448.920 1304.000 1449.270 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1476.860 158.630 1476.920 ;
        RECT 1283.470 1476.860 1283.790 1476.920 ;
        RECT 158.310 1476.720 1283.790 1476.860 ;
        RECT 158.310 1476.660 158.630 1476.720 ;
        RECT 1283.470 1476.660 1283.790 1476.720 ;
      LAYER via ;
        RECT 158.340 1476.660 158.600 1476.920 ;
        RECT 1283.500 1476.660 1283.760 1476.920 ;
      LAYER met2 ;
        RECT 1283.490 1481.195 1283.770 1481.565 ;
        RECT 1283.560 1476.950 1283.700 1481.195 ;
        RECT 158.340 1476.630 158.600 1476.950 ;
        RECT 1283.500 1476.630 1283.760 1476.950 ;
        RECT 158.400 17.410 158.540 1476.630 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1481.240 1283.770 1481.520 ;
      LAYER met3 ;
        RECT 1283.465 1481.530 1283.795 1481.545 ;
        RECT 1283.465 1481.480 1300.420 1481.530 ;
        RECT 1283.465 1481.230 1304.000 1481.480 ;
        RECT 1283.465 1481.215 1283.795 1481.230 ;
        RECT 1300.000 1480.880 1304.000 1481.230 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 179.010 1511.200 179.330 1511.260 ;
        RECT 1283.470 1511.200 1283.790 1511.260 ;
        RECT 179.010 1511.060 1283.790 1511.200 ;
        RECT 179.010 1511.000 179.330 1511.060 ;
        RECT 1283.470 1511.000 1283.790 1511.060 ;
        RECT 174.870 17.920 175.190 17.980 ;
        RECT 179.010 17.920 179.330 17.980 ;
        RECT 174.870 17.780 179.330 17.920 ;
        RECT 174.870 17.720 175.190 17.780 ;
        RECT 179.010 17.720 179.330 17.780 ;
      LAYER via ;
        RECT 179.040 1511.000 179.300 1511.260 ;
        RECT 1283.500 1511.000 1283.760 1511.260 ;
        RECT 174.900 17.720 175.160 17.980 ;
        RECT 179.040 17.720 179.300 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1512.475 1283.770 1512.845 ;
        RECT 1283.560 1511.290 1283.700 1512.475 ;
        RECT 179.040 1510.970 179.300 1511.290 ;
        RECT 1283.500 1510.970 1283.760 1511.290 ;
        RECT 179.100 18.010 179.240 1510.970 ;
        RECT 174.900 17.690 175.160 18.010 ;
        RECT 179.040 17.690 179.300 18.010 ;
        RECT 174.960 2.400 175.100 17.690 ;
        RECT 174.750 -4.800 175.310 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1512.520 1283.770 1512.800 ;
      LAYER met3 ;
        RECT 1283.465 1512.810 1283.795 1512.825 ;
        RECT 1283.465 1512.760 1300.420 1512.810 ;
        RECT 1283.465 1512.510 1304.000 1512.760 ;
        RECT 1283.465 1512.495 1283.795 1512.510 ;
        RECT 1300.000 1512.160 1304.000 1512.510 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 192.810 1539.080 193.130 1539.140 ;
        RECT 1283.470 1539.080 1283.790 1539.140 ;
        RECT 192.810 1538.940 1283.790 1539.080 ;
        RECT 192.810 1538.880 193.130 1538.940 ;
        RECT 1283.470 1538.880 1283.790 1538.940 ;
      LAYER via ;
        RECT 192.840 1538.880 193.100 1539.140 ;
        RECT 1283.500 1538.880 1283.760 1539.140 ;
      LAYER met2 ;
        RECT 1283.490 1544.435 1283.770 1544.805 ;
        RECT 1283.560 1539.170 1283.700 1544.435 ;
        RECT 192.840 1538.850 193.100 1539.170 ;
        RECT 1283.500 1538.850 1283.760 1539.170 ;
        RECT 192.900 2.400 193.040 1538.850 ;
        RECT 192.690 -4.800 193.250 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1544.480 1283.770 1544.760 ;
      LAYER met3 ;
        RECT 1283.465 1544.770 1283.795 1544.785 ;
        RECT 1283.465 1544.720 1300.420 1544.770 ;
        RECT 1283.465 1544.470 1304.000 1544.720 ;
        RECT 1283.465 1544.455 1283.795 1544.470 ;
        RECT 1300.000 1544.120 1304.000 1544.470 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1573.420 213.830 1573.480 ;
        RECT 1283.470 1573.420 1283.790 1573.480 ;
        RECT 213.510 1573.280 1283.790 1573.420 ;
        RECT 213.510 1573.220 213.830 1573.280 ;
        RECT 1283.470 1573.220 1283.790 1573.280 ;
        RECT 210.750 17.920 211.070 17.980 ;
        RECT 213.510 17.920 213.830 17.980 ;
        RECT 210.750 17.780 213.830 17.920 ;
        RECT 210.750 17.720 211.070 17.780 ;
        RECT 213.510 17.720 213.830 17.780 ;
      LAYER via ;
        RECT 213.540 1573.220 213.800 1573.480 ;
        RECT 1283.500 1573.220 1283.760 1573.480 ;
        RECT 210.780 17.720 211.040 17.980 ;
        RECT 213.540 17.720 213.800 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1576.395 1283.770 1576.765 ;
        RECT 1283.560 1573.510 1283.700 1576.395 ;
        RECT 213.540 1573.190 213.800 1573.510 ;
        RECT 1283.500 1573.190 1283.760 1573.510 ;
        RECT 213.600 18.010 213.740 1573.190 ;
        RECT 210.780 17.690 211.040 18.010 ;
        RECT 213.540 17.690 213.800 18.010 ;
        RECT 210.840 2.400 210.980 17.690 ;
        RECT 210.630 -4.800 211.190 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1576.440 1283.770 1576.720 ;
      LAYER met3 ;
        RECT 1283.465 1576.730 1283.795 1576.745 ;
        RECT 1283.465 1576.680 1300.420 1576.730 ;
        RECT 1283.465 1576.430 1304.000 1576.680 ;
        RECT 1283.465 1576.415 1283.795 1576.430 ;
        RECT 1300.000 1576.080 1304.000 1576.430 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 234.210 1608.100 234.530 1608.160 ;
        RECT 1283.470 1608.100 1283.790 1608.160 ;
        RECT 234.210 1607.960 1283.790 1608.100 ;
        RECT 234.210 1607.900 234.530 1607.960 ;
        RECT 1283.470 1607.900 1283.790 1607.960 ;
        RECT 228.690 17.920 229.010 17.980 ;
        RECT 234.210 17.920 234.530 17.980 ;
        RECT 228.690 17.780 234.530 17.920 ;
        RECT 228.690 17.720 229.010 17.780 ;
        RECT 234.210 17.720 234.530 17.780 ;
      LAYER via ;
        RECT 234.240 1607.900 234.500 1608.160 ;
        RECT 1283.500 1607.900 1283.760 1608.160 ;
        RECT 228.720 17.720 228.980 17.980 ;
        RECT 234.240 17.720 234.500 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1608.355 1283.770 1608.725 ;
        RECT 1283.560 1608.190 1283.700 1608.355 ;
        RECT 234.240 1607.870 234.500 1608.190 ;
        RECT 1283.500 1607.870 1283.760 1608.190 ;
        RECT 234.300 18.010 234.440 1607.870 ;
        RECT 228.720 17.690 228.980 18.010 ;
        RECT 234.240 17.690 234.500 18.010 ;
        RECT 228.780 2.400 228.920 17.690 ;
        RECT 228.570 -4.800 229.130 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1608.400 1283.770 1608.680 ;
      LAYER met3 ;
        RECT 1283.465 1608.690 1283.795 1608.705 ;
        RECT 1283.465 1608.640 1300.420 1608.690 ;
        RECT 1283.465 1608.390 1304.000 1608.640 ;
        RECT 1283.465 1608.375 1283.795 1608.390 ;
        RECT 1300.000 1608.040 1304.000 1608.390 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 54.810 1283.740 55.130 1283.800 ;
        RECT 1283.470 1283.740 1283.790 1283.800 ;
        RECT 54.810 1283.600 1283.790 1283.740 ;
        RECT 54.810 1283.540 55.130 1283.600 ;
        RECT 1283.470 1283.540 1283.790 1283.600 ;
        RECT 50.210 17.920 50.530 17.980 ;
        RECT 54.810 17.920 55.130 17.980 ;
        RECT 50.210 17.780 55.130 17.920 ;
        RECT 50.210 17.720 50.530 17.780 ;
        RECT 54.810 17.720 55.130 17.780 ;
      LAYER via ;
        RECT 54.840 1283.540 55.100 1283.800 ;
        RECT 1283.500 1283.540 1283.760 1283.800 ;
        RECT 50.240 17.720 50.500 17.980 ;
        RECT 54.840 17.720 55.100 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1289.435 1283.770 1289.805 ;
        RECT 1283.560 1283.830 1283.700 1289.435 ;
        RECT 54.840 1283.510 55.100 1283.830 ;
        RECT 1283.500 1283.510 1283.760 1283.830 ;
        RECT 54.900 18.010 55.040 1283.510 ;
        RECT 50.240 17.690 50.500 18.010 ;
        RECT 54.840 17.690 55.100 18.010 ;
        RECT 50.300 2.400 50.440 17.690 ;
        RECT 50.090 -4.800 50.650 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1289.480 1283.770 1289.760 ;
      LAYER met3 ;
        RECT 1283.465 1289.770 1283.795 1289.785 ;
        RECT 1283.465 1289.720 1300.420 1289.770 ;
        RECT 1283.465 1289.470 1304.000 1289.720 ;
        RECT 1283.465 1289.455 1283.795 1289.470 ;
        RECT 1300.000 1289.120 1304.000 1289.470 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1649.240 255.230 1649.300 ;
        RECT 1283.470 1649.240 1283.790 1649.300 ;
        RECT 254.910 1649.100 1283.790 1649.240 ;
        RECT 254.910 1649.040 255.230 1649.100 ;
        RECT 1283.470 1649.040 1283.790 1649.100 ;
        RECT 252.610 17.920 252.930 17.980 ;
        RECT 254.910 17.920 255.230 17.980 ;
        RECT 252.610 17.780 255.230 17.920 ;
        RECT 252.610 17.720 252.930 17.780 ;
        RECT 254.910 17.720 255.230 17.780 ;
      LAYER via ;
        RECT 254.940 1649.040 255.200 1649.300 ;
        RECT 1283.500 1649.040 1283.760 1649.300 ;
        RECT 252.640 17.720 252.900 17.980 ;
        RECT 254.940 17.720 255.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1651.195 1283.770 1651.565 ;
        RECT 1283.560 1649.330 1283.700 1651.195 ;
        RECT 254.940 1649.010 255.200 1649.330 ;
        RECT 1283.500 1649.010 1283.760 1649.330 ;
        RECT 255.000 18.010 255.140 1649.010 ;
        RECT 252.640 17.690 252.900 18.010 ;
        RECT 254.940 17.690 255.200 18.010 ;
        RECT 252.700 2.400 252.840 17.690 ;
        RECT 252.490 -4.800 253.050 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1651.240 1283.770 1651.520 ;
      LAYER met3 ;
        RECT 1283.465 1651.530 1283.795 1651.545 ;
        RECT 1283.465 1651.480 1300.420 1651.530 ;
        RECT 1283.465 1651.230 1304.000 1651.480 ;
        RECT 1283.465 1651.215 1283.795 1651.230 ;
        RECT 1300.000 1650.880 1304.000 1651.230 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 275.610 1676.780 275.930 1676.840 ;
        RECT 1283.470 1676.780 1283.790 1676.840 ;
        RECT 275.610 1676.640 1283.790 1676.780 ;
        RECT 275.610 1676.580 275.930 1676.640 ;
        RECT 1283.470 1676.580 1283.790 1676.640 ;
        RECT 270.090 17.920 270.410 17.980 ;
        RECT 275.610 17.920 275.930 17.980 ;
        RECT 270.090 17.780 275.930 17.920 ;
        RECT 270.090 17.720 270.410 17.780 ;
        RECT 275.610 17.720 275.930 17.780 ;
      LAYER via ;
        RECT 275.640 1676.580 275.900 1676.840 ;
        RECT 1283.500 1676.580 1283.760 1676.840 ;
        RECT 270.120 17.720 270.380 17.980 ;
        RECT 275.640 17.720 275.900 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1682.475 1283.770 1682.845 ;
        RECT 1283.560 1676.870 1283.700 1682.475 ;
        RECT 275.640 1676.550 275.900 1676.870 ;
        RECT 1283.500 1676.550 1283.760 1676.870 ;
        RECT 275.700 18.010 275.840 1676.550 ;
        RECT 270.120 17.690 270.380 18.010 ;
        RECT 275.640 17.690 275.900 18.010 ;
        RECT 270.180 2.400 270.320 17.690 ;
        RECT 269.970 -4.800 270.530 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1682.520 1283.770 1682.800 ;
      LAYER met3 ;
        RECT 1283.465 1682.810 1283.795 1682.825 ;
        RECT 1283.465 1682.760 1300.420 1682.810 ;
        RECT 1283.465 1682.510 1304.000 1682.760 ;
        RECT 1283.465 1682.495 1283.795 1682.510 ;
        RECT 1300.000 1682.160 1304.000 1682.510 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 289.410 1711.460 289.730 1711.520 ;
        RECT 1283.470 1711.460 1283.790 1711.520 ;
        RECT 289.410 1711.320 1283.790 1711.460 ;
        RECT 289.410 1711.260 289.730 1711.320 ;
        RECT 1283.470 1711.260 1283.790 1711.320 ;
      LAYER via ;
        RECT 289.440 1711.260 289.700 1711.520 ;
        RECT 1283.500 1711.260 1283.760 1711.520 ;
      LAYER met2 ;
        RECT 1283.490 1714.435 1283.770 1714.805 ;
        RECT 1283.560 1711.550 1283.700 1714.435 ;
        RECT 289.440 1711.230 289.700 1711.550 ;
        RECT 1283.500 1711.230 1283.760 1711.550 ;
        RECT 289.500 17.410 289.640 1711.230 ;
        RECT 288.120 17.270 289.640 17.410 ;
        RECT 288.120 2.400 288.260 17.270 ;
        RECT 287.910 -4.800 288.470 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1714.480 1283.770 1714.760 ;
      LAYER met3 ;
        RECT 1283.465 1714.770 1283.795 1714.785 ;
        RECT 1283.465 1714.720 1300.420 1714.770 ;
        RECT 1283.465 1714.470 1304.000 1714.720 ;
        RECT 1283.465 1714.455 1283.795 1714.470 ;
        RECT 1300.000 1714.120 1304.000 1714.470 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 310.110 1745.800 310.430 1745.860 ;
        RECT 1283.470 1745.800 1283.790 1745.860 ;
        RECT 310.110 1745.660 1283.790 1745.800 ;
        RECT 310.110 1745.600 310.430 1745.660 ;
        RECT 1283.470 1745.600 1283.790 1745.660 ;
        RECT 305.970 17.920 306.290 17.980 ;
        RECT 310.110 17.920 310.430 17.980 ;
        RECT 305.970 17.780 310.430 17.920 ;
        RECT 305.970 17.720 306.290 17.780 ;
        RECT 310.110 17.720 310.430 17.780 ;
      LAYER via ;
        RECT 310.140 1745.600 310.400 1745.860 ;
        RECT 1283.500 1745.600 1283.760 1745.860 ;
        RECT 306.000 17.720 306.260 17.980 ;
        RECT 310.140 17.720 310.400 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1746.395 1283.770 1746.765 ;
        RECT 1283.560 1745.890 1283.700 1746.395 ;
        RECT 310.140 1745.570 310.400 1745.890 ;
        RECT 1283.500 1745.570 1283.760 1745.890 ;
        RECT 310.200 18.010 310.340 1745.570 ;
        RECT 306.000 17.690 306.260 18.010 ;
        RECT 310.140 17.690 310.400 18.010 ;
        RECT 306.060 2.400 306.200 17.690 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1746.440 1283.770 1746.720 ;
      LAYER met3 ;
        RECT 1283.465 1746.730 1283.795 1746.745 ;
        RECT 1283.465 1746.680 1300.420 1746.730 ;
        RECT 1283.465 1746.430 1304.000 1746.680 ;
        RECT 1283.465 1746.415 1283.795 1746.430 ;
        RECT 1300.000 1746.080 1304.000 1746.430 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 323.910 1773.680 324.230 1773.740 ;
        RECT 1283.470 1773.680 1283.790 1773.740 ;
        RECT 323.910 1773.540 1283.790 1773.680 ;
        RECT 323.910 1773.480 324.230 1773.540 ;
        RECT 1283.470 1773.480 1283.790 1773.540 ;
      LAYER via ;
        RECT 323.940 1773.480 324.200 1773.740 ;
        RECT 1283.500 1773.480 1283.760 1773.740 ;
      LAYER met2 ;
        RECT 1283.490 1778.355 1283.770 1778.725 ;
        RECT 1283.560 1773.770 1283.700 1778.355 ;
        RECT 323.940 1773.450 324.200 1773.770 ;
        RECT 1283.500 1773.450 1283.760 1773.770 ;
        RECT 324.000 2.400 324.140 1773.450 ;
        RECT 323.790 -4.800 324.350 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1778.400 1283.770 1778.680 ;
      LAYER met3 ;
        RECT 1283.465 1778.690 1283.795 1778.705 ;
        RECT 1283.465 1778.640 1300.420 1778.690 ;
        RECT 1283.465 1778.390 1304.000 1778.640 ;
        RECT 1283.465 1778.375 1283.795 1778.390 ;
        RECT 1300.000 1778.040 1304.000 1778.390 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 344.610 1808.020 344.930 1808.080 ;
        RECT 1283.470 1808.020 1283.790 1808.080 ;
        RECT 344.610 1807.880 1283.790 1808.020 ;
        RECT 344.610 1807.820 344.930 1807.880 ;
        RECT 1283.470 1807.820 1283.790 1807.880 ;
        RECT 341.390 17.920 341.710 17.980 ;
        RECT 344.610 17.920 344.930 17.980 ;
        RECT 341.390 17.780 344.930 17.920 ;
        RECT 341.390 17.720 341.710 17.780 ;
        RECT 344.610 17.720 344.930 17.780 ;
      LAYER via ;
        RECT 344.640 1807.820 344.900 1808.080 ;
        RECT 1283.500 1807.820 1283.760 1808.080 ;
        RECT 341.420 17.720 341.680 17.980 ;
        RECT 344.640 17.720 344.900 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1810.315 1283.770 1810.685 ;
        RECT 1283.560 1808.110 1283.700 1810.315 ;
        RECT 344.640 1807.790 344.900 1808.110 ;
        RECT 1283.500 1807.790 1283.760 1808.110 ;
        RECT 344.700 18.010 344.840 1807.790 ;
        RECT 341.420 17.690 341.680 18.010 ;
        RECT 344.640 17.690 344.900 18.010 ;
        RECT 341.480 2.400 341.620 17.690 ;
        RECT 341.270 -4.800 341.830 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1810.360 1283.770 1810.640 ;
      LAYER met3 ;
        RECT 1283.465 1810.650 1283.795 1810.665 ;
        RECT 1283.465 1810.600 1300.420 1810.650 ;
        RECT 1283.465 1810.350 1304.000 1810.600 ;
        RECT 1283.465 1810.335 1283.795 1810.350 ;
        RECT 1300.000 1810.000 1304.000 1810.350 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 1842.700 365.170 1842.760 ;
        RECT 1283.470 1842.700 1283.790 1842.760 ;
        RECT 364.850 1842.560 1283.790 1842.700 ;
        RECT 364.850 1842.500 365.170 1842.560 ;
        RECT 1283.470 1842.500 1283.790 1842.560 ;
        RECT 359.330 17.920 359.650 17.980 ;
        RECT 364.850 17.920 365.170 17.980 ;
        RECT 359.330 17.780 365.170 17.920 ;
        RECT 359.330 17.720 359.650 17.780 ;
        RECT 364.850 17.720 365.170 17.780 ;
      LAYER via ;
        RECT 364.880 1842.500 365.140 1842.760 ;
        RECT 1283.500 1842.500 1283.760 1842.760 ;
        RECT 359.360 17.720 359.620 17.980 ;
        RECT 364.880 17.720 365.140 17.980 ;
      LAYER met2 ;
        RECT 364.880 1842.470 365.140 1842.790 ;
        RECT 1283.500 1842.645 1283.760 1842.790 ;
        RECT 364.940 18.010 365.080 1842.470 ;
        RECT 1283.490 1842.275 1283.770 1842.645 ;
        RECT 359.360 17.690 359.620 18.010 ;
        RECT 364.880 17.690 365.140 18.010 ;
        RECT 359.420 2.400 359.560 17.690 ;
        RECT 359.210 -4.800 359.770 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1842.320 1283.770 1842.600 ;
      LAYER met3 ;
        RECT 1283.465 1842.610 1283.795 1842.625 ;
        RECT 1283.465 1842.560 1300.420 1842.610 ;
        RECT 1283.465 1842.310 1304.000 1842.560 ;
        RECT 1283.465 1842.295 1283.795 1842.310 ;
        RECT 1300.000 1841.960 1304.000 1842.310 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 379.110 1870.240 379.430 1870.300 ;
        RECT 1283.470 1870.240 1283.790 1870.300 ;
        RECT 379.110 1870.100 1283.790 1870.240 ;
        RECT 379.110 1870.040 379.430 1870.100 ;
        RECT 1283.470 1870.040 1283.790 1870.100 ;
      LAYER via ;
        RECT 379.140 1870.040 379.400 1870.300 ;
        RECT 1283.500 1870.040 1283.760 1870.300 ;
      LAYER met2 ;
        RECT 1283.490 1874.235 1283.770 1874.605 ;
        RECT 1283.560 1870.330 1283.700 1874.235 ;
        RECT 379.140 1870.010 379.400 1870.330 ;
        RECT 1283.500 1870.010 1283.760 1870.330 ;
        RECT 379.200 17.410 379.340 1870.010 ;
        RECT 377.360 17.270 379.340 17.410 ;
        RECT 377.360 2.400 377.500 17.270 ;
        RECT 377.150 -4.800 377.710 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1874.280 1283.770 1874.560 ;
      LAYER met3 ;
        RECT 1283.465 1874.570 1283.795 1874.585 ;
        RECT 1283.465 1874.520 1300.420 1874.570 ;
        RECT 1283.465 1874.270 1304.000 1874.520 ;
        RECT 1283.465 1874.255 1283.795 1874.270 ;
        RECT 1300.000 1873.920 1304.000 1874.270 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 399.810 1904.580 400.130 1904.640 ;
        RECT 1283.470 1904.580 1283.790 1904.640 ;
        RECT 399.810 1904.440 1283.790 1904.580 ;
        RECT 399.810 1904.380 400.130 1904.440 ;
        RECT 1283.470 1904.380 1283.790 1904.440 ;
        RECT 395.210 17.920 395.530 17.980 ;
        RECT 399.810 17.920 400.130 17.980 ;
        RECT 395.210 17.780 400.130 17.920 ;
        RECT 395.210 17.720 395.530 17.780 ;
        RECT 399.810 17.720 400.130 17.780 ;
      LAYER via ;
        RECT 399.840 1904.380 400.100 1904.640 ;
        RECT 1283.500 1904.380 1283.760 1904.640 ;
        RECT 395.240 17.720 395.500 17.980 ;
        RECT 399.840 17.720 400.100 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1905.515 1283.770 1905.885 ;
        RECT 1283.560 1904.670 1283.700 1905.515 ;
        RECT 399.840 1904.350 400.100 1904.670 ;
        RECT 1283.500 1904.350 1283.760 1904.670 ;
        RECT 399.900 18.010 400.040 1904.350 ;
        RECT 395.240 17.690 395.500 18.010 ;
        RECT 399.840 17.690 400.100 18.010 ;
        RECT 395.300 2.400 395.440 17.690 ;
        RECT 395.090 -4.800 395.650 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1905.560 1283.770 1905.840 ;
      LAYER met3 ;
        RECT 1283.465 1905.850 1283.795 1905.865 ;
        RECT 1283.465 1905.800 1300.420 1905.850 ;
        RECT 1283.465 1905.550 1304.000 1905.800 ;
        RECT 1283.465 1905.535 1283.795 1905.550 ;
        RECT 1300.000 1905.200 1304.000 1905.550 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 413.610 1932.120 413.930 1932.180 ;
        RECT 1283.470 1932.120 1283.790 1932.180 ;
        RECT 413.610 1931.980 1283.790 1932.120 ;
        RECT 413.610 1931.920 413.930 1931.980 ;
        RECT 1283.470 1931.920 1283.790 1931.980 ;
      LAYER via ;
        RECT 413.640 1931.920 413.900 1932.180 ;
        RECT 1283.500 1931.920 1283.760 1932.180 ;
      LAYER met2 ;
        RECT 1283.490 1937.475 1283.770 1937.845 ;
        RECT 1283.560 1932.210 1283.700 1937.475 ;
        RECT 413.640 1931.890 413.900 1932.210 ;
        RECT 1283.500 1931.890 1283.760 1932.210 ;
        RECT 413.700 17.410 413.840 1931.890 ;
        RECT 413.240 17.270 413.840 17.410 ;
        RECT 413.240 2.400 413.380 17.270 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1937.520 1283.770 1937.800 ;
      LAYER met3 ;
        RECT 1283.465 1937.810 1283.795 1937.825 ;
        RECT 1283.465 1937.760 1300.420 1937.810 ;
        RECT 1283.465 1937.510 1304.000 1937.760 ;
        RECT 1283.465 1937.495 1283.795 1937.510 ;
        RECT 1300.000 1937.160 1304.000 1937.510 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 75.510 1332.020 75.830 1332.080 ;
        RECT 1283.470 1332.020 1283.790 1332.080 ;
        RECT 75.510 1331.880 1283.790 1332.020 ;
        RECT 75.510 1331.820 75.830 1331.880 ;
        RECT 1283.470 1331.820 1283.790 1331.880 ;
      LAYER via ;
        RECT 75.540 1331.820 75.800 1332.080 ;
        RECT 1283.500 1331.820 1283.760 1332.080 ;
      LAYER met2 ;
        RECT 1283.490 1332.275 1283.770 1332.645 ;
        RECT 1283.560 1332.110 1283.700 1332.275 ;
        RECT 75.540 1331.790 75.800 1332.110 ;
        RECT 1283.500 1331.790 1283.760 1332.110 ;
        RECT 75.600 17.410 75.740 1331.790 ;
        RECT 74.220 17.270 75.740 17.410 ;
        RECT 74.220 2.400 74.360 17.270 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1332.320 1283.770 1332.600 ;
      LAYER met3 ;
        RECT 1283.465 1332.610 1283.795 1332.625 ;
        RECT 1283.465 1332.560 1300.420 1332.610 ;
        RECT 1283.465 1332.310 1304.000 1332.560 ;
        RECT 1283.465 1332.295 1283.795 1332.310 ;
        RECT 1300.000 1331.960 1304.000 1332.310 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 434.310 1966.800 434.630 1966.860 ;
        RECT 1283.470 1966.800 1283.790 1966.860 ;
        RECT 434.310 1966.660 1283.790 1966.800 ;
        RECT 434.310 1966.600 434.630 1966.660 ;
        RECT 1283.470 1966.600 1283.790 1966.660 ;
        RECT 430.630 17.920 430.950 17.980 ;
        RECT 434.310 17.920 434.630 17.980 ;
        RECT 430.630 17.780 434.630 17.920 ;
        RECT 430.630 17.720 430.950 17.780 ;
        RECT 434.310 17.720 434.630 17.780 ;
      LAYER via ;
        RECT 434.340 1966.600 434.600 1966.860 ;
        RECT 1283.500 1966.600 1283.760 1966.860 ;
        RECT 430.660 17.720 430.920 17.980 ;
        RECT 434.340 17.720 434.600 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1969.435 1283.770 1969.805 ;
        RECT 1283.560 1966.890 1283.700 1969.435 ;
        RECT 434.340 1966.570 434.600 1966.890 ;
        RECT 1283.500 1966.570 1283.760 1966.890 ;
        RECT 434.400 18.010 434.540 1966.570 ;
        RECT 430.660 17.690 430.920 18.010 ;
        RECT 434.340 17.690 434.600 18.010 ;
        RECT 430.720 2.400 430.860 17.690 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1969.480 1283.770 1969.760 ;
      LAYER met3 ;
        RECT 1283.465 1969.770 1283.795 1969.785 ;
        RECT 1283.465 1969.720 1300.420 1969.770 ;
        RECT 1283.465 1969.470 1304.000 1969.720 ;
        RECT 1283.465 1969.455 1283.795 1969.470 ;
        RECT 1300.000 1969.120 1304.000 1969.470 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 454.550 2001.140 454.870 2001.200 ;
        RECT 1283.470 2001.140 1283.790 2001.200 ;
        RECT 454.550 2001.000 1283.790 2001.140 ;
        RECT 454.550 2000.940 454.870 2001.000 ;
        RECT 1283.470 2000.940 1283.790 2001.000 ;
        RECT 448.570 17.920 448.890 17.980 ;
        RECT 454.550 17.920 454.870 17.980 ;
        RECT 448.570 17.780 454.870 17.920 ;
        RECT 448.570 17.720 448.890 17.780 ;
        RECT 454.550 17.720 454.870 17.780 ;
      LAYER via ;
        RECT 454.580 2000.940 454.840 2001.200 ;
        RECT 1283.500 2000.940 1283.760 2001.200 ;
        RECT 448.600 17.720 448.860 17.980 ;
        RECT 454.580 17.720 454.840 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2001.395 1283.770 2001.765 ;
        RECT 1283.560 2001.230 1283.700 2001.395 ;
        RECT 454.580 2000.910 454.840 2001.230 ;
        RECT 1283.500 2000.910 1283.760 2001.230 ;
        RECT 454.640 18.010 454.780 2000.910 ;
        RECT 448.600 17.690 448.860 18.010 ;
        RECT 454.580 17.690 454.840 18.010 ;
        RECT 448.660 2.400 448.800 17.690 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2001.440 1283.770 2001.720 ;
      LAYER met3 ;
        RECT 1283.465 2001.730 1283.795 2001.745 ;
        RECT 1283.465 2001.680 1300.420 2001.730 ;
        RECT 1283.465 2001.430 1304.000 2001.680 ;
        RECT 1283.465 2001.415 1283.795 2001.430 ;
        RECT 1300.000 2001.080 1304.000 2001.430 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 468.810 2028.680 469.130 2028.740 ;
        RECT 1283.470 2028.680 1283.790 2028.740 ;
        RECT 468.810 2028.540 1283.790 2028.680 ;
        RECT 468.810 2028.480 469.130 2028.540 ;
        RECT 1283.470 2028.480 1283.790 2028.540 ;
        RECT 466.510 17.920 466.830 17.980 ;
        RECT 468.810 17.920 469.130 17.980 ;
        RECT 466.510 17.780 469.130 17.920 ;
        RECT 466.510 17.720 466.830 17.780 ;
        RECT 468.810 17.720 469.130 17.780 ;
      LAYER via ;
        RECT 468.840 2028.480 469.100 2028.740 ;
        RECT 1283.500 2028.480 1283.760 2028.740 ;
        RECT 466.540 17.720 466.800 17.980 ;
        RECT 468.840 17.720 469.100 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2033.355 1283.770 2033.725 ;
        RECT 1283.560 2028.770 1283.700 2033.355 ;
        RECT 468.840 2028.450 469.100 2028.770 ;
        RECT 1283.500 2028.450 1283.760 2028.770 ;
        RECT 468.900 18.010 469.040 2028.450 ;
        RECT 466.540 17.690 466.800 18.010 ;
        RECT 468.840 17.690 469.100 18.010 ;
        RECT 466.600 2.400 466.740 17.690 ;
        RECT 466.390 -4.800 466.950 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2033.400 1283.770 2033.680 ;
      LAYER met3 ;
        RECT 1283.465 2033.690 1283.795 2033.705 ;
        RECT 1283.465 2033.640 1300.420 2033.690 ;
        RECT 1283.465 2033.390 1304.000 2033.640 ;
        RECT 1283.465 2033.375 1283.795 2033.390 ;
        RECT 1300.000 2033.040 1304.000 2033.390 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 489.510 2063.360 489.830 2063.420 ;
        RECT 1283.470 2063.360 1283.790 2063.420 ;
        RECT 489.510 2063.220 1283.790 2063.360 ;
        RECT 489.510 2063.160 489.830 2063.220 ;
        RECT 1283.470 2063.160 1283.790 2063.220 ;
        RECT 484.450 17.920 484.770 17.980 ;
        RECT 489.510 17.920 489.830 17.980 ;
        RECT 484.450 17.780 489.830 17.920 ;
        RECT 484.450 17.720 484.770 17.780 ;
        RECT 489.510 17.720 489.830 17.780 ;
      LAYER via ;
        RECT 489.540 2063.160 489.800 2063.420 ;
        RECT 1283.500 2063.160 1283.760 2063.420 ;
        RECT 484.480 17.720 484.740 17.980 ;
        RECT 489.540 17.720 489.800 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2065.315 1283.770 2065.685 ;
        RECT 1283.560 2063.450 1283.700 2065.315 ;
        RECT 489.540 2063.130 489.800 2063.450 ;
        RECT 1283.500 2063.130 1283.760 2063.450 ;
        RECT 489.600 18.010 489.740 2063.130 ;
        RECT 484.480 17.690 484.740 18.010 ;
        RECT 489.540 17.690 489.800 18.010 ;
        RECT 484.540 2.400 484.680 17.690 ;
        RECT 484.330 -4.800 484.890 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2065.360 1283.770 2065.640 ;
      LAYER met3 ;
        RECT 1283.465 2065.650 1283.795 2065.665 ;
        RECT 1283.465 2065.600 1300.420 2065.650 ;
        RECT 1283.465 2065.350 1304.000 2065.600 ;
        RECT 1283.465 2065.335 1283.795 2065.350 ;
        RECT 1300.000 2065.000 1304.000 2065.350 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 2090.900 503.630 2090.960 ;
        RECT 1283.470 2090.900 1283.790 2090.960 ;
        RECT 503.310 2090.760 1283.790 2090.900 ;
        RECT 503.310 2090.700 503.630 2090.760 ;
        RECT 1283.470 2090.700 1283.790 2090.760 ;
      LAYER via ;
        RECT 503.340 2090.700 503.600 2090.960 ;
        RECT 1283.500 2090.700 1283.760 2090.960 ;
      LAYER met2 ;
        RECT 1283.490 2097.275 1283.770 2097.645 ;
        RECT 1283.560 2090.990 1283.700 2097.275 ;
        RECT 503.340 2090.670 503.600 2090.990 ;
        RECT 1283.500 2090.670 1283.760 2090.990 ;
        RECT 503.400 17.410 503.540 2090.670 ;
        RECT 502.480 17.270 503.540 17.410 ;
        RECT 502.480 2.400 502.620 17.270 ;
        RECT 502.270 -4.800 502.830 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2097.320 1283.770 2097.600 ;
      LAYER met3 ;
        RECT 1283.465 2097.610 1283.795 2097.625 ;
        RECT 1283.465 2097.560 1300.420 2097.610 ;
        RECT 1283.465 2097.310 1304.000 2097.560 ;
        RECT 1283.465 2097.295 1283.795 2097.310 ;
        RECT 1300.000 2096.960 1304.000 2097.310 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 524.010 2125.580 524.330 2125.640 ;
        RECT 1283.470 2125.580 1283.790 2125.640 ;
        RECT 524.010 2125.440 1283.790 2125.580 ;
        RECT 524.010 2125.380 524.330 2125.440 ;
        RECT 1283.470 2125.380 1283.790 2125.440 ;
        RECT 519.870 17.920 520.190 17.980 ;
        RECT 524.010 17.920 524.330 17.980 ;
        RECT 519.870 17.780 524.330 17.920 ;
        RECT 519.870 17.720 520.190 17.780 ;
        RECT 524.010 17.720 524.330 17.780 ;
      LAYER via ;
        RECT 524.040 2125.380 524.300 2125.640 ;
        RECT 1283.500 2125.380 1283.760 2125.640 ;
        RECT 519.900 17.720 520.160 17.980 ;
        RECT 524.040 17.720 524.300 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2128.555 1283.770 2128.925 ;
        RECT 1283.560 2125.670 1283.700 2128.555 ;
        RECT 524.040 2125.350 524.300 2125.670 ;
        RECT 1283.500 2125.350 1283.760 2125.670 ;
        RECT 524.100 18.010 524.240 2125.350 ;
        RECT 519.900 17.690 520.160 18.010 ;
        RECT 524.040 17.690 524.300 18.010 ;
        RECT 519.960 2.400 520.100 17.690 ;
        RECT 519.750 -4.800 520.310 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2128.600 1283.770 2128.880 ;
      LAYER met3 ;
        RECT 1283.465 2128.890 1283.795 2128.905 ;
        RECT 1283.465 2128.840 1300.420 2128.890 ;
        RECT 1283.465 2128.590 1304.000 2128.840 ;
        RECT 1283.465 2128.575 1283.795 2128.590 ;
        RECT 1300.000 2128.240 1304.000 2128.590 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 2159.920 538.130 2159.980 ;
        RECT 1283.470 2159.920 1283.790 2159.980 ;
        RECT 537.810 2159.780 1283.790 2159.920 ;
        RECT 537.810 2159.720 538.130 2159.780 ;
        RECT 1283.470 2159.720 1283.790 2159.780 ;
      LAYER via ;
        RECT 537.840 2159.720 538.100 2159.980 ;
        RECT 1283.500 2159.720 1283.760 2159.980 ;
      LAYER met2 ;
        RECT 1283.490 2160.515 1283.770 2160.885 ;
        RECT 1283.560 2160.010 1283.700 2160.515 ;
        RECT 537.840 2159.690 538.100 2160.010 ;
        RECT 1283.500 2159.690 1283.760 2160.010 ;
        RECT 537.900 2.400 538.040 2159.690 ;
        RECT 537.690 -4.800 538.250 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2160.560 1283.770 2160.840 ;
      LAYER met3 ;
        RECT 1283.465 2160.850 1283.795 2160.865 ;
        RECT 1283.465 2160.800 1300.420 2160.850 ;
        RECT 1283.465 2160.550 1304.000 2160.800 ;
        RECT 1283.465 2160.535 1283.795 2160.550 ;
        RECT 1300.000 2160.200 1304.000 2160.550 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 558.510 2187.460 558.830 2187.520 ;
        RECT 1283.470 2187.460 1283.790 2187.520 ;
        RECT 558.510 2187.320 1283.790 2187.460 ;
        RECT 558.510 2187.260 558.830 2187.320 ;
        RECT 1283.470 2187.260 1283.790 2187.320 ;
        RECT 555.750 17.920 556.070 17.980 ;
        RECT 558.510 17.920 558.830 17.980 ;
        RECT 555.750 17.780 558.830 17.920 ;
        RECT 555.750 17.720 556.070 17.780 ;
        RECT 558.510 17.720 558.830 17.780 ;
      LAYER via ;
        RECT 558.540 2187.260 558.800 2187.520 ;
        RECT 1283.500 2187.260 1283.760 2187.520 ;
        RECT 555.780 17.720 556.040 17.980 ;
        RECT 558.540 17.720 558.800 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2192.475 1283.770 2192.845 ;
        RECT 1283.560 2187.550 1283.700 2192.475 ;
        RECT 558.540 2187.230 558.800 2187.550 ;
        RECT 1283.500 2187.230 1283.760 2187.550 ;
        RECT 558.600 18.010 558.740 2187.230 ;
        RECT 555.780 17.690 556.040 18.010 ;
        RECT 558.540 17.690 558.800 18.010 ;
        RECT 555.840 2.400 555.980 17.690 ;
        RECT 555.630 -4.800 556.190 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2192.520 1283.770 2192.800 ;
      LAYER met3 ;
        RECT 1283.465 2192.810 1283.795 2192.825 ;
        RECT 1283.465 2192.760 1300.420 2192.810 ;
        RECT 1283.465 2192.510 1304.000 2192.760 ;
        RECT 1283.465 2192.495 1283.795 2192.510 ;
        RECT 1300.000 2192.160 1304.000 2192.510 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 579.210 2222.140 579.530 2222.200 ;
        RECT 1283.470 2222.140 1283.790 2222.200 ;
        RECT 579.210 2222.000 1283.790 2222.140 ;
        RECT 579.210 2221.940 579.530 2222.000 ;
        RECT 1283.470 2221.940 1283.790 2222.000 ;
        RECT 573.690 17.920 574.010 17.980 ;
        RECT 579.210 17.920 579.530 17.980 ;
        RECT 573.690 17.780 579.530 17.920 ;
        RECT 573.690 17.720 574.010 17.780 ;
        RECT 579.210 17.720 579.530 17.780 ;
      LAYER via ;
        RECT 579.240 2221.940 579.500 2222.200 ;
        RECT 1283.500 2221.940 1283.760 2222.200 ;
        RECT 573.720 17.720 573.980 17.980 ;
        RECT 579.240 17.720 579.500 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2224.435 1283.770 2224.805 ;
        RECT 1283.560 2222.230 1283.700 2224.435 ;
        RECT 579.240 2221.910 579.500 2222.230 ;
        RECT 1283.500 2221.910 1283.760 2222.230 ;
        RECT 579.300 18.010 579.440 2221.910 ;
        RECT 573.720 17.690 573.980 18.010 ;
        RECT 579.240 17.690 579.500 18.010 ;
        RECT 573.780 2.400 573.920 17.690 ;
        RECT 573.570 -4.800 574.130 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2224.480 1283.770 2224.760 ;
      LAYER met3 ;
        RECT 1283.465 2224.770 1283.795 2224.785 ;
        RECT 1283.465 2224.720 1300.420 2224.770 ;
        RECT 1283.465 2224.470 1304.000 2224.720 ;
        RECT 1283.465 2224.455 1283.795 2224.470 ;
        RECT 1300.000 2224.120 1304.000 2224.470 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 2256.480 593.330 2256.540 ;
        RECT 1283.470 2256.480 1283.790 2256.540 ;
        RECT 593.010 2256.340 1283.790 2256.480 ;
        RECT 593.010 2256.280 593.330 2256.340 ;
        RECT 1283.470 2256.280 1283.790 2256.340 ;
      LAYER via ;
        RECT 593.040 2256.280 593.300 2256.540 ;
        RECT 1283.500 2256.280 1283.760 2256.540 ;
      LAYER met2 ;
        RECT 593.040 2256.250 593.300 2256.570 ;
        RECT 1283.490 2256.395 1283.770 2256.765 ;
        RECT 1283.500 2256.250 1283.760 2256.395 ;
        RECT 593.100 17.410 593.240 2256.250 ;
        RECT 591.260 17.270 593.240 17.410 ;
        RECT 591.260 2.400 591.400 17.270 ;
        RECT 591.050 -4.800 591.610 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2256.440 1283.770 2256.720 ;
      LAYER met3 ;
        RECT 1283.465 2256.730 1283.795 2256.745 ;
        RECT 1283.465 2256.680 1300.420 2256.730 ;
        RECT 1283.465 2256.430 1304.000 2256.680 ;
        RECT 1283.465 2256.415 1283.795 2256.430 ;
        RECT 1300.000 2256.080 1304.000 2256.430 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 103.110 1373.500 103.430 1373.560 ;
        RECT 1283.470 1373.500 1283.790 1373.560 ;
        RECT 103.110 1373.360 1283.790 1373.500 ;
        RECT 103.110 1373.300 103.430 1373.360 ;
        RECT 1283.470 1373.300 1283.790 1373.360 ;
        RECT 97.590 17.920 97.910 17.980 ;
        RECT 103.110 17.920 103.430 17.980 ;
        RECT 97.590 17.780 103.430 17.920 ;
        RECT 97.590 17.720 97.910 17.780 ;
        RECT 103.110 17.720 103.430 17.780 ;
      LAYER via ;
        RECT 103.140 1373.300 103.400 1373.560 ;
        RECT 1283.500 1373.300 1283.760 1373.560 ;
        RECT 97.620 17.720 97.880 17.980 ;
        RECT 103.140 17.720 103.400 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1374.435 1283.770 1374.805 ;
        RECT 1283.560 1373.590 1283.700 1374.435 ;
        RECT 103.140 1373.270 103.400 1373.590 ;
        RECT 1283.500 1373.270 1283.760 1373.590 ;
        RECT 103.200 18.010 103.340 1373.270 ;
        RECT 97.620 17.690 97.880 18.010 ;
        RECT 103.140 17.690 103.400 18.010 ;
        RECT 97.680 2.400 97.820 17.690 ;
        RECT 97.470 -4.800 98.030 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1374.480 1283.770 1374.760 ;
      LAYER met3 ;
        RECT 1283.465 1374.770 1283.795 1374.785 ;
        RECT 1283.465 1374.720 1300.420 1374.770 ;
        RECT 1283.465 1374.470 1304.000 1374.720 ;
        RECT 1283.465 1374.455 1283.795 1374.470 ;
        RECT 1300.000 1374.120 1304.000 1374.470 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 613.710 2284.020 614.030 2284.080 ;
        RECT 1283.470 2284.020 1283.790 2284.080 ;
        RECT 613.710 2283.880 1283.790 2284.020 ;
        RECT 613.710 2283.820 614.030 2283.880 ;
        RECT 1283.470 2283.820 1283.790 2283.880 ;
        RECT 609.110 17.920 609.430 17.980 ;
        RECT 613.710 17.920 614.030 17.980 ;
        RECT 609.110 17.780 614.030 17.920 ;
        RECT 609.110 17.720 609.430 17.780 ;
        RECT 613.710 17.720 614.030 17.780 ;
      LAYER via ;
        RECT 613.740 2283.820 614.000 2284.080 ;
        RECT 1283.500 2283.820 1283.760 2284.080 ;
        RECT 609.140 17.720 609.400 17.980 ;
        RECT 613.740 17.720 614.000 17.980 ;
      LAYER met2 ;
        RECT 1283.490 2288.355 1283.770 2288.725 ;
        RECT 1283.560 2284.110 1283.700 2288.355 ;
        RECT 613.740 2283.790 614.000 2284.110 ;
        RECT 1283.500 2283.790 1283.760 2284.110 ;
        RECT 613.800 18.010 613.940 2283.790 ;
        RECT 609.140 17.690 609.400 18.010 ;
        RECT 613.740 17.690 614.000 18.010 ;
        RECT 609.200 2.400 609.340 17.690 ;
        RECT 608.990 -4.800 609.550 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2288.400 1283.770 2288.680 ;
      LAYER met3 ;
        RECT 1283.465 2288.690 1283.795 2288.705 ;
        RECT 1283.465 2288.640 1300.420 2288.690 ;
        RECT 1283.465 2288.390 1304.000 2288.640 ;
        RECT 1283.465 2288.375 1283.795 2288.390 ;
        RECT 1300.000 2288.040 1304.000 2288.390 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 2318.700 627.830 2318.760 ;
        RECT 1283.470 2318.700 1283.790 2318.760 ;
        RECT 627.510 2318.560 1283.790 2318.700 ;
        RECT 627.510 2318.500 627.830 2318.560 ;
        RECT 1283.470 2318.500 1283.790 2318.560 ;
      LAYER via ;
        RECT 627.540 2318.500 627.800 2318.760 ;
        RECT 1283.500 2318.500 1283.760 2318.760 ;
      LAYER met2 ;
        RECT 1283.490 2320.315 1283.770 2320.685 ;
        RECT 1283.560 2318.790 1283.700 2320.315 ;
        RECT 627.540 2318.470 627.800 2318.790 ;
        RECT 1283.500 2318.470 1283.760 2318.790 ;
        RECT 627.600 17.410 627.740 2318.470 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
      LAYER via2 ;
        RECT 1283.490 2320.360 1283.770 2320.640 ;
      LAYER met3 ;
        RECT 1283.465 2320.650 1283.795 2320.665 ;
        RECT 1283.465 2320.600 1300.420 2320.650 ;
        RECT 1283.465 2320.350 1304.000 2320.600 ;
        RECT 1283.465 2320.335 1283.795 2320.350 ;
        RECT 1300.000 2320.000 1304.000 2320.350 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 123.810 1414.640 124.130 1414.700 ;
        RECT 1283.470 1414.640 1283.790 1414.700 ;
        RECT 123.810 1414.500 1283.790 1414.640 ;
        RECT 123.810 1414.440 124.130 1414.500 ;
        RECT 1283.470 1414.440 1283.790 1414.500 ;
        RECT 121.510 17.920 121.830 17.980 ;
        RECT 123.810 17.920 124.130 17.980 ;
        RECT 121.510 17.780 124.130 17.920 ;
        RECT 121.510 17.720 121.830 17.780 ;
        RECT 123.810 17.720 124.130 17.780 ;
      LAYER via ;
        RECT 123.840 1414.440 124.100 1414.700 ;
        RECT 1283.500 1414.440 1283.760 1414.700 ;
        RECT 121.540 17.720 121.800 17.980 ;
        RECT 123.840 17.720 124.100 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1417.275 1283.770 1417.645 ;
        RECT 1283.560 1414.730 1283.700 1417.275 ;
        RECT 123.840 1414.410 124.100 1414.730 ;
        RECT 1283.500 1414.410 1283.760 1414.730 ;
        RECT 123.900 18.010 124.040 1414.410 ;
        RECT 121.540 17.690 121.800 18.010 ;
        RECT 123.840 17.690 124.100 18.010 ;
        RECT 121.600 2.400 121.740 17.690 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1417.320 1283.770 1417.600 ;
      LAYER met3 ;
        RECT 1283.465 1417.610 1283.795 1417.625 ;
        RECT 1283.465 1417.560 1300.420 1417.610 ;
        RECT 1283.465 1417.310 1304.000 1417.560 ;
        RECT 1283.465 1417.295 1283.795 1417.310 ;
        RECT 1300.000 1416.960 1304.000 1417.310 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 150.950 1456.120 151.270 1456.180 ;
        RECT 1283.470 1456.120 1283.790 1456.180 ;
        RECT 150.950 1455.980 1283.790 1456.120 ;
        RECT 150.950 1455.920 151.270 1455.980 ;
        RECT 1283.470 1455.920 1283.790 1455.980 ;
        RECT 145.430 17.920 145.750 17.980 ;
        RECT 150.950 17.920 151.270 17.980 ;
        RECT 145.430 17.780 151.270 17.920 ;
        RECT 145.430 17.720 145.750 17.780 ;
        RECT 150.950 17.720 151.270 17.780 ;
      LAYER via ;
        RECT 150.980 1455.920 151.240 1456.180 ;
        RECT 1283.500 1455.920 1283.760 1456.180 ;
        RECT 145.460 17.720 145.720 17.980 ;
        RECT 150.980 17.720 151.240 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1459.435 1283.770 1459.805 ;
        RECT 1283.560 1456.210 1283.700 1459.435 ;
        RECT 150.980 1455.890 151.240 1456.210 ;
        RECT 1283.500 1455.890 1283.760 1456.210 ;
        RECT 151.040 18.010 151.180 1455.890 ;
        RECT 145.460 17.690 145.720 18.010 ;
        RECT 150.980 17.690 151.240 18.010 ;
        RECT 145.520 2.400 145.660 17.690 ;
        RECT 145.310 -4.800 145.870 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1459.480 1283.770 1459.760 ;
      LAYER met3 ;
        RECT 1283.465 1459.770 1283.795 1459.785 ;
        RECT 1283.465 1459.720 1300.420 1459.770 ;
        RECT 1283.465 1459.470 1304.000 1459.720 ;
        RECT 1283.465 1459.455 1283.795 1459.470 ;
        RECT 1300.000 1459.120 1304.000 1459.470 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 165.210 1490.800 165.530 1490.860 ;
        RECT 1283.470 1490.800 1283.790 1490.860 ;
        RECT 165.210 1490.660 1283.790 1490.800 ;
        RECT 165.210 1490.600 165.530 1490.660 ;
        RECT 1283.470 1490.600 1283.790 1490.660 ;
      LAYER via ;
        RECT 165.240 1490.600 165.500 1490.860 ;
        RECT 1283.500 1490.600 1283.760 1490.860 ;
      LAYER met2 ;
        RECT 1283.490 1491.395 1283.770 1491.765 ;
        RECT 1283.560 1490.890 1283.700 1491.395 ;
        RECT 165.240 1490.570 165.500 1490.890 ;
        RECT 1283.500 1490.570 1283.760 1490.890 ;
        RECT 165.300 17.410 165.440 1490.570 ;
        RECT 163.460 17.270 165.440 17.410 ;
        RECT 163.460 2.400 163.600 17.270 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1491.440 1283.770 1491.720 ;
      LAYER met3 ;
        RECT 1283.465 1491.730 1283.795 1491.745 ;
        RECT 1283.465 1491.680 1300.420 1491.730 ;
        RECT 1283.465 1491.430 1304.000 1491.680 ;
        RECT 1283.465 1491.415 1283.795 1491.430 ;
        RECT 1300.000 1491.080 1304.000 1491.430 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 185.910 1518.340 186.230 1518.400 ;
        RECT 1283.470 1518.340 1283.790 1518.400 ;
        RECT 185.910 1518.200 1283.790 1518.340 ;
        RECT 185.910 1518.140 186.230 1518.200 ;
        RECT 1283.470 1518.140 1283.790 1518.200 ;
        RECT 180.850 17.920 181.170 17.980 ;
        RECT 185.910 17.920 186.230 17.980 ;
        RECT 180.850 17.780 186.230 17.920 ;
        RECT 180.850 17.720 181.170 17.780 ;
        RECT 185.910 17.720 186.230 17.780 ;
      LAYER via ;
        RECT 185.940 1518.140 186.200 1518.400 ;
        RECT 1283.500 1518.140 1283.760 1518.400 ;
        RECT 180.880 17.720 181.140 17.980 ;
        RECT 185.940 17.720 186.200 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1523.355 1283.770 1523.725 ;
        RECT 1283.560 1518.430 1283.700 1523.355 ;
        RECT 185.940 1518.110 186.200 1518.430 ;
        RECT 1283.500 1518.110 1283.760 1518.430 ;
        RECT 186.000 18.010 186.140 1518.110 ;
        RECT 180.880 17.690 181.140 18.010 ;
        RECT 185.940 17.690 186.200 18.010 ;
        RECT 180.940 2.400 181.080 17.690 ;
        RECT 180.730 -4.800 181.290 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1523.400 1283.770 1523.680 ;
      LAYER met3 ;
        RECT 1283.465 1523.690 1283.795 1523.705 ;
        RECT 1283.465 1523.640 1300.420 1523.690 ;
        RECT 1283.465 1523.390 1304.000 1523.640 ;
        RECT 1283.465 1523.375 1283.795 1523.390 ;
        RECT 1300.000 1523.040 1304.000 1523.390 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 199.710 1552.680 200.030 1552.740 ;
        RECT 1283.470 1552.680 1283.790 1552.740 ;
        RECT 199.710 1552.540 1283.790 1552.680 ;
        RECT 199.710 1552.480 200.030 1552.540 ;
        RECT 1283.470 1552.480 1283.790 1552.540 ;
      LAYER via ;
        RECT 199.740 1552.480 200.000 1552.740 ;
        RECT 1283.500 1552.480 1283.760 1552.740 ;
      LAYER met2 ;
        RECT 1283.490 1555.315 1283.770 1555.685 ;
        RECT 1283.560 1552.770 1283.700 1555.315 ;
        RECT 199.740 1552.450 200.000 1552.770 ;
        RECT 1283.500 1552.450 1283.760 1552.770 ;
        RECT 199.800 17.410 199.940 1552.450 ;
        RECT 198.880 17.270 199.940 17.410 ;
        RECT 198.880 2.400 199.020 17.270 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1555.360 1283.770 1555.640 ;
      LAYER met3 ;
        RECT 1283.465 1555.650 1283.795 1555.665 ;
        RECT 1283.465 1555.600 1300.420 1555.650 ;
        RECT 1283.465 1555.350 1304.000 1555.600 ;
        RECT 1283.465 1555.335 1283.795 1555.350 ;
        RECT 1300.000 1555.000 1304.000 1555.350 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 220.410 1587.360 220.730 1587.420 ;
        RECT 1283.470 1587.360 1283.790 1587.420 ;
        RECT 220.410 1587.220 1283.790 1587.360 ;
        RECT 220.410 1587.160 220.730 1587.220 ;
        RECT 1283.470 1587.160 1283.790 1587.220 ;
        RECT 216.730 17.920 217.050 17.980 ;
        RECT 220.410 17.920 220.730 17.980 ;
        RECT 216.730 17.780 220.730 17.920 ;
        RECT 216.730 17.720 217.050 17.780 ;
        RECT 220.410 17.720 220.730 17.780 ;
      LAYER via ;
        RECT 220.440 1587.160 220.700 1587.420 ;
        RECT 1283.500 1587.160 1283.760 1587.420 ;
        RECT 216.760 17.720 217.020 17.980 ;
        RECT 220.440 17.720 220.700 17.980 ;
      LAYER met2 ;
        RECT 220.440 1587.130 220.700 1587.450 ;
        RECT 1283.490 1587.275 1283.770 1587.645 ;
        RECT 1283.500 1587.130 1283.760 1587.275 ;
        RECT 220.500 18.010 220.640 1587.130 ;
        RECT 216.760 17.690 217.020 18.010 ;
        RECT 220.440 17.690 220.700 18.010 ;
        RECT 216.820 2.400 216.960 17.690 ;
        RECT 216.610 -4.800 217.170 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1587.320 1283.770 1587.600 ;
      LAYER met3 ;
        RECT 1283.465 1587.610 1283.795 1587.625 ;
        RECT 1283.465 1587.560 1300.420 1587.610 ;
        RECT 1283.465 1587.310 1304.000 1587.560 ;
        RECT 1283.465 1587.295 1283.795 1587.310 ;
        RECT 1300.000 1586.960 1304.000 1587.310 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 240.650 1614.900 240.970 1614.960 ;
        RECT 1283.470 1614.900 1283.790 1614.960 ;
        RECT 240.650 1614.760 1283.790 1614.900 ;
        RECT 240.650 1614.700 240.970 1614.760 ;
        RECT 1283.470 1614.700 1283.790 1614.760 ;
        RECT 234.670 17.920 234.990 17.980 ;
        RECT 240.650 17.920 240.970 17.980 ;
        RECT 234.670 17.780 240.970 17.920 ;
        RECT 234.670 17.720 234.990 17.780 ;
        RECT 240.650 17.720 240.970 17.780 ;
      LAYER via ;
        RECT 240.680 1614.700 240.940 1614.960 ;
        RECT 1283.500 1614.700 1283.760 1614.960 ;
        RECT 234.700 17.720 234.960 17.980 ;
        RECT 240.680 17.720 240.940 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1619.235 1283.770 1619.605 ;
        RECT 1283.560 1614.990 1283.700 1619.235 ;
        RECT 240.680 1614.670 240.940 1614.990 ;
        RECT 1283.500 1614.670 1283.760 1614.990 ;
        RECT 240.740 468.930 240.880 1614.670 ;
        RECT 240.280 468.790 240.880 468.930 ;
        RECT 240.280 434.930 240.420 468.790 ;
        RECT 240.280 434.790 240.880 434.930 ;
        RECT 240.740 18.010 240.880 434.790 ;
        RECT 234.700 17.690 234.960 18.010 ;
        RECT 240.680 17.690 240.940 18.010 ;
        RECT 234.760 2.400 234.900 17.690 ;
        RECT 234.550 -4.800 235.110 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1619.280 1283.770 1619.560 ;
      LAYER met3 ;
        RECT 1283.465 1619.570 1283.795 1619.585 ;
        RECT 1283.465 1619.520 1300.420 1619.570 ;
        RECT 1283.465 1619.270 1304.000 1619.520 ;
        RECT 1283.465 1619.255 1283.795 1619.270 ;
        RECT 1300.000 1618.920 1304.000 1619.270 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 61.710 1297.340 62.030 1297.400 ;
        RECT 1283.470 1297.340 1283.790 1297.400 ;
        RECT 61.710 1297.200 1283.790 1297.340 ;
        RECT 61.710 1297.140 62.030 1297.200 ;
        RECT 1283.470 1297.140 1283.790 1297.200 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 61.710 17.920 62.030 17.980 ;
        RECT 56.190 17.780 62.030 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 61.710 17.720 62.030 17.780 ;
      LAYER via ;
        RECT 61.740 1297.140 62.000 1297.400 ;
        RECT 1283.500 1297.140 1283.760 1297.400 ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 61.740 17.720 62.000 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1300.315 1283.770 1300.685 ;
        RECT 1283.560 1297.430 1283.700 1300.315 ;
        RECT 61.740 1297.110 62.000 1297.430 ;
        RECT 1283.500 1297.110 1283.760 1297.430 ;
        RECT 61.800 18.010 61.940 1297.110 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 61.740 17.690 62.000 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1300.360 1283.770 1300.640 ;
      LAYER met3 ;
        RECT 1283.465 1300.650 1283.795 1300.665 ;
        RECT 1283.465 1300.600 1300.420 1300.650 ;
        RECT 1283.465 1300.350 1304.000 1300.600 ;
        RECT 1283.465 1300.335 1283.795 1300.350 ;
        RECT 1300.000 1300.000 1304.000 1300.350 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 82.410 1338.820 82.730 1338.880 ;
        RECT 1283.470 1338.820 1283.790 1338.880 ;
        RECT 82.410 1338.680 1283.790 1338.820 ;
        RECT 82.410 1338.620 82.730 1338.680 ;
        RECT 1283.470 1338.620 1283.790 1338.680 ;
        RECT 80.110 17.920 80.430 17.980 ;
        RECT 82.410 17.920 82.730 17.980 ;
        RECT 80.110 17.780 82.730 17.920 ;
        RECT 80.110 17.720 80.430 17.780 ;
        RECT 82.410 17.720 82.730 17.780 ;
      LAYER via ;
        RECT 82.440 1338.620 82.700 1338.880 ;
        RECT 1283.500 1338.620 1283.760 1338.880 ;
        RECT 80.140 17.720 80.400 17.980 ;
        RECT 82.440 17.720 82.700 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1343.155 1283.770 1343.525 ;
        RECT 1283.560 1338.910 1283.700 1343.155 ;
        RECT 82.440 1338.590 82.700 1338.910 ;
        RECT 1283.500 1338.590 1283.760 1338.910 ;
        RECT 82.500 18.010 82.640 1338.590 ;
        RECT 80.140 17.690 80.400 18.010 ;
        RECT 82.440 17.690 82.700 18.010 ;
        RECT 80.200 2.400 80.340 17.690 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1343.200 1283.770 1343.480 ;
      LAYER met3 ;
        RECT 1283.465 1343.490 1283.795 1343.505 ;
        RECT 1283.465 1343.440 1300.420 1343.490 ;
        RECT 1283.465 1343.190 1304.000 1343.440 ;
        RECT 1283.465 1343.175 1283.795 1343.190 ;
        RECT 1300.000 1342.840 1304.000 1343.190 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 1380.300 109.870 1380.360 ;
        RECT 1283.470 1380.300 1283.790 1380.360 ;
        RECT 109.550 1380.160 1283.790 1380.300 ;
        RECT 109.550 1380.100 109.870 1380.160 ;
        RECT 1283.470 1380.100 1283.790 1380.160 ;
        RECT 103.570 17.920 103.890 17.980 ;
        RECT 109.550 17.920 109.870 17.980 ;
        RECT 103.570 17.780 109.870 17.920 ;
        RECT 103.570 17.720 103.890 17.780 ;
        RECT 109.550 17.720 109.870 17.780 ;
      LAYER via ;
        RECT 109.580 1380.100 109.840 1380.360 ;
        RECT 1283.500 1380.100 1283.760 1380.360 ;
        RECT 103.600 17.720 103.860 17.980 ;
        RECT 109.580 17.720 109.840 17.980 ;
      LAYER met2 ;
        RECT 1283.490 1385.315 1283.770 1385.685 ;
        RECT 1283.560 1380.390 1283.700 1385.315 ;
        RECT 109.580 1380.070 109.840 1380.390 ;
        RECT 1283.500 1380.070 1283.760 1380.390 ;
        RECT 109.640 18.010 109.780 1380.070 ;
        RECT 103.600 17.690 103.860 18.010 ;
        RECT 109.580 17.690 109.840 18.010 ;
        RECT 103.660 2.400 103.800 17.690 ;
        RECT 103.450 -4.800 104.010 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1385.360 1283.770 1385.640 ;
      LAYER met3 ;
        RECT 1283.465 1385.650 1283.795 1385.665 ;
        RECT 1283.465 1385.600 1300.420 1385.650 ;
        RECT 1283.465 1385.350 1304.000 1385.600 ;
        RECT 1283.465 1385.335 1283.795 1385.350 ;
        RECT 1300.000 1385.000 1304.000 1385.350 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 130.710 1428.580 131.030 1428.640 ;
        RECT 1283.470 1428.580 1283.790 1428.640 ;
        RECT 130.710 1428.440 1283.790 1428.580 ;
        RECT 130.710 1428.380 131.030 1428.440 ;
        RECT 1283.470 1428.380 1283.790 1428.440 ;
        RECT 127.490 17.920 127.810 17.980 ;
        RECT 130.710 17.920 131.030 17.980 ;
        RECT 127.490 17.780 131.030 17.920 ;
        RECT 127.490 17.720 127.810 17.780 ;
        RECT 130.710 17.720 131.030 17.780 ;
      LAYER via ;
        RECT 130.740 1428.380 131.000 1428.640 ;
        RECT 1283.500 1428.380 1283.760 1428.640 ;
        RECT 127.520 17.720 127.780 17.980 ;
        RECT 130.740 17.720 131.000 17.980 ;
      LAYER met2 ;
        RECT 130.740 1428.350 131.000 1428.670 ;
        RECT 1283.500 1428.525 1283.760 1428.670 ;
        RECT 130.800 18.010 130.940 1428.350 ;
        RECT 1283.490 1428.155 1283.770 1428.525 ;
        RECT 127.520 17.690 127.780 18.010 ;
        RECT 130.740 17.690 131.000 18.010 ;
        RECT 127.580 2.400 127.720 17.690 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1428.200 1283.770 1428.480 ;
      LAYER met3 ;
        RECT 1283.465 1428.490 1283.795 1428.505 ;
        RECT 1283.465 1428.440 1300.420 1428.490 ;
        RECT 1283.465 1428.190 1304.000 1428.440 ;
        RECT 1283.465 1428.175 1283.795 1428.190 ;
        RECT 1300.000 1427.840 1304.000 1428.190 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 27.210 1242.260 27.530 1242.320 ;
        RECT 1283.470 1242.260 1283.790 1242.320 ;
        RECT 27.210 1242.120 1283.790 1242.260 ;
        RECT 27.210 1242.060 27.530 1242.120 ;
        RECT 1283.470 1242.060 1283.790 1242.120 ;
        RECT 26.290 2.960 26.610 3.020 ;
        RECT 27.210 2.960 27.530 3.020 ;
        RECT 26.290 2.820 27.530 2.960 ;
        RECT 26.290 2.760 26.610 2.820 ;
        RECT 27.210 2.760 27.530 2.820 ;
      LAYER via ;
        RECT 27.240 1242.060 27.500 1242.320 ;
        RECT 1283.500 1242.060 1283.760 1242.320 ;
        RECT 26.320 2.760 26.580 3.020 ;
        RECT 27.240 2.760 27.500 3.020 ;
      LAYER met2 ;
        RECT 1283.490 1247.275 1283.770 1247.645 ;
        RECT 1283.560 1242.350 1283.700 1247.275 ;
        RECT 27.240 1242.030 27.500 1242.350 ;
        RECT 1283.500 1242.030 1283.760 1242.350 ;
        RECT 27.300 3.050 27.440 1242.030 ;
        RECT 26.320 2.730 26.580 3.050 ;
        RECT 27.240 2.730 27.500 3.050 ;
        RECT 26.380 2.400 26.520 2.730 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1247.320 1283.770 1247.600 ;
      LAYER met3 ;
        RECT 1283.465 1247.610 1283.795 1247.625 ;
        RECT 1283.465 1247.560 1300.420 1247.610 ;
        RECT 1283.465 1247.310 1304.000 1247.560 ;
        RECT 1283.465 1247.295 1283.795 1247.310 ;
        RECT 1300.000 1246.960 1304.000 1247.310 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 34.110 1256.200 34.430 1256.260 ;
        RECT 1283.470 1256.200 1283.790 1256.260 ;
        RECT 34.110 1256.060 1283.790 1256.200 ;
        RECT 34.110 1256.000 34.430 1256.060 ;
        RECT 1283.470 1256.000 1283.790 1256.060 ;
      LAYER via ;
        RECT 34.140 1256.000 34.400 1256.260 ;
        RECT 1283.500 1256.000 1283.760 1256.260 ;
      LAYER met2 ;
        RECT 1283.490 1258.155 1283.770 1258.525 ;
        RECT 1283.560 1256.290 1283.700 1258.155 ;
        RECT 34.140 1255.970 34.400 1256.290 ;
        RECT 1283.500 1255.970 1283.760 1256.290 ;
        RECT 34.200 3.130 34.340 1255.970 ;
        RECT 32.360 2.990 34.340 3.130 ;
        RECT 32.360 2.400 32.500 2.990 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 1283.490 1258.200 1283.770 1258.480 ;
      LAYER met3 ;
        RECT 1283.465 1258.490 1283.795 1258.505 ;
        RECT 1283.465 1258.440 1300.420 1258.490 ;
        RECT 1283.465 1258.190 1304.000 1258.440 ;
        RECT 1283.465 1258.175 1283.795 1258.190 ;
        RECT 1300.000 1257.840 1304.000 1258.190 ;
    END
  END wbs_we_i
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.010 1192.620 1306.330 1192.680 ;
        RECT 1486.790 1192.620 1487.110 1192.680 ;
        RECT 1306.010 1192.480 1487.110 1192.620 ;
        RECT 1306.010 1192.420 1306.330 1192.480 ;
        RECT 1486.790 1192.420 1487.110 1192.480 ;
        RECT 1486.790 1014.120 1487.110 1014.180 ;
        RECT 1489.550 1014.120 1489.870 1014.180 ;
        RECT 1486.790 1013.980 1489.870 1014.120 ;
        RECT 1486.790 1013.920 1487.110 1013.980 ;
        RECT 1489.550 1013.920 1489.870 1013.980 ;
        RECT 1489.550 1007.660 1489.870 1007.720 ;
        RECT 2087.090 1007.660 2087.410 1007.720 ;
        RECT 1489.550 1007.520 2087.410 1007.660 ;
        RECT 1489.550 1007.460 1489.870 1007.520 ;
        RECT 2087.090 1007.460 2087.410 1007.520 ;
        RECT 1489.550 544.580 1489.870 544.640 ;
        RECT 1518.070 544.580 1518.390 544.640 ;
        RECT 1528.190 544.580 1528.510 544.640 ;
        RECT 1538.770 544.580 1539.090 544.640 ;
        RECT 1489.550 544.440 1539.090 544.580 ;
        RECT 1489.550 544.380 1489.870 544.440 ;
        RECT 1518.070 544.380 1518.390 544.440 ;
        RECT 1528.190 544.380 1528.510 544.440 ;
        RECT 1538.770 544.380 1539.090 544.440 ;
        RECT 2090.310 544.580 2090.630 544.640 ;
        RECT 2121.130 544.580 2121.450 544.640 ;
        RECT 2139.070 544.580 2139.390 544.640 ;
        RECT 2090.310 544.440 2139.390 544.580 ;
        RECT 2090.310 544.380 2090.630 544.440 ;
        RECT 2121.130 544.380 2121.450 544.440 ;
        RECT 2139.070 544.380 2139.390 544.440 ;
        RECT 710.310 14.180 710.630 14.240 ;
        RECT 728.250 14.180 728.570 14.240 ;
        RECT 746.190 14.180 746.510 14.240 ;
        RECT 763.670 14.180 763.990 14.240 ;
        RECT 781.610 14.180 781.930 14.240 ;
        RECT 799.550 14.180 799.870 14.240 ;
        RECT 817.490 14.180 817.810 14.240 ;
        RECT 835.430 14.180 835.750 14.240 ;
        RECT 852.910 14.180 853.230 14.240 ;
        RECT 870.850 14.180 871.170 14.240 ;
        RECT 888.790 14.180 889.110 14.240 ;
        RECT 906.730 14.180 907.050 14.240 ;
        RECT 924.210 14.180 924.530 14.240 ;
        RECT 942.150 14.180 942.470 14.240 ;
        RECT 960.090 14.180 960.410 14.240 ;
        RECT 978.030 14.180 978.350 14.240 ;
        RECT 995.970 14.180 996.290 14.240 ;
        RECT 1013.450 14.180 1013.770 14.240 ;
        RECT 1031.390 14.180 1031.710 14.240 ;
        RECT 1049.330 14.180 1049.650 14.240 ;
        RECT 1067.270 14.180 1067.590 14.240 ;
        RECT 1085.210 14.180 1085.530 14.240 ;
        RECT 1102.690 14.180 1103.010 14.240 ;
        RECT 1120.630 14.180 1120.950 14.240 ;
        RECT 1138.570 14.180 1138.890 14.240 ;
        RECT 1156.510 14.180 1156.830 14.240 ;
        RECT 1173.990 14.180 1174.310 14.240 ;
        RECT 1191.930 14.180 1192.250 14.240 ;
        RECT 1209.870 14.180 1210.190 14.240 ;
        RECT 1227.810 14.180 1228.130 14.240 ;
        RECT 1245.750 14.180 1246.070 14.240 ;
        RECT 1263.230 14.180 1263.550 14.240 ;
        RECT 1281.170 14.180 1281.490 14.240 ;
        RECT 1299.110 14.180 1299.430 14.240 ;
        RECT 1317.050 14.180 1317.370 14.240 ;
        RECT 1334.990 14.180 1335.310 14.240 ;
        RECT 1352.470 14.180 1352.790 14.240 ;
        RECT 1370.410 14.180 1370.730 14.240 ;
        RECT 1388.350 14.180 1388.670 14.240 ;
        RECT 1406.290 14.180 1406.610 14.240 ;
        RECT 1423.770 14.180 1424.090 14.240 ;
        RECT 1441.710 14.180 1442.030 14.240 ;
        RECT 1459.650 14.180 1459.970 14.240 ;
        RECT 1477.590 14.180 1477.910 14.240 ;
        RECT 1495.530 14.180 1495.850 14.240 ;
        RECT 1513.010 14.180 1513.330 14.240 ;
        RECT 1528.190 14.180 1528.510 14.240 ;
        RECT 1530.950 14.180 1531.270 14.240 ;
        RECT 1548.890 14.180 1549.210 14.240 ;
        RECT 1566.830 14.180 1567.150 14.240 ;
        RECT 1584.770 14.180 1585.090 14.240 ;
        RECT 1602.250 14.180 1602.570 14.240 ;
        RECT 1620.190 14.180 1620.510 14.240 ;
        RECT 1638.130 14.180 1638.450 14.240 ;
        RECT 1656.070 14.180 1656.390 14.240 ;
        RECT 1673.550 14.180 1673.870 14.240 ;
        RECT 1691.490 14.180 1691.810 14.240 ;
        RECT 1709.430 14.180 1709.750 14.240 ;
        RECT 1727.370 14.180 1727.690 14.240 ;
        RECT 1745.310 14.180 1745.630 14.240 ;
        RECT 1762.790 14.180 1763.110 14.240 ;
        RECT 1780.730 14.180 1781.050 14.240 ;
        RECT 1798.670 14.180 1798.990 14.240 ;
        RECT 1816.610 14.180 1816.930 14.240 ;
        RECT 1834.550 14.180 1834.870 14.240 ;
        RECT 1852.030 14.180 1852.350 14.240 ;
        RECT 1869.970 14.180 1870.290 14.240 ;
        RECT 1887.910 14.180 1888.230 14.240 ;
        RECT 1905.850 14.180 1906.170 14.240 ;
        RECT 1923.330 14.180 1923.650 14.240 ;
        RECT 1941.270 14.180 1941.590 14.240 ;
        RECT 1959.210 14.180 1959.530 14.240 ;
        RECT 1977.150 14.180 1977.470 14.240 ;
        RECT 1995.090 14.180 1995.410 14.240 ;
        RECT 2012.570 14.180 2012.890 14.240 ;
        RECT 2030.510 14.180 2030.830 14.240 ;
        RECT 2048.450 14.180 2048.770 14.240 ;
        RECT 2066.390 14.180 2066.710 14.240 ;
        RECT 2084.330 14.180 2084.650 14.240 ;
        RECT 2101.810 14.180 2102.130 14.240 ;
        RECT 2119.750 14.180 2120.070 14.240 ;
        RECT 2137.690 14.180 2138.010 14.240 ;
        RECT 2155.630 14.180 2155.950 14.240 ;
        RECT 2173.110 14.180 2173.430 14.240 ;
        RECT 2191.050 14.180 2191.370 14.240 ;
        RECT 2208.990 14.180 2209.310 14.240 ;
        RECT 2226.930 14.180 2227.250 14.240 ;
        RECT 2244.870 14.180 2245.190 14.240 ;
        RECT 2262.350 14.180 2262.670 14.240 ;
        RECT 2280.290 14.180 2280.610 14.240 ;
        RECT 2298.230 14.180 2298.550 14.240 ;
        RECT 2316.170 14.180 2316.490 14.240 ;
        RECT 2334.110 14.180 2334.430 14.240 ;
        RECT 2351.590 14.180 2351.910 14.240 ;
        RECT 2369.530 14.180 2369.850 14.240 ;
        RECT 2387.470 14.180 2387.790 14.240 ;
        RECT 2405.410 14.180 2405.730 14.240 ;
        RECT 2422.890 14.180 2423.210 14.240 ;
        RECT 2440.830 14.180 2441.150 14.240 ;
        RECT 2458.770 14.180 2459.090 14.240 ;
        RECT 2476.710 14.180 2477.030 14.240 ;
        RECT 2494.650 14.180 2494.970 14.240 ;
        RECT 2512.130 14.180 2512.450 14.240 ;
        RECT 2530.070 14.180 2530.390 14.240 ;
        RECT 2548.010 14.180 2548.330 14.240 ;
        RECT 2565.950 14.180 2566.270 14.240 ;
        RECT 2583.890 14.180 2584.210 14.240 ;
        RECT 2601.370 14.180 2601.690 14.240 ;
        RECT 2619.310 14.180 2619.630 14.240 ;
        RECT 2637.250 14.180 2637.570 14.240 ;
        RECT 2655.190 14.180 2655.510 14.240 ;
        RECT 2672.670 14.180 2672.990 14.240 ;
        RECT 2690.610 14.180 2690.930 14.240 ;
        RECT 2708.550 14.180 2708.870 14.240 ;
        RECT 2726.490 14.180 2726.810 14.240 ;
        RECT 2744.430 14.180 2744.750 14.240 ;
        RECT 2761.910 14.180 2762.230 14.240 ;
        RECT 2779.850 14.180 2780.170 14.240 ;
        RECT 2797.790 14.180 2798.110 14.240 ;
        RECT 2815.730 14.180 2816.050 14.240 ;
        RECT 2833.670 14.180 2833.990 14.240 ;
        RECT 2851.150 14.180 2851.470 14.240 ;
        RECT 2869.090 14.180 2869.410 14.240 ;
        RECT 2887.030 14.180 2887.350 14.240 ;
        RECT 2904.970 14.180 2905.290 14.240 ;
        RECT 710.310 14.040 2905.290 14.180 ;
        RECT 710.310 13.980 710.630 14.040 ;
        RECT 728.250 13.980 728.570 14.040 ;
        RECT 746.190 13.980 746.510 14.040 ;
        RECT 763.670 13.980 763.990 14.040 ;
        RECT 781.610 13.980 781.930 14.040 ;
        RECT 799.550 13.980 799.870 14.040 ;
        RECT 817.490 13.980 817.810 14.040 ;
        RECT 835.430 13.980 835.750 14.040 ;
        RECT 852.910 13.980 853.230 14.040 ;
        RECT 870.850 13.980 871.170 14.040 ;
        RECT 888.790 13.980 889.110 14.040 ;
        RECT 906.730 13.980 907.050 14.040 ;
        RECT 924.210 13.980 924.530 14.040 ;
        RECT 942.150 13.980 942.470 14.040 ;
        RECT 960.090 13.980 960.410 14.040 ;
        RECT 978.030 13.980 978.350 14.040 ;
        RECT 995.970 13.980 996.290 14.040 ;
        RECT 1013.450 13.980 1013.770 14.040 ;
        RECT 1031.390 13.980 1031.710 14.040 ;
        RECT 1049.330 13.980 1049.650 14.040 ;
        RECT 1067.270 13.980 1067.590 14.040 ;
        RECT 1085.210 13.980 1085.530 14.040 ;
        RECT 1102.690 13.980 1103.010 14.040 ;
        RECT 1120.630 13.980 1120.950 14.040 ;
        RECT 1138.570 13.980 1138.890 14.040 ;
        RECT 1156.510 13.980 1156.830 14.040 ;
        RECT 1173.990 13.980 1174.310 14.040 ;
        RECT 1191.930 13.980 1192.250 14.040 ;
        RECT 1209.870 13.980 1210.190 14.040 ;
        RECT 1227.810 13.980 1228.130 14.040 ;
        RECT 1245.750 13.980 1246.070 14.040 ;
        RECT 1263.230 13.980 1263.550 14.040 ;
        RECT 1281.170 13.980 1281.490 14.040 ;
        RECT 1299.110 13.980 1299.430 14.040 ;
        RECT 1317.050 13.980 1317.370 14.040 ;
        RECT 1334.990 13.980 1335.310 14.040 ;
        RECT 1352.470 13.980 1352.790 14.040 ;
        RECT 1370.410 13.980 1370.730 14.040 ;
        RECT 1388.350 13.980 1388.670 14.040 ;
        RECT 1406.290 13.980 1406.610 14.040 ;
        RECT 1423.770 13.980 1424.090 14.040 ;
        RECT 1441.710 13.980 1442.030 14.040 ;
        RECT 1459.650 13.980 1459.970 14.040 ;
        RECT 1477.590 13.980 1477.910 14.040 ;
        RECT 1495.530 13.980 1495.850 14.040 ;
        RECT 1513.010 13.980 1513.330 14.040 ;
        RECT 1528.190 13.980 1528.510 14.040 ;
        RECT 1530.950 13.980 1531.270 14.040 ;
        RECT 1548.890 13.980 1549.210 14.040 ;
        RECT 1566.830 13.980 1567.150 14.040 ;
        RECT 1584.770 13.980 1585.090 14.040 ;
        RECT 1602.250 13.980 1602.570 14.040 ;
        RECT 1620.190 13.980 1620.510 14.040 ;
        RECT 1638.130 13.980 1638.450 14.040 ;
        RECT 1656.070 13.980 1656.390 14.040 ;
        RECT 1673.550 13.980 1673.870 14.040 ;
        RECT 1691.490 13.980 1691.810 14.040 ;
        RECT 1709.430 13.980 1709.750 14.040 ;
        RECT 1727.370 13.980 1727.690 14.040 ;
        RECT 1745.310 13.980 1745.630 14.040 ;
        RECT 1762.790 13.980 1763.110 14.040 ;
        RECT 1780.730 13.980 1781.050 14.040 ;
        RECT 1798.670 13.980 1798.990 14.040 ;
        RECT 1816.610 13.980 1816.930 14.040 ;
        RECT 1834.550 13.980 1834.870 14.040 ;
        RECT 1852.030 13.980 1852.350 14.040 ;
        RECT 1869.970 13.980 1870.290 14.040 ;
        RECT 1887.910 13.980 1888.230 14.040 ;
        RECT 1905.850 13.980 1906.170 14.040 ;
        RECT 1923.330 13.980 1923.650 14.040 ;
        RECT 1941.270 13.980 1941.590 14.040 ;
        RECT 1959.210 13.980 1959.530 14.040 ;
        RECT 1977.150 13.980 1977.470 14.040 ;
        RECT 1995.090 13.980 1995.410 14.040 ;
        RECT 2012.570 13.980 2012.890 14.040 ;
        RECT 2030.510 13.980 2030.830 14.040 ;
        RECT 2048.450 13.980 2048.770 14.040 ;
        RECT 2066.390 13.980 2066.710 14.040 ;
        RECT 2084.330 13.980 2084.650 14.040 ;
        RECT 2101.810 13.980 2102.130 14.040 ;
        RECT 2119.750 13.980 2120.070 14.040 ;
        RECT 2137.690 13.980 2138.010 14.040 ;
        RECT 2155.630 13.980 2155.950 14.040 ;
        RECT 2173.110 13.980 2173.430 14.040 ;
        RECT 2191.050 13.980 2191.370 14.040 ;
        RECT 2208.990 13.980 2209.310 14.040 ;
        RECT 2226.930 13.980 2227.250 14.040 ;
        RECT 2244.870 13.980 2245.190 14.040 ;
        RECT 2262.350 13.980 2262.670 14.040 ;
        RECT 2280.290 13.980 2280.610 14.040 ;
        RECT 2298.230 13.980 2298.550 14.040 ;
        RECT 2316.170 13.980 2316.490 14.040 ;
        RECT 2334.110 13.980 2334.430 14.040 ;
        RECT 2351.590 13.980 2351.910 14.040 ;
        RECT 2369.530 13.980 2369.850 14.040 ;
        RECT 2387.470 13.980 2387.790 14.040 ;
        RECT 2405.410 13.980 2405.730 14.040 ;
        RECT 2422.890 13.980 2423.210 14.040 ;
        RECT 2440.830 13.980 2441.150 14.040 ;
        RECT 2458.770 13.980 2459.090 14.040 ;
        RECT 2476.710 13.980 2477.030 14.040 ;
        RECT 2494.650 13.980 2494.970 14.040 ;
        RECT 2512.130 13.980 2512.450 14.040 ;
        RECT 2530.070 13.980 2530.390 14.040 ;
        RECT 2548.010 13.980 2548.330 14.040 ;
        RECT 2565.950 13.980 2566.270 14.040 ;
        RECT 2583.890 13.980 2584.210 14.040 ;
        RECT 2601.370 13.980 2601.690 14.040 ;
        RECT 2619.310 13.980 2619.630 14.040 ;
        RECT 2637.250 13.980 2637.570 14.040 ;
        RECT 2655.190 13.980 2655.510 14.040 ;
        RECT 2672.670 13.980 2672.990 14.040 ;
        RECT 2690.610 13.980 2690.930 14.040 ;
        RECT 2708.550 13.980 2708.870 14.040 ;
        RECT 2726.490 13.980 2726.810 14.040 ;
        RECT 2744.430 13.980 2744.750 14.040 ;
        RECT 2761.910 13.980 2762.230 14.040 ;
        RECT 2779.850 13.980 2780.170 14.040 ;
        RECT 2797.790 13.980 2798.110 14.040 ;
        RECT 2815.730 13.980 2816.050 14.040 ;
        RECT 2833.670 13.980 2833.990 14.040 ;
        RECT 2851.150 13.980 2851.470 14.040 ;
        RECT 2869.090 13.980 2869.410 14.040 ;
        RECT 2887.030 13.980 2887.350 14.040 ;
        RECT 2904.970 13.980 2905.290 14.040 ;
        RECT 692.370 2.960 692.690 3.020 ;
        RECT 710.310 2.960 710.630 3.020 ;
        RECT 692.370 2.820 710.630 2.960 ;
        RECT 692.370 2.760 692.690 2.820 ;
        RECT 710.310 2.760 710.630 2.820 ;
      LAYER via ;
        RECT 1306.040 1192.420 1306.300 1192.680 ;
        RECT 1486.820 1192.420 1487.080 1192.680 ;
        RECT 1486.820 1013.920 1487.080 1014.180 ;
        RECT 1489.580 1013.920 1489.840 1014.180 ;
        RECT 1489.580 1007.460 1489.840 1007.720 ;
        RECT 2087.120 1007.460 2087.380 1007.720 ;
        RECT 1489.580 544.380 1489.840 544.640 ;
        RECT 1518.100 544.380 1518.360 544.640 ;
        RECT 1528.220 544.380 1528.480 544.640 ;
        RECT 1538.800 544.380 1539.060 544.640 ;
        RECT 2090.340 544.380 2090.600 544.640 ;
        RECT 2121.160 544.380 2121.420 544.640 ;
        RECT 2139.100 544.380 2139.360 544.640 ;
        RECT 710.340 13.980 710.600 14.240 ;
        RECT 728.280 13.980 728.540 14.240 ;
        RECT 746.220 13.980 746.480 14.240 ;
        RECT 763.700 13.980 763.960 14.240 ;
        RECT 781.640 13.980 781.900 14.240 ;
        RECT 799.580 13.980 799.840 14.240 ;
        RECT 817.520 13.980 817.780 14.240 ;
        RECT 835.460 13.980 835.720 14.240 ;
        RECT 852.940 13.980 853.200 14.240 ;
        RECT 870.880 13.980 871.140 14.240 ;
        RECT 888.820 13.980 889.080 14.240 ;
        RECT 906.760 13.980 907.020 14.240 ;
        RECT 924.240 13.980 924.500 14.240 ;
        RECT 942.180 13.980 942.440 14.240 ;
        RECT 960.120 13.980 960.380 14.240 ;
        RECT 978.060 13.980 978.320 14.240 ;
        RECT 996.000 13.980 996.260 14.240 ;
        RECT 1013.480 13.980 1013.740 14.240 ;
        RECT 1031.420 13.980 1031.680 14.240 ;
        RECT 1049.360 13.980 1049.620 14.240 ;
        RECT 1067.300 13.980 1067.560 14.240 ;
        RECT 1085.240 13.980 1085.500 14.240 ;
        RECT 1102.720 13.980 1102.980 14.240 ;
        RECT 1120.660 13.980 1120.920 14.240 ;
        RECT 1138.600 13.980 1138.860 14.240 ;
        RECT 1156.540 13.980 1156.800 14.240 ;
        RECT 1174.020 13.980 1174.280 14.240 ;
        RECT 1191.960 13.980 1192.220 14.240 ;
        RECT 1209.900 13.980 1210.160 14.240 ;
        RECT 1227.840 13.980 1228.100 14.240 ;
        RECT 1245.780 13.980 1246.040 14.240 ;
        RECT 1263.260 13.980 1263.520 14.240 ;
        RECT 1281.200 13.980 1281.460 14.240 ;
        RECT 1299.140 13.980 1299.400 14.240 ;
        RECT 1317.080 13.980 1317.340 14.240 ;
        RECT 1335.020 13.980 1335.280 14.240 ;
        RECT 1352.500 13.980 1352.760 14.240 ;
        RECT 1370.440 13.980 1370.700 14.240 ;
        RECT 1388.380 13.980 1388.640 14.240 ;
        RECT 1406.320 13.980 1406.580 14.240 ;
        RECT 1423.800 13.980 1424.060 14.240 ;
        RECT 1441.740 13.980 1442.000 14.240 ;
        RECT 1459.680 13.980 1459.940 14.240 ;
        RECT 1477.620 13.980 1477.880 14.240 ;
        RECT 1495.560 13.980 1495.820 14.240 ;
        RECT 1513.040 13.980 1513.300 14.240 ;
        RECT 1528.220 13.980 1528.480 14.240 ;
        RECT 1530.980 13.980 1531.240 14.240 ;
        RECT 1548.920 13.980 1549.180 14.240 ;
        RECT 1566.860 13.980 1567.120 14.240 ;
        RECT 1584.800 13.980 1585.060 14.240 ;
        RECT 1602.280 13.980 1602.540 14.240 ;
        RECT 1620.220 13.980 1620.480 14.240 ;
        RECT 1638.160 13.980 1638.420 14.240 ;
        RECT 1656.100 13.980 1656.360 14.240 ;
        RECT 1673.580 13.980 1673.840 14.240 ;
        RECT 1691.520 13.980 1691.780 14.240 ;
        RECT 1709.460 13.980 1709.720 14.240 ;
        RECT 1727.400 13.980 1727.660 14.240 ;
        RECT 1745.340 13.980 1745.600 14.240 ;
        RECT 1762.820 13.980 1763.080 14.240 ;
        RECT 1780.760 13.980 1781.020 14.240 ;
        RECT 1798.700 13.980 1798.960 14.240 ;
        RECT 1816.640 13.980 1816.900 14.240 ;
        RECT 1834.580 13.980 1834.840 14.240 ;
        RECT 1852.060 13.980 1852.320 14.240 ;
        RECT 1870.000 13.980 1870.260 14.240 ;
        RECT 1887.940 13.980 1888.200 14.240 ;
        RECT 1905.880 13.980 1906.140 14.240 ;
        RECT 1923.360 13.980 1923.620 14.240 ;
        RECT 1941.300 13.980 1941.560 14.240 ;
        RECT 1959.240 13.980 1959.500 14.240 ;
        RECT 1977.180 13.980 1977.440 14.240 ;
        RECT 1995.120 13.980 1995.380 14.240 ;
        RECT 2012.600 13.980 2012.860 14.240 ;
        RECT 2030.540 13.980 2030.800 14.240 ;
        RECT 2048.480 13.980 2048.740 14.240 ;
        RECT 2066.420 13.980 2066.680 14.240 ;
        RECT 2084.360 13.980 2084.620 14.240 ;
        RECT 2101.840 13.980 2102.100 14.240 ;
        RECT 2119.780 13.980 2120.040 14.240 ;
        RECT 2137.720 13.980 2137.980 14.240 ;
        RECT 2155.660 13.980 2155.920 14.240 ;
        RECT 2173.140 13.980 2173.400 14.240 ;
        RECT 2191.080 13.980 2191.340 14.240 ;
        RECT 2209.020 13.980 2209.280 14.240 ;
        RECT 2226.960 13.980 2227.220 14.240 ;
        RECT 2244.900 13.980 2245.160 14.240 ;
        RECT 2262.380 13.980 2262.640 14.240 ;
        RECT 2280.320 13.980 2280.580 14.240 ;
        RECT 2298.260 13.980 2298.520 14.240 ;
        RECT 2316.200 13.980 2316.460 14.240 ;
        RECT 2334.140 13.980 2334.400 14.240 ;
        RECT 2351.620 13.980 2351.880 14.240 ;
        RECT 2369.560 13.980 2369.820 14.240 ;
        RECT 2387.500 13.980 2387.760 14.240 ;
        RECT 2405.440 13.980 2405.700 14.240 ;
        RECT 2422.920 13.980 2423.180 14.240 ;
        RECT 2440.860 13.980 2441.120 14.240 ;
        RECT 2458.800 13.980 2459.060 14.240 ;
        RECT 2476.740 13.980 2477.000 14.240 ;
        RECT 2494.680 13.980 2494.940 14.240 ;
        RECT 2512.160 13.980 2512.420 14.240 ;
        RECT 2530.100 13.980 2530.360 14.240 ;
        RECT 2548.040 13.980 2548.300 14.240 ;
        RECT 2565.980 13.980 2566.240 14.240 ;
        RECT 2583.920 13.980 2584.180 14.240 ;
        RECT 2601.400 13.980 2601.660 14.240 ;
        RECT 2619.340 13.980 2619.600 14.240 ;
        RECT 2637.280 13.980 2637.540 14.240 ;
        RECT 2655.220 13.980 2655.480 14.240 ;
        RECT 2672.700 13.980 2672.960 14.240 ;
        RECT 2690.640 13.980 2690.900 14.240 ;
        RECT 2708.580 13.980 2708.840 14.240 ;
        RECT 2726.520 13.980 2726.780 14.240 ;
        RECT 2744.460 13.980 2744.720 14.240 ;
        RECT 2761.940 13.980 2762.200 14.240 ;
        RECT 2779.880 13.980 2780.140 14.240 ;
        RECT 2797.820 13.980 2798.080 14.240 ;
        RECT 2815.760 13.980 2816.020 14.240 ;
        RECT 2833.700 13.980 2833.960 14.240 ;
        RECT 2851.180 13.980 2851.440 14.240 ;
        RECT 2869.120 13.980 2869.380 14.240 ;
        RECT 2887.060 13.980 2887.320 14.240 ;
        RECT 2905.000 13.980 2905.260 14.240 ;
        RECT 692.400 2.760 692.660 3.020 ;
        RECT 710.340 2.760 710.600 3.020 ;
      LAYER met2 ;
        RECT 1306.070 1200.000 1306.350 1204.000 ;
        RECT 1306.100 1192.710 1306.240 1200.000 ;
        RECT 1306.040 1192.390 1306.300 1192.710 ;
        RECT 1486.820 1192.390 1487.080 1192.710 ;
        RECT 1486.880 1014.210 1487.020 1192.390 ;
        RECT 1486.820 1013.890 1487.080 1014.210 ;
        RECT 1489.580 1013.890 1489.840 1014.210 ;
        RECT 1489.640 1007.750 1489.780 1013.890 ;
        RECT 1489.580 1007.430 1489.840 1007.750 ;
        RECT 2087.120 1007.430 2087.380 1007.750 ;
        RECT 1489.640 901.525 1489.780 1007.430 ;
        RECT 2087.180 902.885 2087.320 1007.430 ;
        RECT 2087.110 902.515 2087.390 902.885 ;
        RECT 1489.570 901.155 1489.850 901.525 ;
        RECT 1489.570 858.995 1489.850 859.365 ;
        RECT 1489.640 544.670 1489.780 858.995 ;
        RECT 2090.330 858.315 2090.610 858.685 ;
        RECT 1518.090 544.835 1518.370 545.205 ;
        RECT 1538.790 544.835 1539.070 545.205 ;
        RECT 1518.160 544.670 1518.300 544.835 ;
        RECT 1538.860 544.670 1539.000 544.835 ;
        RECT 2090.400 544.670 2090.540 858.315 ;
        RECT 2121.150 544.835 2121.430 545.205 ;
        RECT 2139.090 544.835 2139.370 545.205 ;
        RECT 2121.220 544.670 2121.360 544.835 ;
        RECT 2139.160 544.670 2139.300 544.835 ;
        RECT 1489.580 544.350 1489.840 544.670 ;
        RECT 1518.100 544.350 1518.360 544.670 ;
        RECT 1528.220 544.350 1528.480 544.670 ;
        RECT 1538.800 544.350 1539.060 544.670 ;
        RECT 2090.340 544.350 2090.600 544.670 ;
        RECT 2121.160 544.350 2121.420 544.670 ;
        RECT 2139.100 544.350 2139.360 544.670 ;
        RECT 1528.280 14.270 1528.420 544.350 ;
        RECT 710.340 13.950 710.600 14.270 ;
        RECT 728.280 13.950 728.540 14.270 ;
        RECT 746.220 13.950 746.480 14.270 ;
        RECT 763.700 13.950 763.960 14.270 ;
        RECT 781.640 13.950 781.900 14.270 ;
        RECT 799.580 13.950 799.840 14.270 ;
        RECT 817.520 13.950 817.780 14.270 ;
        RECT 835.460 13.950 835.720 14.270 ;
        RECT 852.940 13.950 853.200 14.270 ;
        RECT 870.880 13.950 871.140 14.270 ;
        RECT 888.820 13.950 889.080 14.270 ;
        RECT 906.760 13.950 907.020 14.270 ;
        RECT 924.240 13.950 924.500 14.270 ;
        RECT 942.180 13.950 942.440 14.270 ;
        RECT 960.120 13.950 960.380 14.270 ;
        RECT 978.060 13.950 978.320 14.270 ;
        RECT 996.000 13.950 996.260 14.270 ;
        RECT 1013.480 13.950 1013.740 14.270 ;
        RECT 1031.420 13.950 1031.680 14.270 ;
        RECT 1049.360 13.950 1049.620 14.270 ;
        RECT 1067.300 13.950 1067.560 14.270 ;
        RECT 1085.240 13.950 1085.500 14.270 ;
        RECT 1102.720 13.950 1102.980 14.270 ;
        RECT 1120.660 13.950 1120.920 14.270 ;
        RECT 1138.600 13.950 1138.860 14.270 ;
        RECT 1156.540 13.950 1156.800 14.270 ;
        RECT 1174.020 13.950 1174.280 14.270 ;
        RECT 1191.960 13.950 1192.220 14.270 ;
        RECT 1209.900 13.950 1210.160 14.270 ;
        RECT 1227.840 13.950 1228.100 14.270 ;
        RECT 1245.780 13.950 1246.040 14.270 ;
        RECT 1263.260 13.950 1263.520 14.270 ;
        RECT 1281.200 13.950 1281.460 14.270 ;
        RECT 1299.140 13.950 1299.400 14.270 ;
        RECT 1317.080 13.950 1317.340 14.270 ;
        RECT 1335.020 13.950 1335.280 14.270 ;
        RECT 1352.500 13.950 1352.760 14.270 ;
        RECT 1370.440 13.950 1370.700 14.270 ;
        RECT 1388.380 13.950 1388.640 14.270 ;
        RECT 1406.320 13.950 1406.580 14.270 ;
        RECT 1423.800 13.950 1424.060 14.270 ;
        RECT 1441.740 13.950 1442.000 14.270 ;
        RECT 1459.680 13.950 1459.940 14.270 ;
        RECT 1477.620 13.950 1477.880 14.270 ;
        RECT 1495.560 13.950 1495.820 14.270 ;
        RECT 1513.040 13.950 1513.300 14.270 ;
        RECT 1528.220 13.950 1528.480 14.270 ;
        RECT 1530.980 13.950 1531.240 14.270 ;
        RECT 1548.920 13.950 1549.180 14.270 ;
        RECT 1566.860 13.950 1567.120 14.270 ;
        RECT 1584.800 13.950 1585.060 14.270 ;
        RECT 1602.280 13.950 1602.540 14.270 ;
        RECT 1620.220 13.950 1620.480 14.270 ;
        RECT 1638.160 13.950 1638.420 14.270 ;
        RECT 1656.100 13.950 1656.360 14.270 ;
        RECT 1673.580 13.950 1673.840 14.270 ;
        RECT 1691.520 13.950 1691.780 14.270 ;
        RECT 1709.460 13.950 1709.720 14.270 ;
        RECT 1727.400 13.950 1727.660 14.270 ;
        RECT 1745.340 13.950 1745.600 14.270 ;
        RECT 1762.820 13.950 1763.080 14.270 ;
        RECT 1780.760 13.950 1781.020 14.270 ;
        RECT 1798.700 13.950 1798.960 14.270 ;
        RECT 1816.640 13.950 1816.900 14.270 ;
        RECT 1834.580 13.950 1834.840 14.270 ;
        RECT 1852.060 13.950 1852.320 14.270 ;
        RECT 1870.000 13.950 1870.260 14.270 ;
        RECT 1887.940 13.950 1888.200 14.270 ;
        RECT 1905.880 13.950 1906.140 14.270 ;
        RECT 1923.360 13.950 1923.620 14.270 ;
        RECT 1941.300 13.950 1941.560 14.270 ;
        RECT 1959.240 13.950 1959.500 14.270 ;
        RECT 1977.180 13.950 1977.440 14.270 ;
        RECT 1995.120 13.950 1995.380 14.270 ;
        RECT 2012.600 13.950 2012.860 14.270 ;
        RECT 2030.540 13.950 2030.800 14.270 ;
        RECT 2048.480 13.950 2048.740 14.270 ;
        RECT 2066.420 13.950 2066.680 14.270 ;
        RECT 2084.360 13.950 2084.620 14.270 ;
        RECT 2101.840 13.950 2102.100 14.270 ;
        RECT 2119.780 13.950 2120.040 14.270 ;
        RECT 2137.720 13.950 2137.980 14.270 ;
        RECT 2155.660 13.950 2155.920 14.270 ;
        RECT 2173.140 13.950 2173.400 14.270 ;
        RECT 2191.080 13.950 2191.340 14.270 ;
        RECT 2209.020 13.950 2209.280 14.270 ;
        RECT 2226.960 13.950 2227.220 14.270 ;
        RECT 2244.900 13.950 2245.160 14.270 ;
        RECT 2262.380 13.950 2262.640 14.270 ;
        RECT 2280.320 13.950 2280.580 14.270 ;
        RECT 2298.260 13.950 2298.520 14.270 ;
        RECT 2316.200 13.950 2316.460 14.270 ;
        RECT 2334.140 13.950 2334.400 14.270 ;
        RECT 2351.620 13.950 2351.880 14.270 ;
        RECT 2369.560 13.950 2369.820 14.270 ;
        RECT 2387.500 13.950 2387.760 14.270 ;
        RECT 2405.440 13.950 2405.700 14.270 ;
        RECT 2422.920 13.950 2423.180 14.270 ;
        RECT 2440.860 13.950 2441.120 14.270 ;
        RECT 2458.800 13.950 2459.060 14.270 ;
        RECT 2476.740 13.950 2477.000 14.270 ;
        RECT 2494.680 13.950 2494.940 14.270 ;
        RECT 2512.160 13.950 2512.420 14.270 ;
        RECT 2530.100 13.950 2530.360 14.270 ;
        RECT 2548.040 13.950 2548.300 14.270 ;
        RECT 2565.980 13.950 2566.240 14.270 ;
        RECT 2583.920 13.950 2584.180 14.270 ;
        RECT 2601.400 13.950 2601.660 14.270 ;
        RECT 2619.340 13.950 2619.600 14.270 ;
        RECT 2637.280 13.950 2637.540 14.270 ;
        RECT 2655.220 13.950 2655.480 14.270 ;
        RECT 2672.700 13.950 2672.960 14.270 ;
        RECT 2690.640 13.950 2690.900 14.270 ;
        RECT 2708.580 13.950 2708.840 14.270 ;
        RECT 2726.520 13.950 2726.780 14.270 ;
        RECT 2744.460 13.950 2744.720 14.270 ;
        RECT 2761.940 13.950 2762.200 14.270 ;
        RECT 2779.880 13.950 2780.140 14.270 ;
        RECT 2797.820 13.950 2798.080 14.270 ;
        RECT 2815.760 13.950 2816.020 14.270 ;
        RECT 2833.700 13.950 2833.960 14.270 ;
        RECT 2851.180 13.950 2851.440 14.270 ;
        RECT 2869.120 13.950 2869.380 14.270 ;
        RECT 2887.060 13.950 2887.320 14.270 ;
        RECT 2905.000 13.950 2905.260 14.270 ;
        RECT 710.400 3.050 710.540 13.950 ;
        RECT 692.400 2.730 692.660 3.050 ;
        RECT 710.340 2.730 710.600 3.050 ;
        RECT 692.460 2.400 692.600 2.730 ;
        RECT 710.400 2.400 710.540 2.730 ;
        RECT 728.340 2.400 728.480 13.950 ;
        RECT 746.280 2.400 746.420 13.950 ;
        RECT 763.760 2.400 763.900 13.950 ;
        RECT 781.700 2.400 781.840 13.950 ;
        RECT 799.640 2.400 799.780 13.950 ;
        RECT 817.580 2.400 817.720 13.950 ;
        RECT 835.520 2.400 835.660 13.950 ;
        RECT 853.000 2.400 853.140 13.950 ;
        RECT 870.940 2.400 871.080 13.950 ;
        RECT 888.880 2.400 889.020 13.950 ;
        RECT 906.820 2.400 906.960 13.950 ;
        RECT 924.300 2.400 924.440 13.950 ;
        RECT 942.240 2.400 942.380 13.950 ;
        RECT 960.180 2.400 960.320 13.950 ;
        RECT 978.120 2.400 978.260 13.950 ;
        RECT 996.060 2.400 996.200 13.950 ;
        RECT 1013.540 2.400 1013.680 13.950 ;
        RECT 1031.480 2.400 1031.620 13.950 ;
        RECT 1049.420 2.400 1049.560 13.950 ;
        RECT 1067.360 2.400 1067.500 13.950 ;
        RECT 1085.300 2.400 1085.440 13.950 ;
        RECT 1102.780 2.400 1102.920 13.950 ;
        RECT 1120.720 2.400 1120.860 13.950 ;
        RECT 1138.660 2.400 1138.800 13.950 ;
        RECT 1156.600 2.400 1156.740 13.950 ;
        RECT 1174.080 2.400 1174.220 13.950 ;
        RECT 1192.020 2.400 1192.160 13.950 ;
        RECT 1209.960 2.400 1210.100 13.950 ;
        RECT 1227.900 2.400 1228.040 13.950 ;
        RECT 1245.840 2.400 1245.980 13.950 ;
        RECT 1263.320 2.400 1263.460 13.950 ;
        RECT 1281.260 2.400 1281.400 13.950 ;
        RECT 1299.200 2.400 1299.340 13.950 ;
        RECT 1317.140 2.400 1317.280 13.950 ;
        RECT 1335.080 2.400 1335.220 13.950 ;
        RECT 1352.560 2.400 1352.700 13.950 ;
        RECT 1370.500 2.400 1370.640 13.950 ;
        RECT 1388.440 2.400 1388.580 13.950 ;
        RECT 1406.380 2.400 1406.520 13.950 ;
        RECT 1423.860 2.400 1424.000 13.950 ;
        RECT 1441.800 2.400 1441.940 13.950 ;
        RECT 1459.740 2.400 1459.880 13.950 ;
        RECT 1477.680 2.400 1477.820 13.950 ;
        RECT 1495.620 2.400 1495.760 13.950 ;
        RECT 1513.100 2.400 1513.240 13.950 ;
        RECT 1531.040 2.400 1531.180 13.950 ;
        RECT 1548.980 2.400 1549.120 13.950 ;
        RECT 1566.920 2.400 1567.060 13.950 ;
        RECT 1584.860 2.400 1585.000 13.950 ;
        RECT 1602.340 2.400 1602.480 13.950 ;
        RECT 1620.280 2.400 1620.420 13.950 ;
        RECT 1638.220 2.400 1638.360 13.950 ;
        RECT 1656.160 2.400 1656.300 13.950 ;
        RECT 1673.640 2.400 1673.780 13.950 ;
        RECT 1691.580 2.400 1691.720 13.950 ;
        RECT 1709.520 2.400 1709.660 13.950 ;
        RECT 1727.460 2.400 1727.600 13.950 ;
        RECT 1745.400 2.400 1745.540 13.950 ;
        RECT 1762.880 2.400 1763.020 13.950 ;
        RECT 1780.820 2.400 1780.960 13.950 ;
        RECT 1798.760 2.400 1798.900 13.950 ;
        RECT 1816.700 2.400 1816.840 13.950 ;
        RECT 1834.640 2.400 1834.780 13.950 ;
        RECT 1852.120 2.400 1852.260 13.950 ;
        RECT 1870.060 2.400 1870.200 13.950 ;
        RECT 1888.000 2.400 1888.140 13.950 ;
        RECT 1905.940 2.400 1906.080 13.950 ;
        RECT 1923.420 2.400 1923.560 13.950 ;
        RECT 1941.360 2.400 1941.500 13.950 ;
        RECT 1959.300 2.400 1959.440 13.950 ;
        RECT 1977.240 2.400 1977.380 13.950 ;
        RECT 1995.180 2.400 1995.320 13.950 ;
        RECT 2012.660 2.400 2012.800 13.950 ;
        RECT 2030.600 2.400 2030.740 13.950 ;
        RECT 2048.540 2.400 2048.680 13.950 ;
        RECT 2066.480 2.400 2066.620 13.950 ;
        RECT 2084.420 2.400 2084.560 13.950 ;
        RECT 2101.900 2.400 2102.040 13.950 ;
        RECT 2119.840 2.400 2119.980 13.950 ;
        RECT 2137.780 2.400 2137.920 13.950 ;
        RECT 2155.720 2.400 2155.860 13.950 ;
        RECT 2173.200 2.400 2173.340 13.950 ;
        RECT 2191.140 2.400 2191.280 13.950 ;
        RECT 2209.080 2.400 2209.220 13.950 ;
        RECT 2227.020 2.400 2227.160 13.950 ;
        RECT 2244.960 2.400 2245.100 13.950 ;
        RECT 2262.440 2.400 2262.580 13.950 ;
        RECT 2280.380 2.400 2280.520 13.950 ;
        RECT 2298.320 2.400 2298.460 13.950 ;
        RECT 2316.260 2.400 2316.400 13.950 ;
        RECT 2334.200 2.400 2334.340 13.950 ;
        RECT 2351.680 2.400 2351.820 13.950 ;
        RECT 2369.620 2.400 2369.760 13.950 ;
        RECT 2387.560 2.400 2387.700 13.950 ;
        RECT 2405.500 2.400 2405.640 13.950 ;
        RECT 2422.980 2.400 2423.120 13.950 ;
        RECT 2440.920 2.400 2441.060 13.950 ;
        RECT 2458.860 2.400 2459.000 13.950 ;
        RECT 2476.800 2.400 2476.940 13.950 ;
        RECT 2494.740 2.400 2494.880 13.950 ;
        RECT 2512.220 2.400 2512.360 13.950 ;
        RECT 2530.160 2.400 2530.300 13.950 ;
        RECT 2548.100 2.400 2548.240 13.950 ;
        RECT 2566.040 2.400 2566.180 13.950 ;
        RECT 2583.980 2.400 2584.120 13.950 ;
        RECT 2601.460 2.400 2601.600 13.950 ;
        RECT 2619.400 2.400 2619.540 13.950 ;
        RECT 2637.340 2.400 2637.480 13.950 ;
        RECT 2655.280 2.400 2655.420 13.950 ;
        RECT 2672.760 2.400 2672.900 13.950 ;
        RECT 2690.700 2.400 2690.840 13.950 ;
        RECT 2708.640 2.400 2708.780 13.950 ;
        RECT 2726.580 2.400 2726.720 13.950 ;
        RECT 2744.520 2.400 2744.660 13.950 ;
        RECT 2762.000 2.400 2762.140 13.950 ;
        RECT 2779.940 2.400 2780.080 13.950 ;
        RECT 2797.880 2.400 2798.020 13.950 ;
        RECT 2815.820 2.400 2815.960 13.950 ;
        RECT 2833.760 2.400 2833.900 13.950 ;
        RECT 2851.240 2.400 2851.380 13.950 ;
        RECT 2869.180 2.400 2869.320 13.950 ;
        RECT 2887.120 2.400 2887.260 13.950 ;
        RECT 2905.060 2.400 2905.200 13.950 ;
        RECT 692.250 -4.800 692.810 2.400 ;
        RECT 710.190 -4.800 710.750 2.400 ;
        RECT 728.130 -4.800 728.690 2.400 ;
        RECT 746.070 -4.800 746.630 2.400 ;
        RECT 763.550 -4.800 764.110 2.400 ;
        RECT 781.490 -4.800 782.050 2.400 ;
        RECT 799.430 -4.800 799.990 2.400 ;
        RECT 817.370 -4.800 817.930 2.400 ;
        RECT 835.310 -4.800 835.870 2.400 ;
        RECT 852.790 -4.800 853.350 2.400 ;
        RECT 870.730 -4.800 871.290 2.400 ;
        RECT 888.670 -4.800 889.230 2.400 ;
        RECT 906.610 -4.800 907.170 2.400 ;
        RECT 924.090 -4.800 924.650 2.400 ;
        RECT 942.030 -4.800 942.590 2.400 ;
        RECT 959.970 -4.800 960.530 2.400 ;
        RECT 977.910 -4.800 978.470 2.400 ;
        RECT 995.850 -4.800 996.410 2.400 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2087.110 902.560 2087.390 902.840 ;
        RECT 1489.570 901.200 1489.850 901.480 ;
        RECT 1489.570 859.040 1489.850 859.320 ;
        RECT 2090.330 858.360 2090.610 858.640 ;
        RECT 1518.090 544.880 1518.370 545.160 ;
        RECT 1538.790 544.880 1539.070 545.160 ;
        RECT 2121.150 544.880 2121.430 545.160 ;
        RECT 2139.090 544.880 2139.370 545.160 ;
      LAYER met3 ;
        RECT 2087.085 902.850 2087.415 902.865 ;
        RECT 2087.085 902.550 2101.890 902.850 ;
        RECT 2087.085 902.535 2087.415 902.550 ;
        RECT 2101.590 901.745 2101.890 902.550 ;
        RECT 1489.545 901.490 1489.875 901.505 ;
        RECT 1500.000 901.490 1504.600 901.745 ;
        RECT 1489.545 901.445 1504.600 901.490 ;
        RECT 2100.000 901.445 2104.600 901.745 ;
        RECT 1489.545 901.190 1501.130 901.445 ;
        RECT 1489.545 901.175 1489.875 901.190 ;
        RECT 1500.830 896.105 1501.130 901.190 ;
        RECT 2101.590 896.105 2101.890 901.445 ;
        RECT 1500.000 895.805 1504.600 896.105 ;
        RECT 2100.000 895.805 2104.600 896.105 ;
        RECT 1500.830 887.605 1501.130 895.805 ;
        RECT 2101.590 887.605 2101.890 895.805 ;
        RECT 1500.000 887.305 1504.600 887.605 ;
        RECT 2100.000 887.305 2104.600 887.605 ;
        RECT 1500.830 881.965 1501.130 887.305 ;
        RECT 2101.590 881.965 2101.890 887.305 ;
        RECT 1500.000 881.665 1504.600 881.965 ;
        RECT 2100.000 881.665 2104.600 881.965 ;
        RECT 1500.830 873.465 1501.130 881.665 ;
        RECT 2101.590 873.465 2101.890 881.665 ;
        RECT 1500.000 873.165 1504.600 873.465 ;
        RECT 2100.000 873.165 2104.600 873.465 ;
        RECT 1500.830 867.825 1501.130 873.165 ;
        RECT 2101.590 867.825 2101.890 873.165 ;
        RECT 1500.000 867.525 1504.600 867.825 ;
        RECT 2100.000 867.525 2104.600 867.825 ;
        RECT 1489.545 859.330 1489.875 859.345 ;
        RECT 1489.545 859.325 1498.370 859.330 ;
        RECT 1500.830 859.325 1501.130 867.525 ;
        RECT 2101.590 859.325 2101.890 867.525 ;
        RECT 1489.545 859.030 1504.600 859.325 ;
        RECT 1489.545 859.015 1489.875 859.030 ;
        RECT 1498.070 859.025 1504.600 859.030 ;
        RECT 2100.000 859.025 2104.600 859.325 ;
        RECT 2090.305 858.650 2090.635 858.665 ;
        RECT 2100.670 858.650 2100.970 859.025 ;
        RECT 2090.305 858.350 2100.970 858.650 ;
        RECT 2090.305 858.335 2090.635 858.350 ;
        RECT 1518.065 545.180 1518.395 545.185 ;
        RECT 1518.065 545.170 1518.650 545.180 ;
        RECT 1538.765 545.170 1539.095 545.185 ;
        RECT 2121.125 545.180 2121.455 545.185 ;
        RECT 1540.350 545.170 1540.730 545.180 ;
        RECT 2120.870 545.170 2121.455 545.180 ;
        RECT 1518.065 544.870 1518.850 545.170 ;
        RECT 1538.765 544.870 1540.730 545.170 ;
        RECT 2120.670 544.870 2121.455 545.170 ;
        RECT 1518.065 544.860 1518.650 544.870 ;
        RECT 1518.065 544.855 1518.395 544.860 ;
        RECT 1538.765 544.855 1539.095 544.870 ;
        RECT 1540.350 544.860 1540.730 544.870 ;
        RECT 2120.870 544.860 2121.455 544.870 ;
        RECT 2121.125 544.855 2121.455 544.860 ;
        RECT 2139.065 545.170 2139.395 545.185 ;
        RECT 2140.190 545.170 2140.570 545.180 ;
        RECT 2139.065 544.870 2140.570 545.170 ;
        RECT 2139.065 544.855 2139.395 544.870 ;
        RECT 2140.190 544.860 2140.570 544.870 ;
      LAYER via3 ;
        RECT 1518.300 544.860 1518.620 545.180 ;
        RECT 1540.380 544.860 1540.700 545.180 ;
        RECT 2120.900 544.860 2121.220 545.180 ;
        RECT 2140.220 544.860 2140.540 545.180 ;
      LAYER met4 ;
        RECT 1518.315 550.950 1518.615 554.600 ;
        RECT 1543.290 550.950 1543.590 554.600 ;
        RECT 1518.310 550.000 1518.615 550.950 ;
        RECT 1540.390 550.650 1543.590 550.950 ;
        RECT 1518.310 545.185 1518.610 550.000 ;
        RECT 1540.390 545.185 1540.690 550.650 ;
        RECT 1543.290 550.000 1543.590 550.650 ;
        RECT 2118.315 550.950 2118.615 554.600 ;
        RECT 2143.290 550.950 2143.590 554.600 ;
        RECT 2118.315 550.650 2121.210 550.950 ;
        RECT 2118.315 550.000 2118.615 550.650 ;
        RECT 2120.910 545.185 2121.210 550.650 ;
        RECT 2140.230 550.650 2143.590 550.950 ;
        RECT 2140.230 545.185 2140.530 550.650 ;
        RECT 2143.290 550.000 2143.590 550.650 ;
        RECT 1518.295 544.855 1518.625 545.185 ;
        RECT 1540.375 544.855 1540.705 545.185 ;
        RECT 2120.895 544.855 2121.225 545.185 ;
        RECT 2140.215 544.855 2140.545 545.185 ;
    END
  END la_data_out[100]
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1881.480 3043.600 1884.050 3044.660 ;
        RECT 2481.480 3043.600 2484.050 3044.660 ;
        RECT 1502.430 561.575 1505.000 562.635 ;
        RECT 2102.430 561.575 2105.000 562.635 ;
      LAYER via3 ;
        RECT 1882.500 3043.620 1884.020 3044.630 ;
        RECT 2482.500 3043.620 2484.020 3044.630 ;
        RECT 1502.460 561.605 1503.980 562.615 ;
        RECT 2102.460 561.605 2103.980 562.615 ;
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 -9.320 367.020 3529.000 ;
        RECT 544.020 -9.320 547.020 3529.000 ;
        RECT 724.020 -9.320 727.020 3529.000 ;
        RECT 904.020 -9.320 907.020 3529.000 ;
        RECT 1084.020 -9.320 1087.020 3529.000 ;
        RECT 1264.020 -9.320 1267.020 3529.000 ;
        RECT 1444.020 2415.000 1447.020 3529.000 ;
        RECT 1624.020 3071.235 1627.020 3529.000 ;
        RECT 1804.020 3071.235 1807.020 3529.000 ;
        RECT 1882.470 2603.670 1884.070 3044.680 ;
        RECT 1624.020 2415.000 1627.020 2585.000 ;
        RECT 1804.020 2415.000 1807.020 2585.000 ;
        RECT 1984.020 2415.000 1987.020 3529.000 ;
        RECT 2164.020 3071.235 2167.020 3529.000 ;
        RECT 2344.020 3071.235 2347.020 3529.000 ;
        RECT 2482.470 2603.670 2484.070 3044.680 ;
        RECT 2164.020 2415.000 2167.020 2585.000 ;
        RECT 2344.020 2415.000 2347.020 2585.000 ;
        RECT 2524.020 2415.000 2527.020 3529.000 ;
        RECT 2704.020 2415.000 2707.020 3529.000 ;
        RECT 1321.040 1210.640 1322.640 2388.880 ;
        RECT 1444.020 -9.320 1447.020 1185.000 ;
        RECT 1624.020 1021.235 1627.020 1185.000 ;
        RECT 1804.020 1021.235 1807.020 1185.000 ;
        RECT 1502.410 561.555 1504.010 1002.565 ;
        RECT 1624.020 -9.320 1627.020 535.000 ;
        RECT 1804.020 -9.320 1807.020 535.000 ;
        RECT 1984.020 -9.320 1987.020 1185.000 ;
        RECT 2164.020 1021.235 2167.020 1185.000 ;
        RECT 2344.020 1021.235 2347.020 1185.000 ;
        RECT 2102.410 561.555 2104.010 1002.565 ;
        RECT 2164.020 -9.320 2167.020 535.000 ;
        RECT 2344.020 -9.320 2347.020 535.000 ;
        RECT 2524.020 -9.320 2527.020 1185.000 ;
        RECT 2704.020 -9.320 2707.020 1185.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1882.680 2891.090 1883.860 2892.270 ;
        RECT 1882.680 2889.490 1883.860 2890.670 ;
        RECT 1882.680 2711.090 1883.860 2712.270 ;
        RECT 1882.680 2709.490 1883.860 2710.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 2482.680 2891.090 2483.860 2892.270 ;
        RECT 2482.680 2889.490 2483.860 2890.670 ;
        RECT 2482.680 2711.090 2483.860 2712.270 ;
        RECT 2482.680 2709.490 2483.860 2710.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1321.250 2351.090 1322.430 2352.270 ;
        RECT 1321.250 2349.490 1322.430 2350.670 ;
        RECT 1321.250 2171.090 1322.430 2172.270 ;
        RECT 1321.250 2169.490 1322.430 2170.670 ;
        RECT 1321.250 1991.090 1322.430 1992.270 ;
        RECT 1321.250 1989.490 1322.430 1990.670 ;
        RECT 1321.250 1811.090 1322.430 1812.270 ;
        RECT 1321.250 1809.490 1322.430 1810.670 ;
        RECT 1321.250 1631.090 1322.430 1632.270 ;
        RECT 1321.250 1629.490 1322.430 1630.670 ;
        RECT 1321.250 1451.090 1322.430 1452.270 ;
        RECT 1321.250 1449.490 1322.430 1450.670 ;
        RECT 1321.250 1271.090 1322.430 1272.270 ;
        RECT 1321.250 1269.490 1322.430 1270.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1502.620 911.090 1503.800 912.270 ;
        RECT 1502.620 909.490 1503.800 910.670 ;
        RECT 1502.620 731.090 1503.800 732.270 ;
        RECT 1502.620 729.490 1503.800 730.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 2102.620 911.090 2103.800 912.270 ;
        RECT 2102.620 909.490 2103.800 910.670 ;
        RECT 2102.620 731.090 2103.800 732.270 ;
        RECT 2102.620 729.490 2103.800 730.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1882.470 2892.380 1884.070 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2482.470 2892.380 2484.070 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1882.470 2889.370 1884.070 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2482.470 2889.370 2484.070 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1882.470 2712.380 1884.070 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2482.470 2712.380 2484.070 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1882.470 2709.370 1884.070 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2482.470 2709.370 2484.070 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1321.040 2352.380 1322.640 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1321.040 2349.370 1322.640 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1321.040 2172.380 1322.640 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1321.040 2169.370 1322.640 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1321.040 1992.380 1322.640 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1321.040 1989.370 1322.640 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1321.040 1812.380 1322.640 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1321.040 1809.370 1322.640 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1321.040 1632.380 1322.640 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1321.040 1629.370 1322.640 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1321.040 1452.380 1322.640 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1321.040 1449.370 1322.640 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1321.040 1272.380 1322.640 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1321.040 1269.370 1322.640 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1502.410 912.380 1504.010 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2102.410 912.380 2104.010 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1502.410 909.370 1504.010 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2102.410 909.370 2104.010 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1502.410 732.380 1504.010 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2102.410 732.380 2104.010 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1502.410 729.370 1504.010 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2102.410 729.370 2104.010 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1881.040 3051.235 1886.300 3052.140 ;
        RECT 2481.040 3051.235 2486.300 3052.140 ;
        RECT 1881.480 3050.400 1886.300 3051.235 ;
        RECT 2481.480 3050.400 2486.300 3051.235 ;
        RECT 1500.180 555.000 1505.000 555.835 ;
        RECT 2100.180 555.000 2105.000 555.835 ;
        RECT 1500.180 554.095 1505.440 555.000 ;
        RECT 2100.180 554.095 2105.440 555.000 ;
      LAYER via3 ;
        RECT 1884.720 3050.440 1886.240 3052.050 ;
        RECT 2484.720 3050.440 2486.240 3052.050 ;
        RECT 1500.240 554.185 1501.760 555.795 ;
        RECT 2100.240 554.185 2101.760 555.795 ;
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 -9.320 457.020 3529.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 -9.320 817.020 3529.000 ;
        RECT 994.020 -9.320 997.020 3529.000 ;
        RECT 1174.020 -9.320 1177.020 3529.000 ;
        RECT 1354.020 2415.000 1357.020 3529.000 ;
        RECT 1534.020 3071.235 1537.020 3529.000 ;
        RECT 1714.020 3071.235 1717.020 3529.000 ;
        RECT 1894.020 3071.235 1897.020 3529.000 ;
        RECT 1884.690 2604.060 1886.310 3052.140 ;
        RECT 1534.020 2415.000 1537.020 2585.000 ;
        RECT 1714.020 2415.000 1717.020 2585.000 ;
        RECT 1894.020 2415.000 1897.020 2585.000 ;
        RECT 2074.020 2415.000 2077.020 3529.000 ;
        RECT 2254.020 3071.235 2257.020 3529.000 ;
        RECT 2434.020 3071.235 2437.020 3529.000 ;
        RECT 2484.690 2604.060 2486.310 3052.140 ;
        RECT 2254.020 2415.000 2257.020 2585.000 ;
        RECT 2434.020 2415.000 2437.020 2585.000 ;
        RECT 2614.020 2415.000 2617.020 3529.000 ;
        RECT 1397.840 1210.640 1399.440 2388.880 ;
        RECT 1354.020 -9.320 1357.020 1185.000 ;
        RECT 1534.020 1021.235 1537.020 1185.000 ;
        RECT 1714.020 1021.235 1717.020 1185.000 ;
        RECT 1894.020 1021.235 1897.020 1185.000 ;
        RECT 1500.170 554.095 1501.790 1002.175 ;
        RECT 1534.020 -9.320 1537.020 535.000 ;
        RECT 1714.020 -9.320 1717.020 535.000 ;
        RECT 1894.020 -9.320 1897.020 535.000 ;
        RECT 2074.020 -9.320 2077.020 1185.000 ;
        RECT 2254.020 1021.235 2257.020 1185.000 ;
        RECT 2434.020 1021.235 2437.020 1185.000 ;
        RECT 2100.170 554.095 2101.790 1002.175 ;
        RECT 2254.020 -9.320 2257.020 535.000 ;
        RECT 2434.020 -9.320 2437.020 535.000 ;
        RECT 2614.020 -9.320 2617.020 1185.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1884.910 2981.090 1886.090 2982.270 ;
        RECT 1884.910 2979.490 1886.090 2980.670 ;
        RECT 1884.910 2801.090 1886.090 2802.270 ;
        RECT 1884.910 2799.490 1886.090 2800.670 ;
        RECT 1884.910 2621.090 1886.090 2622.270 ;
        RECT 1884.910 2619.490 1886.090 2620.670 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 2484.910 2981.090 2486.090 2982.270 ;
        RECT 2484.910 2979.490 2486.090 2980.670 ;
        RECT 2484.910 2801.090 2486.090 2802.270 ;
        RECT 2484.910 2799.490 2486.090 2800.670 ;
        RECT 2484.910 2621.090 2486.090 2622.270 ;
        RECT 2484.910 2619.490 2486.090 2620.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1398.050 2261.090 1399.230 2262.270 ;
        RECT 1398.050 2259.490 1399.230 2260.670 ;
        RECT 1398.050 2081.090 1399.230 2082.270 ;
        RECT 1398.050 2079.490 1399.230 2080.670 ;
        RECT 1398.050 1901.090 1399.230 1902.270 ;
        RECT 1398.050 1899.490 1399.230 1900.670 ;
        RECT 1398.050 1721.090 1399.230 1722.270 ;
        RECT 1398.050 1719.490 1399.230 1720.670 ;
        RECT 1398.050 1541.090 1399.230 1542.270 ;
        RECT 1398.050 1539.490 1399.230 1540.670 ;
        RECT 1398.050 1361.090 1399.230 1362.270 ;
        RECT 1398.050 1359.490 1399.230 1360.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1500.390 821.090 1501.570 822.270 ;
        RECT 1500.390 819.490 1501.570 820.670 ;
        RECT 1500.390 641.090 1501.570 642.270 ;
        RECT 1500.390 639.490 1501.570 640.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2100.390 821.090 2101.570 822.270 ;
        RECT 2100.390 819.490 2101.570 820.670 ;
        RECT 2100.390 641.090 2101.570 642.270 ;
        RECT 2100.390 639.490 2101.570 640.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1884.690 2982.380 1886.310 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2484.690 2982.380 2486.310 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1884.690 2979.370 1886.310 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2484.690 2979.370 2486.310 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1884.690 2802.380 1886.310 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2484.690 2802.380 2486.310 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1884.690 2799.370 1886.310 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2484.690 2799.370 2486.310 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1884.690 2622.380 1886.310 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2484.690 2622.380 2486.310 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1884.690 2619.370 1886.310 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2484.690 2619.370 2486.310 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1397.840 2262.380 1399.440 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1397.840 2259.370 1399.440 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1397.840 2082.380 1399.440 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1397.840 2079.370 1399.440 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1397.840 1902.380 1399.440 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1397.840 1899.370 1399.440 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1397.840 1722.380 1399.440 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1397.840 1719.370 1399.440 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1397.840 1542.380 1399.440 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1397.840 1539.370 1399.440 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1397.840 1362.380 1399.440 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1397.840 1359.370 1399.440 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1500.170 822.380 1501.790 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2100.170 822.380 2101.790 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1500.170 819.370 1501.790 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2100.170 819.370 2101.790 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1500.170 642.380 1501.790 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2100.170 642.380 2101.790 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1500.170 639.370 1501.790 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2100.170 639.370 2101.790 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 -18.720 385.020 3538.400 ;
        RECT 562.020 -18.720 565.020 3538.400 ;
        RECT 742.020 -18.720 745.020 3538.400 ;
        RECT 922.020 -18.720 925.020 3538.400 ;
        RECT 1102.020 -18.720 1105.020 3538.400 ;
        RECT 1282.020 2415.000 1285.020 3538.400 ;
        RECT 1462.020 2415.000 1465.020 3538.400 ;
        RECT 1642.020 3071.235 1645.020 3538.400 ;
        RECT 1822.020 3071.235 1825.020 3538.400 ;
        RECT 1642.020 2415.000 1645.020 2585.000 ;
        RECT 1822.020 2415.000 1825.020 2585.000 ;
        RECT 2002.020 2415.000 2005.020 3538.400 ;
        RECT 2182.020 3071.235 2185.020 3538.400 ;
        RECT 2362.020 3071.235 2365.020 3538.400 ;
        RECT 2182.020 2415.000 2185.020 2585.000 ;
        RECT 2362.020 2415.000 2365.020 2585.000 ;
        RECT 2542.020 2415.000 2545.020 3538.400 ;
        RECT 1282.020 -18.720 1285.020 1185.000 ;
        RECT 1462.020 -18.720 1465.020 1185.000 ;
        RECT 1642.020 1021.235 1645.020 1185.000 ;
        RECT 1822.020 1021.235 1825.020 1185.000 ;
        RECT 1642.020 -18.720 1645.020 535.000 ;
        RECT 1822.020 -18.720 1825.020 535.000 ;
        RECT 2002.020 -18.720 2005.020 1185.000 ;
        RECT 2182.020 1021.235 2185.020 1185.000 ;
        RECT 2362.020 1021.235 2365.020 1185.000 ;
        RECT 2182.020 -18.720 2185.020 535.000 ;
        RECT 2362.020 -18.720 2365.020 535.000 ;
        RECT 2542.020 -18.720 2545.020 1185.000 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 -18.720 475.020 3538.400 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 -18.720 835.020 3538.400 ;
        RECT 1012.020 -18.720 1015.020 3538.400 ;
        RECT 1192.020 -18.720 1195.020 3538.400 ;
        RECT 1372.020 2415.000 1375.020 3538.400 ;
        RECT 1552.020 3071.235 1555.020 3538.400 ;
        RECT 1732.020 3071.235 1735.020 3538.400 ;
        RECT 1552.020 2415.000 1555.020 2585.000 ;
        RECT 1732.020 2415.000 1735.020 2585.000 ;
        RECT 1912.020 2415.000 1915.020 3538.400 ;
        RECT 2092.020 3071.235 2095.020 3538.400 ;
        RECT 2272.020 3071.235 2275.020 3538.400 ;
        RECT 2452.020 3071.235 2455.020 3538.400 ;
        RECT 2092.020 2415.000 2095.020 2585.000 ;
        RECT 2272.020 2415.000 2275.020 2585.000 ;
        RECT 2452.020 2415.000 2455.020 2585.000 ;
        RECT 2632.020 2415.000 2635.020 3538.400 ;
        RECT 1372.020 -18.720 1375.020 1185.000 ;
        RECT 1552.020 -18.720 1555.020 535.000 ;
        RECT 1732.020 -18.720 1735.020 535.000 ;
        RECT 1912.020 -18.720 1915.020 1185.000 ;
        RECT 2092.020 -18.720 2095.020 535.000 ;
        RECT 2272.020 -18.720 2275.020 535.000 ;
        RECT 2452.020 -18.720 2455.020 535.000 ;
        RECT 2632.020 -18.720 2635.020 1185.000 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 -28.120 403.020 3547.800 ;
        RECT 580.020 -28.120 583.020 3547.800 ;
        RECT 760.020 -28.120 763.020 3547.800 ;
        RECT 940.020 -28.120 943.020 3547.800 ;
        RECT 1120.020 -28.120 1123.020 3547.800 ;
        RECT 1300.020 2415.000 1303.020 3547.800 ;
        RECT 1480.020 2415.000 1483.020 3547.800 ;
        RECT 1660.020 3071.235 1663.020 3547.800 ;
        RECT 1840.020 3071.235 1843.020 3547.800 ;
        RECT 1660.020 2415.000 1663.020 2585.000 ;
        RECT 1840.020 2415.000 1843.020 2585.000 ;
        RECT 2020.020 2415.000 2023.020 3547.800 ;
        RECT 2200.020 3071.235 2203.020 3547.800 ;
        RECT 2380.020 3071.235 2383.020 3547.800 ;
        RECT 2200.020 2415.000 2203.020 2585.000 ;
        RECT 2380.020 2415.000 2383.020 2585.000 ;
        RECT 2560.020 2415.000 2563.020 3547.800 ;
        RECT 1300.020 -28.120 1303.020 1185.000 ;
        RECT 1480.020 -28.120 1483.020 1185.000 ;
        RECT 1660.020 1021.235 1663.020 1185.000 ;
        RECT 1840.020 1021.235 1843.020 1185.000 ;
        RECT 1660.020 -28.120 1663.020 535.000 ;
        RECT 1840.020 -28.120 1843.020 535.000 ;
        RECT 2020.020 -28.120 2023.020 1185.000 ;
        RECT 2200.020 1021.235 2203.020 1185.000 ;
        RECT 2380.020 1021.235 2383.020 1185.000 ;
        RECT 2200.020 -28.120 2203.020 535.000 ;
        RECT 2380.020 -28.120 2383.020 535.000 ;
        RECT 2560.020 -28.120 2563.020 1185.000 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 -28.120 493.020 3547.800 ;
        RECT 670.020 -28.120 673.020 3547.800 ;
        RECT 850.020 -28.120 853.020 3547.800 ;
        RECT 1030.020 -28.120 1033.020 3547.800 ;
        RECT 1210.020 -28.120 1213.020 3547.800 ;
        RECT 1390.020 2415.000 1393.020 3547.800 ;
        RECT 1570.020 3071.235 1573.020 3547.800 ;
        RECT 1750.020 3071.235 1753.020 3547.800 ;
        RECT 1570.020 2415.000 1573.020 2585.000 ;
        RECT 1750.020 2415.000 1753.020 2585.000 ;
        RECT 1930.020 2415.000 1933.020 3547.800 ;
        RECT 2110.020 3071.235 2113.020 3547.800 ;
        RECT 2290.020 3071.235 2293.020 3547.800 ;
        RECT 2470.020 3071.235 2473.020 3547.800 ;
        RECT 2110.020 2415.000 2113.020 2585.000 ;
        RECT 2290.020 2415.000 2293.020 2585.000 ;
        RECT 2470.020 2415.000 2473.020 2585.000 ;
        RECT 2650.020 2415.000 2653.020 3547.800 ;
        RECT 1390.020 -28.120 1393.020 1185.000 ;
        RECT 1570.020 1021.235 1573.020 1185.000 ;
        RECT 1750.020 1021.235 1753.020 1185.000 ;
        RECT 1570.020 -28.120 1573.020 535.000 ;
        RECT 1750.020 -28.120 1753.020 535.000 ;
        RECT 1930.020 -28.120 1933.020 1185.000 ;
        RECT 2110.020 1021.235 2113.020 1185.000 ;
        RECT 2290.020 1021.235 2293.020 1185.000 ;
        RECT 2470.020 1021.235 2473.020 1185.000 ;
        RECT 2110.020 -28.120 2113.020 535.000 ;
        RECT 2290.020 -28.120 2293.020 535.000 ;
        RECT 2470.020 -28.120 2473.020 535.000 ;
        RECT 2650.020 -28.120 2653.020 1185.000 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 -37.520 421.020 3557.200 ;
        RECT 598.020 -37.520 601.020 3557.200 ;
        RECT 778.020 -37.520 781.020 3557.200 ;
        RECT 958.020 -37.520 961.020 3557.200 ;
        RECT 1138.020 -37.520 1141.020 3557.200 ;
        RECT 1318.020 2415.000 1321.020 3557.200 ;
        RECT 1498.020 3071.235 1501.020 3557.200 ;
        RECT 1678.020 3071.235 1681.020 3557.200 ;
        RECT 1858.020 3071.235 1861.020 3557.200 ;
        RECT 2038.020 2415.000 2041.020 3557.200 ;
        RECT 2218.020 3071.235 2221.020 3557.200 ;
        RECT 2398.020 3071.235 2401.020 3557.200 ;
        RECT 2578.020 2415.000 2581.020 3557.200 ;
        RECT 1318.020 -37.520 1321.020 1185.000 ;
        RECT 1498.020 1021.235 1501.020 1185.000 ;
        RECT 1678.020 1021.235 1681.020 1185.000 ;
        RECT 1858.020 1021.235 1861.020 1185.000 ;
        RECT 1498.020 -37.520 1501.020 535.000 ;
        RECT 1678.020 -37.520 1681.020 535.000 ;
        RECT 1858.020 -37.520 1861.020 535.000 ;
        RECT 2038.020 -37.520 2041.020 1185.000 ;
        RECT 2218.020 1021.235 2221.020 1185.000 ;
        RECT 2398.020 1021.235 2401.020 1185.000 ;
        RECT 2218.020 -37.520 2221.020 535.000 ;
        RECT 2398.020 -37.520 2401.020 535.000 ;
        RECT 2578.020 -37.520 2581.020 1185.000 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 -37.520 511.020 3557.200 ;
        RECT 688.020 -37.520 691.020 3557.200 ;
        RECT 868.020 -37.520 871.020 3557.200 ;
        RECT 1048.020 -37.520 1051.020 3557.200 ;
        RECT 1228.020 -37.520 1231.020 3557.200 ;
        RECT 1408.020 2415.000 1411.020 3557.200 ;
        RECT 1588.020 3071.235 1591.020 3557.200 ;
        RECT 1768.020 3071.235 1771.020 3557.200 ;
        RECT 1588.020 2415.000 1591.020 2585.000 ;
        RECT 1768.020 2415.000 1771.020 2585.000 ;
        RECT 1948.020 2415.000 1951.020 3557.200 ;
        RECT 2128.020 3071.235 2131.020 3557.200 ;
        RECT 2308.020 3071.235 2311.020 3557.200 ;
        RECT 2488.020 3071.235 2491.020 3557.200 ;
        RECT 2128.020 2415.000 2131.020 2585.000 ;
        RECT 2308.020 2415.000 2311.020 2585.000 ;
        RECT 2488.020 2415.000 2491.020 2585.000 ;
        RECT 2668.020 2415.000 2671.020 3557.200 ;
        RECT 1408.020 -37.520 1411.020 1185.000 ;
        RECT 1588.020 1021.235 1591.020 1185.000 ;
        RECT 1768.020 1021.235 1771.020 1185.000 ;
        RECT 1588.020 -37.520 1591.020 535.000 ;
        RECT 1768.020 -37.520 1771.020 535.000 ;
        RECT 1948.020 -37.520 1951.020 1185.000 ;
        RECT 2128.020 1021.235 2131.020 1185.000 ;
        RECT 2308.020 1021.235 2311.020 1185.000 ;
        RECT 2488.020 1021.235 2491.020 1185.000 ;
        RECT 2128.020 -37.520 2131.020 535.000 ;
        RECT 2308.020 -37.520 2311.020 535.000 ;
        RECT 2488.020 -37.520 2491.020 535.000 ;
        RECT 2668.020 -37.520 2671.020 1185.000 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
        RECT 1305.520 1205.865 2694.260 2388.725 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met1 ;
        RECT 2442.670 3067.040 2442.990 3067.100 ;
        RECT 2469.810 3067.040 2470.130 3067.100 ;
        RECT 2442.670 3066.900 2470.130 3067.040 ;
        RECT 2442.670 3066.840 2442.990 3066.900 ;
        RECT 2469.810 3066.840 2470.130 3066.900 ;
        RECT 1868.130 3063.980 1868.450 3064.040 ;
        RECT 1898.030 3063.980 1898.350 3064.040 ;
        RECT 2442.670 3063.980 2442.990 3064.040 ;
        RECT 1868.130 3063.840 2442.990 3063.980 ;
        RECT 1868.130 3063.780 1868.450 3063.840 ;
        RECT 1898.030 3063.780 1898.350 3063.840 ;
        RECT 2442.670 3063.780 2442.990 3063.840 ;
        RECT 2469.810 3063.980 2470.130 3064.040 ;
        RECT 2497.870 3063.980 2498.190 3064.040 ;
        RECT 2469.810 3063.840 2498.190 3063.980 ;
        RECT 2469.810 3063.780 2470.130 3063.840 ;
        RECT 2497.870 3063.780 2498.190 3063.840 ;
        RECT 1899.870 3052.080 1900.190 3052.140 ;
        RECT 2482.230 3052.080 2482.550 3052.140 ;
        RECT 1899.870 3051.940 2482.550 3052.080 ;
        RECT 1899.870 3051.880 1900.190 3051.940 ;
        RECT 2482.230 3051.880 2482.550 3051.940 ;
      LAYER met1 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
      LAYER met1 ;
        RECT 1938.510 3029.300 1938.830 3029.360 ;
        RECT 2083.870 3029.300 2084.190 3029.360 ;
        RECT 1938.510 3029.160 2084.190 3029.300 ;
        RECT 1938.510 3029.100 1938.830 3029.160 ;
        RECT 2083.870 3029.100 2084.190 3029.160 ;
        RECT 1924.710 3022.500 1925.030 3022.560 ;
        RECT 2083.870 3022.500 2084.190 3022.560 ;
        RECT 1924.710 3022.360 2084.190 3022.500 ;
        RECT 1924.710 3022.300 1925.030 3022.360 ;
        RECT 2083.870 3022.300 2084.190 3022.360 ;
        RECT 1910.910 3015.700 1911.230 3015.760 ;
        RECT 2083.870 3015.700 2084.190 3015.760 ;
        RECT 1910.910 3015.560 2084.190 3015.700 ;
        RECT 1910.910 3015.500 1911.230 3015.560 ;
        RECT 2083.870 3015.500 2084.190 3015.560 ;
        RECT 1897.110 3008.560 1897.430 3008.620 ;
        RECT 2083.870 3008.560 2084.190 3008.620 ;
        RECT 1897.110 3008.420 2084.190 3008.560 ;
        RECT 1897.110 3008.360 1897.430 3008.420 ;
        RECT 2083.870 3008.360 2084.190 3008.420 ;
        RECT 1890.210 3001.760 1890.530 3001.820 ;
        RECT 2083.870 3001.760 2084.190 3001.820 ;
        RECT 1890.210 3001.620 2084.190 3001.760 ;
        RECT 1890.210 3001.560 1890.530 3001.620 ;
        RECT 2083.870 3001.560 2084.190 3001.620 ;
        RECT 2069.610 2698.140 2069.930 2698.200 ;
        RECT 2084.790 2698.140 2085.110 2698.200 ;
        RECT 2069.610 2698.000 2085.110 2698.140 ;
        RECT 2069.610 2697.940 2069.930 2698.000 ;
        RECT 2084.790 2697.940 2085.110 2698.000 ;
        RECT 1897.570 2691.340 1897.890 2691.400 ;
        RECT 1898.950 2691.340 1899.270 2691.400 ;
        RECT 1897.570 2691.200 1899.270 2691.340 ;
        RECT 1897.570 2691.140 1897.890 2691.200 ;
        RECT 1898.950 2691.140 1899.270 2691.200 ;
        RECT 2052.590 2691.340 2052.910 2691.400 ;
        RECT 2083.870 2691.340 2084.190 2691.400 ;
        RECT 2052.590 2691.200 2084.190 2691.340 ;
        RECT 2052.590 2691.140 2052.910 2691.200 ;
        RECT 2083.870 2691.140 2084.190 2691.200 ;
        RECT 1897.570 2680.460 1897.890 2680.520 ;
        RECT 1898.950 2680.460 1899.270 2680.520 ;
        RECT 1897.570 2680.320 1899.270 2680.460 ;
        RECT 1897.570 2680.260 1897.890 2680.320 ;
        RECT 1898.950 2680.260 1899.270 2680.320 ;
        RECT 2049.370 2608.040 2049.690 2608.100 ;
        RECT 2052.590 2608.040 2052.910 2608.100 ;
        RECT 2049.370 2607.900 2052.910 2608.040 ;
        RECT 2049.370 2607.840 2049.690 2607.900 ;
        RECT 2052.590 2607.840 2052.910 2607.900 ;
      LAYER met1 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met1 ;
        RECT 1486.330 2604.640 1486.650 2604.700 ;
        RECT 2049.370 2604.640 2049.690 2604.700 ;
        RECT 1486.330 2604.500 2049.690 2604.640 ;
        RECT 1486.330 2604.440 1486.650 2604.500 ;
        RECT 2049.370 2604.440 2049.690 2604.500 ;
        RECT 1898.030 2594.780 1898.350 2594.840 ;
        RECT 1898.950 2594.780 1899.270 2594.840 ;
        RECT 1898.030 2594.640 1899.270 2594.780 ;
        RECT 1898.030 2594.580 1898.350 2594.640 ;
        RECT 1898.950 2594.580 1899.270 2594.640 ;
        RECT 1600.410 2594.440 1600.730 2594.500 ;
        RECT 1644.570 2594.440 1644.890 2594.500 ;
        RECT 1648.250 2594.440 1648.570 2594.500 ;
        RECT 1600.410 2594.300 1648.570 2594.440 ;
        RECT 1600.410 2594.240 1600.730 2594.300 ;
        RECT 1644.570 2594.240 1644.890 2594.300 ;
        RECT 1648.250 2594.240 1648.570 2594.300 ;
        RECT 1744.850 2594.440 1745.170 2594.500 ;
        RECT 2277.070 2594.440 2277.390 2594.500 ;
        RECT 1744.850 2594.300 2277.390 2594.440 ;
        RECT 1744.850 2594.240 1745.170 2594.300 ;
        RECT 2277.070 2594.240 2277.390 2594.300 ;
        RECT 1448.610 2594.100 1448.930 2594.160 ;
        RECT 1614.670 2594.100 1614.990 2594.160 ;
        RECT 1448.610 2593.960 1614.990 2594.100 ;
        RECT 1448.610 2593.900 1448.930 2593.960 ;
        RECT 1614.670 2593.900 1614.990 2593.960 ;
        RECT 1636.750 2594.100 1637.070 2594.160 ;
        RECT 1684.590 2594.100 1684.910 2594.160 ;
        RECT 1636.750 2593.960 1684.910 2594.100 ;
        RECT 1636.750 2593.900 1637.070 2593.960 ;
        RECT 1684.590 2593.900 1684.910 2593.960 ;
        RECT 1726.450 2594.100 1726.770 2594.160 ;
        RECT 2242.570 2594.100 2242.890 2594.160 ;
        RECT 1726.450 2593.960 2242.890 2594.100 ;
        RECT 1726.450 2593.900 1726.770 2593.960 ;
        RECT 2242.570 2593.900 2242.890 2593.960 ;
        RECT 2243.490 2594.100 2243.810 2594.160 ;
        RECT 2291.790 2594.100 2292.110 2594.160 ;
        RECT 2243.490 2593.960 2292.110 2594.100 ;
        RECT 2243.490 2593.900 2243.810 2593.960 ;
        RECT 2291.790 2593.900 2292.110 2593.960 ;
        RECT 1538.310 2593.760 1538.630 2593.820 ;
        RECT 1656.530 2593.760 1656.850 2593.820 ;
        RECT 1538.310 2593.620 1656.850 2593.760 ;
        RECT 1538.310 2593.560 1538.630 2593.620 ;
        RECT 1656.530 2593.560 1656.850 2593.620 ;
        RECT 1656.990 2593.760 1657.310 2593.820 ;
        RECT 1702.990 2593.760 1703.310 2593.820 ;
        RECT 1656.990 2593.620 1703.310 2593.760 ;
        RECT 1656.990 2593.560 1657.310 2593.620 ;
        RECT 1702.990 2593.560 1703.310 2593.620 ;
        RECT 1732.890 2593.760 1733.210 2593.820 ;
        RECT 2249.470 2593.760 2249.790 2593.820 ;
        RECT 1732.890 2593.620 2249.790 2593.760 ;
        RECT 1732.890 2593.560 1733.210 2593.620 ;
        RECT 2249.470 2593.560 2249.790 2593.620 ;
        RECT 2256.370 2593.760 2256.690 2593.820 ;
        RECT 2297.770 2593.760 2298.090 2593.820 ;
        RECT 2256.370 2593.620 2298.090 2593.760 ;
        RECT 2256.370 2593.560 2256.690 2593.620 ;
        RECT 2297.770 2593.560 2298.090 2593.620 ;
        RECT 1572.810 2593.420 1573.130 2593.480 ;
        RECT 1615.590 2593.420 1615.910 2593.480 ;
        RECT 1662.050 2593.420 1662.370 2593.480 ;
        RECT 1707.590 2593.420 1707.910 2593.480 ;
        RECT 1572.810 2593.280 1707.910 2593.420 ;
        RECT 1572.810 2593.220 1573.130 2593.280 ;
        RECT 1615.590 2593.220 1615.910 2593.280 ;
        RECT 1662.050 2593.220 1662.370 2593.280 ;
        RECT 1707.590 2593.220 1707.910 2593.280 ;
        RECT 2215.890 2593.420 2216.210 2593.480 ;
        RECT 2262.810 2593.420 2263.130 2593.480 ;
        RECT 2285.350 2593.420 2285.670 2593.480 ;
        RECT 2332.270 2593.420 2332.590 2593.480 ;
        RECT 2215.890 2593.280 2263.960 2593.420 ;
        RECT 2215.890 2593.220 2216.210 2593.280 ;
        RECT 2262.810 2593.220 2263.130 2593.280 ;
        RECT 1593.510 2593.080 1593.830 2593.140 ;
        RECT 1636.750 2593.080 1637.070 2593.140 ;
        RECT 1593.510 2592.940 1637.070 2593.080 ;
        RECT 1593.510 2592.880 1593.830 2592.940 ;
        RECT 1636.750 2592.880 1637.070 2592.940 ;
        RECT 1648.250 2593.080 1648.570 2593.140 ;
        RECT 1690.570 2593.080 1690.890 2593.140 ;
        RECT 1738.410 2593.080 1738.730 2593.140 ;
        RECT 2263.270 2593.080 2263.590 2593.140 ;
        RECT 1648.250 2592.940 2263.590 2593.080 ;
        RECT 1648.250 2592.880 1648.570 2592.940 ;
        RECT 1690.570 2592.880 1690.890 2592.940 ;
        RECT 1738.410 2592.880 1738.730 2592.940 ;
        RECT 2263.270 2592.880 2263.590 2592.940 ;
        RECT 1605.470 2592.740 1605.790 2592.800 ;
        RECT 1650.550 2592.740 1650.870 2592.800 ;
        RECT 1697.470 2592.740 1697.790 2592.800 ;
        RECT 1744.850 2592.740 1745.170 2592.800 ;
        RECT 1605.470 2592.600 1745.170 2592.740 ;
        RECT 1605.470 2592.540 1605.790 2592.600 ;
        RECT 1650.550 2592.540 1650.870 2592.600 ;
        RECT 1697.470 2592.540 1697.790 2592.600 ;
        RECT 1744.850 2592.540 1745.170 2592.600 ;
        RECT 2212.670 2592.740 2212.990 2592.800 ;
        RECT 2256.370 2592.740 2256.690 2592.800 ;
        RECT 2212.670 2592.600 2256.690 2592.740 ;
        RECT 2263.820 2592.740 2263.960 2593.280 ;
        RECT 2285.350 2593.280 2332.590 2593.420 ;
        RECT 2285.350 2593.220 2285.670 2593.280 ;
        RECT 2332.270 2593.220 2332.590 2593.280 ;
        RECT 2305.130 2592.740 2305.450 2592.800 ;
        RECT 2263.820 2592.600 2305.450 2592.740 ;
        RECT 2212.670 2592.540 2212.990 2592.600 ;
        RECT 2256.370 2592.540 2256.690 2592.600 ;
        RECT 2305.130 2592.540 2305.450 2592.600 ;
        RECT 1372.710 2592.400 1373.030 2592.460 ;
        RECT 1580.170 2592.400 1580.490 2592.460 ;
        RECT 1372.710 2592.260 1580.490 2592.400 ;
        RECT 1372.710 2592.200 1373.030 2592.260 ;
        RECT 1580.170 2592.200 1580.490 2592.260 ;
        RECT 1586.610 2592.400 1586.930 2592.460 ;
        RECT 1632.150 2592.400 1632.470 2592.460 ;
        RECT 1679.070 2592.400 1679.390 2592.460 ;
        RECT 1726.450 2592.400 1726.770 2592.460 ;
        RECT 1586.610 2592.260 1726.770 2592.400 ;
        RECT 1586.610 2592.200 1586.930 2592.260 ;
        RECT 1632.150 2592.200 1632.470 2592.260 ;
        RECT 1679.070 2592.200 1679.390 2592.260 ;
        RECT 1726.450 2592.200 1726.770 2592.260 ;
        RECT 2239.810 2592.400 2240.130 2592.460 ;
        RECT 2285.350 2592.400 2285.670 2592.460 ;
        RECT 2239.810 2592.260 2285.670 2592.400 ;
        RECT 2239.810 2592.200 2240.130 2592.260 ;
        RECT 2285.350 2592.200 2285.670 2592.260 ;
        RECT 2291.790 2592.400 2292.110 2592.460 ;
        RECT 2332.270 2592.400 2332.590 2592.460 ;
        RECT 2291.790 2592.260 2332.590 2592.400 ;
        RECT 2291.790 2592.200 2292.110 2592.260 ;
        RECT 2332.270 2592.200 2332.590 2592.260 ;
        RECT 1565.910 2592.060 1566.230 2592.120 ;
        RECT 1586.150 2592.060 1586.470 2592.120 ;
        RECT 1627.090 2592.060 1627.410 2592.120 ;
        RECT 1565.910 2591.920 1585.460 2592.060 ;
        RECT 1565.910 2591.860 1566.230 2591.920 ;
        RECT 1358.910 2591.720 1359.230 2591.780 ;
        RECT 1573.270 2591.720 1573.590 2591.780 ;
        RECT 1358.910 2591.580 1573.590 2591.720 ;
        RECT 1585.320 2591.720 1585.460 2591.920 ;
        RECT 1586.150 2591.920 1627.410 2592.060 ;
        RECT 1586.150 2591.860 1586.470 2591.920 ;
        RECT 1627.090 2591.860 1627.410 2591.920 ;
        RECT 1627.550 2592.060 1627.870 2592.120 ;
        RECT 1656.990 2592.060 1657.310 2592.120 ;
        RECT 1627.550 2591.920 1657.310 2592.060 ;
        RECT 1627.550 2591.860 1627.870 2591.920 ;
        RECT 1656.990 2591.860 1657.310 2591.920 ;
        RECT 1668.950 2592.060 1669.270 2592.120 ;
        RECT 1714.950 2592.060 1715.270 2592.120 ;
        RECT 1668.950 2591.920 1715.270 2592.060 ;
        RECT 1668.950 2591.860 1669.270 2591.920 ;
        RECT 1714.950 2591.860 1715.270 2591.920 ;
        RECT 1848.810 2592.060 1849.130 2592.120 ;
        RECT 2132.170 2592.060 2132.490 2592.120 ;
        RECT 1848.810 2591.920 2132.490 2592.060 ;
        RECT 1848.810 2591.860 1849.130 2591.920 ;
        RECT 2132.170 2591.860 2132.490 2591.920 ;
        RECT 2221.410 2592.060 2221.730 2592.120 ;
        RECT 2268.790 2592.060 2269.110 2592.120 ;
        RECT 2311.570 2592.060 2311.890 2592.120 ;
        RECT 2221.410 2591.920 2311.890 2592.060 ;
        RECT 2221.410 2591.860 2221.730 2591.920 ;
        RECT 2268.790 2591.860 2269.110 2591.920 ;
        RECT 2311.570 2591.860 2311.890 2591.920 ;
        RECT 1593.970 2591.720 1594.290 2591.780 ;
        RECT 1585.320 2591.580 1594.290 2591.720 ;
        RECT 1358.910 2591.520 1359.230 2591.580 ;
        RECT 1573.270 2591.520 1573.590 2591.580 ;
        RECT 1593.970 2591.520 1594.290 2591.580 ;
        RECT 1684.590 2591.720 1684.910 2591.780 ;
        RECT 1732.890 2591.720 1733.210 2591.780 ;
        RECT 1684.590 2591.580 1733.210 2591.720 ;
        RECT 1684.590 2591.520 1684.910 2591.580 ;
        RECT 1732.890 2591.520 1733.210 2591.580 ;
        RECT 1786.710 2591.720 1787.030 2591.780 ;
        RECT 2152.870 2591.720 2153.190 2591.780 ;
        RECT 1786.710 2591.580 2153.190 2591.720 ;
        RECT 1786.710 2591.520 1787.030 2591.580 ;
        RECT 2152.870 2591.520 2153.190 2591.580 ;
        RECT 2179.550 2591.720 2179.870 2591.780 ;
        RECT 2221.500 2591.720 2221.640 2591.860 ;
        RECT 2179.550 2591.580 2221.640 2591.720 ;
        RECT 2226.930 2591.720 2227.250 2591.780 ;
        RECT 2276.610 2591.720 2276.930 2591.780 ;
        RECT 2318.470 2591.720 2318.790 2591.780 ;
        RECT 2226.930 2591.580 2318.790 2591.720 ;
        RECT 2179.550 2591.520 2179.870 2591.580 ;
        RECT 2226.930 2591.520 2227.250 2591.580 ;
        RECT 2276.610 2591.520 2276.930 2591.580 ;
        RECT 2318.470 2591.520 2318.790 2591.580 ;
        RECT 1345.110 2591.380 1345.430 2591.440 ;
        RECT 1566.370 2591.380 1566.690 2591.440 ;
        RECT 1345.110 2591.240 1566.690 2591.380 ;
        RECT 1345.110 2591.180 1345.430 2591.240 ;
        RECT 1566.370 2591.180 1566.690 2591.240 ;
        RECT 1579.250 2591.380 1579.570 2591.440 ;
        RECT 1600.870 2591.380 1601.190 2591.440 ;
        RECT 1579.250 2591.240 1601.190 2591.380 ;
        RECT 1579.250 2591.180 1579.570 2591.240 ;
        RECT 1600.870 2591.180 1601.190 2591.240 ;
        RECT 1627.090 2591.380 1627.410 2591.440 ;
        RECT 1673.550 2591.380 1673.870 2591.440 ;
        RECT 1718.630 2591.380 1718.950 2591.440 ;
        RECT 1721.850 2591.380 1722.170 2591.440 ;
        RECT 1627.090 2591.240 1722.170 2591.380 ;
        RECT 1627.090 2591.180 1627.410 2591.240 ;
        RECT 1673.550 2591.180 1673.870 2591.240 ;
        RECT 1718.630 2591.180 1718.950 2591.240 ;
        RECT 1721.850 2591.180 1722.170 2591.240 ;
        RECT 1772.910 2591.380 1773.230 2591.440 ;
        RECT 2146.430 2591.380 2146.750 2591.440 ;
        RECT 1772.910 2591.240 2146.750 2591.380 ;
        RECT 1772.910 2591.180 1773.230 2591.240 ;
        RECT 2146.430 2591.180 2146.750 2591.240 ;
        RECT 2184.610 2591.040 2184.930 2591.100 ;
        RECT 2227.020 2591.040 2227.160 2591.520 ;
        RECT 2231.990 2591.380 2232.310 2591.440 ;
        RECT 2280.290 2591.380 2280.610 2591.440 ;
        RECT 2325.370 2591.380 2325.690 2591.440 ;
        RECT 2231.990 2591.240 2325.690 2591.380 ;
        RECT 2231.990 2591.180 2232.310 2591.240 ;
        RECT 2280.290 2591.180 2280.610 2591.240 ;
        RECT 2325.370 2591.180 2325.690 2591.240 ;
        RECT 2250.850 2591.040 2251.170 2591.100 ;
        RECT 2297.770 2591.040 2298.090 2591.100 ;
        RECT 2339.170 2591.040 2339.490 2591.100 ;
        RECT 2184.610 2590.900 2227.160 2591.040 ;
        RECT 2238.980 2590.900 2339.490 2591.040 ;
        RECT 2184.610 2590.840 2184.930 2590.900 ;
        RECT 1434.810 2590.700 1435.130 2590.760 ;
        RECT 1608.690 2590.700 1609.010 2590.760 ;
        RECT 1434.810 2590.560 1609.010 2590.700 ;
        RECT 1434.810 2590.500 1435.130 2590.560 ;
        RECT 1608.690 2590.500 1609.010 2590.560 ;
        RECT 1655.610 2590.700 1655.930 2590.760 ;
        RECT 1704.370 2590.700 1704.690 2590.760 ;
        RECT 1655.610 2590.560 1704.690 2590.700 ;
        RECT 1655.610 2590.500 1655.930 2590.560 ;
        RECT 1704.370 2590.500 1704.690 2590.560 ;
        RECT 1759.110 2590.700 1759.430 2590.760 ;
        RECT 2145.970 2590.700 2146.290 2590.760 ;
        RECT 1759.110 2590.560 2146.290 2590.700 ;
        RECT 1759.110 2590.500 1759.430 2590.560 ;
        RECT 2145.970 2590.500 2146.290 2590.560 ;
        RECT 2204.390 2590.700 2204.710 2590.760 ;
        RECT 2238.980 2590.700 2239.120 2590.900 ;
        RECT 2250.850 2590.840 2251.170 2590.900 ;
        RECT 2297.770 2590.840 2298.090 2590.900 ;
        RECT 2339.170 2590.840 2339.490 2590.900 ;
        RECT 2204.390 2590.560 2239.120 2590.700 ;
        RECT 2204.390 2590.500 2204.710 2590.560 ;
        RECT 1427.910 2590.360 1428.230 2590.420 ;
        RECT 1579.250 2590.360 1579.570 2590.420 ;
        RECT 1427.910 2590.220 1579.570 2590.360 ;
        RECT 1427.910 2590.160 1428.230 2590.220 ;
        RECT 1579.250 2590.160 1579.570 2590.220 ;
        RECT 1579.710 2590.360 1580.030 2590.420 ;
        RECT 1621.570 2590.360 1621.890 2590.420 ;
        RECT 1627.550 2590.360 1627.870 2590.420 ;
        RECT 1579.710 2590.220 1627.870 2590.360 ;
        RECT 1579.710 2590.160 1580.030 2590.220 ;
        RECT 1621.570 2590.160 1621.890 2590.220 ;
        RECT 1627.550 2590.160 1627.870 2590.220 ;
        RECT 1628.010 2590.360 1628.330 2590.420 ;
        RECT 1697.470 2590.360 1697.790 2590.420 ;
        RECT 1628.010 2590.220 1697.790 2590.360 ;
        RECT 1628.010 2590.160 1628.330 2590.220 ;
        RECT 1697.470 2590.160 1697.790 2590.220 ;
        RECT 1745.310 2590.360 1745.630 2590.420 ;
        RECT 2126.650 2590.360 2126.970 2590.420 ;
        RECT 1745.310 2590.220 2126.970 2590.360 ;
        RECT 1745.310 2590.160 1745.630 2590.220 ;
        RECT 2126.650 2590.160 2126.970 2590.220 ;
        RECT 2162.990 2590.360 2163.310 2590.420 ;
        RECT 2212.670 2590.360 2212.990 2590.420 ;
        RECT 2162.990 2590.220 2212.990 2590.360 ;
        RECT 2162.990 2590.160 2163.310 2590.220 ;
        RECT 2212.670 2590.160 2212.990 2590.220 ;
        RECT 1414.110 2590.020 1414.430 2590.080 ;
        RECT 1593.970 2590.020 1594.290 2590.080 ;
        RECT 1414.110 2589.880 1594.290 2590.020 ;
        RECT 1414.110 2589.820 1414.430 2589.880 ;
        RECT 1593.970 2589.820 1594.290 2589.880 ;
        RECT 1641.810 2590.020 1642.130 2590.080 ;
        RECT 1697.930 2590.020 1698.250 2590.080 ;
        RECT 1641.810 2589.880 1698.250 2590.020 ;
        RECT 1641.810 2589.820 1642.130 2589.880 ;
        RECT 1697.930 2589.820 1698.250 2589.880 ;
        RECT 1702.990 2590.020 1703.310 2590.080 ;
        RECT 2187.370 2590.020 2187.690 2590.080 ;
        RECT 1702.990 2589.880 2187.690 2590.020 ;
        RECT 1702.990 2589.820 1703.310 2589.880 ;
        RECT 2187.370 2589.820 2187.690 2589.880 ;
        RECT 2197.490 2590.020 2197.810 2590.080 ;
        RECT 2243.490 2590.020 2243.810 2590.080 ;
        RECT 2197.490 2589.880 2243.810 2590.020 ;
        RECT 2197.490 2589.820 2197.810 2589.880 ;
        RECT 2243.490 2589.820 2243.810 2589.880 ;
        RECT 1400.310 2589.680 1400.630 2589.740 ;
        RECT 1587.530 2589.680 1587.850 2589.740 ;
        RECT 1400.310 2589.540 1587.850 2589.680 ;
        RECT 1400.310 2589.480 1400.630 2589.540 ;
        RECT 1587.530 2589.480 1587.850 2589.540 ;
        RECT 1614.210 2589.680 1614.530 2589.740 ;
        RECT 1690.570 2589.680 1690.890 2589.740 ;
        RECT 1614.210 2589.540 1690.890 2589.680 ;
        RECT 1614.210 2589.480 1614.530 2589.540 ;
        RECT 1690.570 2589.480 1690.890 2589.540 ;
        RECT 1707.590 2589.680 1707.910 2589.740 ;
        RECT 2201.170 2589.680 2201.490 2589.740 ;
        RECT 1707.590 2589.540 2201.490 2589.680 ;
        RECT 1707.590 2589.480 1707.910 2589.540 ;
        RECT 2201.170 2589.480 2201.490 2589.540 ;
        RECT 2220.490 2589.680 2220.810 2589.740 ;
        RECT 2349.290 2589.680 2349.610 2589.740 ;
        RECT 2220.490 2589.540 2349.610 2589.680 ;
        RECT 2220.490 2589.480 2220.810 2589.540 ;
        RECT 2349.290 2589.480 2349.610 2589.540 ;
        RECT 1386.510 2589.340 1386.830 2589.400 ;
        RECT 1587.070 2589.340 1587.390 2589.400 ;
        RECT 1386.510 2589.200 1587.390 2589.340 ;
        RECT 1386.510 2589.140 1386.830 2589.200 ;
        RECT 1587.070 2589.140 1587.390 2589.200 ;
        RECT 1607.310 2589.340 1607.630 2589.400 ;
        RECT 1683.670 2589.340 1683.990 2589.400 ;
        RECT 1607.310 2589.200 1683.990 2589.340 ;
        RECT 1607.310 2589.140 1607.630 2589.200 ;
        RECT 1683.670 2589.140 1683.990 2589.200 ;
        RECT 1714.950 2589.340 1715.270 2589.400 ;
        RECT 2214.970 2589.340 2215.290 2589.400 ;
        RECT 1714.950 2589.200 2215.290 2589.340 ;
        RECT 1714.950 2589.140 1715.270 2589.200 ;
        RECT 2214.970 2589.140 2215.290 2589.200 ;
        RECT 2227.850 2589.340 2228.170 2589.400 ;
        RECT 2383.790 2589.340 2384.110 2589.400 ;
        RECT 2227.850 2589.200 2384.110 2589.340 ;
        RECT 2227.850 2589.140 2228.170 2589.200 ;
        RECT 2383.790 2589.140 2384.110 2589.200 ;
        RECT 1579.710 2589.000 1580.030 2589.060 ;
        RECT 1669.870 2589.000 1670.190 2589.060 ;
        RECT 1579.710 2588.860 1670.190 2589.000 ;
        RECT 1579.710 2588.800 1580.030 2588.860 ;
        RECT 1669.870 2588.800 1670.190 2588.860 ;
        RECT 1721.850 2589.000 1722.170 2589.060 ;
        RECT 2228.770 2589.000 2229.090 2589.060 ;
        RECT 1721.850 2588.860 2229.090 2589.000 ;
        RECT 1721.850 2588.800 1722.170 2588.860 ;
        RECT 2228.770 2588.800 2229.090 2588.860 ;
        RECT 1565.910 2588.660 1566.230 2588.720 ;
        RECT 1663.430 2588.660 1663.750 2588.720 ;
        RECT 1565.910 2588.520 1663.750 2588.660 ;
        RECT 1565.910 2588.460 1566.230 2588.520 ;
        RECT 1663.430 2588.460 1663.750 2588.520 ;
        RECT 1669.410 2588.660 1669.730 2588.720 ;
        RECT 1711.270 2588.660 1711.590 2588.720 ;
        RECT 1669.410 2588.520 1711.590 2588.660 ;
        RECT 1669.410 2588.460 1669.730 2588.520 ;
        RECT 1711.270 2588.460 1711.590 2588.520 ;
        RECT 1721.390 2588.660 1721.710 2588.720 ;
        RECT 1739.330 2588.660 1739.650 2588.720 ;
        RECT 1721.390 2588.520 1739.650 2588.660 ;
        RECT 1721.390 2588.460 1721.710 2588.520 ;
        RECT 1739.330 2588.460 1739.650 2588.520 ;
        RECT 2235.210 2588.660 2235.530 2588.720 ;
        RECT 2369.990 2588.660 2370.310 2588.720 ;
        RECT 2235.210 2588.520 2370.310 2588.660 ;
        RECT 2235.210 2588.460 2235.530 2588.520 ;
        RECT 2369.990 2588.460 2370.310 2588.520 ;
        RECT 1524.510 2588.320 1524.830 2588.380 ;
        RECT 1649.170 2588.320 1649.490 2588.380 ;
        RECT 1524.510 2588.180 1649.490 2588.320 ;
        RECT 1524.510 2588.120 1524.830 2588.180 ;
        RECT 1649.170 2588.120 1649.490 2588.180 ;
        RECT 1686.890 2588.320 1687.210 2588.380 ;
        RECT 1718.170 2588.320 1718.490 2588.380 ;
        RECT 1686.890 2588.180 1718.490 2588.320 ;
        RECT 1686.890 2588.120 1687.210 2588.180 ;
        RECT 1718.170 2588.120 1718.490 2588.180 ;
        RECT 2190.590 2588.320 2190.910 2588.380 ;
        RECT 2235.670 2588.320 2235.990 2588.380 ;
        RECT 2190.590 2588.180 2235.990 2588.320 ;
        RECT 2190.590 2588.120 2190.910 2588.180 ;
        RECT 2235.670 2588.120 2235.990 2588.180 ;
        RECT 2241.650 2588.320 2241.970 2588.380 ;
        RECT 2356.190 2588.320 2356.510 2588.380 ;
        RECT 2241.650 2588.180 2356.510 2588.320 ;
        RECT 2241.650 2588.120 2241.970 2588.180 ;
        RECT 2356.190 2588.120 2356.510 2588.180 ;
        RECT 1552.110 2587.980 1552.430 2588.040 ;
        RECT 1662.970 2587.980 1663.290 2588.040 ;
        RECT 1552.110 2587.840 1663.290 2587.980 ;
        RECT 1552.110 2587.780 1552.430 2587.840 ;
        RECT 1662.970 2587.780 1663.290 2587.840 ;
        RECT 1703.910 2587.980 1704.230 2588.040 ;
        RECT 1731.970 2587.980 1732.290 2588.040 ;
        RECT 1703.910 2587.840 1732.290 2587.980 ;
        RECT 1703.910 2587.780 1704.230 2587.840 ;
        RECT 1731.970 2587.780 1732.290 2587.840 ;
        RECT 2183.690 2587.980 2184.010 2588.040 ;
        RECT 2186.450 2587.980 2186.770 2588.040 ;
        RECT 2231.990 2587.980 2232.310 2588.040 ;
        RECT 2183.690 2587.840 2232.310 2587.980 ;
        RECT 2183.690 2587.780 2184.010 2587.840 ;
        RECT 2186.450 2587.780 2186.770 2587.840 ;
        RECT 2231.990 2587.780 2232.310 2587.840 ;
        RECT 1331.310 2587.640 1331.630 2587.700 ;
        RECT 1560.850 2587.640 1561.170 2587.700 ;
        RECT 1331.310 2587.500 1561.170 2587.640 ;
        RECT 1331.310 2587.440 1331.630 2587.500 ;
        RECT 1560.850 2587.440 1561.170 2587.500 ;
        RECT 1627.550 2587.640 1627.870 2587.700 ;
        RECT 1668.950 2587.640 1669.270 2587.700 ;
        RECT 1627.550 2587.500 1669.270 2587.640 ;
        RECT 1627.550 2587.440 1627.870 2587.500 ;
        RECT 1668.950 2587.440 1669.270 2587.500 ;
        RECT 1697.010 2587.640 1697.330 2587.700 ;
        RECT 1725.990 2587.640 1726.310 2587.700 ;
        RECT 1697.010 2587.500 1726.310 2587.640 ;
        RECT 1697.010 2587.440 1697.330 2587.500 ;
        RECT 1725.990 2587.440 1726.310 2587.500 ;
        RECT 1731.510 2587.640 1731.830 2587.700 ;
        RECT 1738.870 2587.640 1739.190 2587.700 ;
        RECT 1731.510 2587.500 1739.190 2587.640 ;
        RECT 1731.510 2587.440 1731.830 2587.500 ;
        RECT 1738.870 2587.440 1739.190 2587.500 ;
        RECT 2170.810 2587.640 2171.130 2587.700 ;
        RECT 2215.890 2587.640 2216.210 2587.700 ;
        RECT 2170.810 2587.500 2216.210 2587.640 ;
        RECT 2170.810 2587.440 2171.130 2587.500 ;
        RECT 2215.890 2587.440 2216.210 2587.500 ;
        RECT 2227.390 2587.640 2227.710 2587.700 ;
        RECT 2397.590 2587.640 2397.910 2587.700 ;
        RECT 2227.390 2587.500 2397.910 2587.640 ;
        RECT 2227.390 2587.440 2227.710 2587.500 ;
        RECT 2397.590 2587.440 2397.910 2587.500 ;
        RECT 1898.030 2570.300 1898.350 2570.360 ;
        RECT 1898.950 2570.300 1899.270 2570.360 ;
        RECT 1898.030 2570.160 1899.270 2570.300 ;
        RECT 1898.030 2570.100 1898.350 2570.160 ;
        RECT 1898.950 2570.100 1899.270 2570.160 ;
        RECT 2170.350 2560.100 2170.670 2560.160 ;
        RECT 2170.810 2560.100 2171.130 2560.160 ;
        RECT 2170.350 2559.960 2171.130 2560.100 ;
        RECT 2170.350 2559.900 2170.670 2559.960 ;
        RECT 2170.810 2559.900 2171.130 2559.960 ;
        RECT 1898.030 2497.880 1898.350 2497.940 ;
        RECT 1898.950 2497.880 1899.270 2497.940 ;
        RECT 1898.030 2497.740 1899.270 2497.880 ;
        RECT 1898.030 2497.680 1898.350 2497.740 ;
        RECT 1898.950 2497.680 1899.270 2497.740 ;
        RECT 1898.030 2473.740 1898.350 2473.800 ;
        RECT 1898.950 2473.740 1899.270 2473.800 ;
        RECT 1898.030 2473.600 1899.270 2473.740 ;
        RECT 1898.030 2473.540 1898.350 2473.600 ;
        RECT 1898.950 2473.540 1899.270 2473.600 ;
        RECT 2168.050 2463.200 2168.370 2463.260 ;
        RECT 2169.430 2463.200 2169.750 2463.260 ;
        RECT 2168.050 2463.060 2169.750 2463.200 ;
        RECT 2168.050 2463.000 2168.370 2463.060 ;
        RECT 2169.430 2463.000 2169.750 2463.060 ;
        RECT 1408.590 2414.920 1408.910 2414.980 ;
        RECT 1414.110 2414.920 1414.430 2414.980 ;
        RECT 1408.590 2414.780 1414.430 2414.920 ;
        RECT 1408.590 2414.720 1408.910 2414.780 ;
        RECT 1414.110 2414.720 1414.430 2414.780 ;
        RECT 1559.010 2414.920 1559.330 2414.980 ;
        RECT 1832.250 2414.920 1832.570 2414.980 ;
        RECT 1559.010 2414.780 1832.570 2414.920 ;
        RECT 1559.010 2414.720 1559.330 2414.780 ;
        RECT 1832.250 2414.720 1832.570 2414.780 ;
        RECT 1858.010 2414.920 1858.330 2414.980 ;
        RECT 2087.550 2414.920 2087.870 2414.980 ;
        RECT 1858.010 2414.780 2087.870 2414.920 ;
        RECT 1858.010 2414.720 1858.330 2414.780 ;
        RECT 2087.550 2414.720 2087.870 2414.780 ;
        RECT 2165.750 2414.920 2166.070 2414.980 ;
        RECT 2197.490 2414.920 2197.810 2414.980 ;
        RECT 2165.750 2414.780 2197.810 2414.920 ;
        RECT 2165.750 2414.720 2166.070 2414.780 ;
        RECT 2197.490 2414.720 2197.810 2414.780 ;
        RECT 2276.610 2414.920 2276.930 2414.980 ;
        RECT 2538.810 2414.920 2539.130 2414.980 ;
        RECT 2276.610 2414.780 2539.130 2414.920 ;
        RECT 2276.610 2414.720 2276.930 2414.780 ;
        RECT 2538.810 2414.720 2539.130 2414.780 ;
        RECT 1537.850 2414.580 1538.170 2414.640 ;
        RECT 1934.830 2414.580 1935.150 2414.640 ;
        RECT 1938.510 2414.580 1938.830 2414.640 ;
        RECT 1537.850 2414.440 1933.220 2414.580 ;
        RECT 1537.850 2414.380 1538.170 2414.440 ;
        RECT 1487.250 2414.240 1487.570 2414.300 ;
        RECT 1932.530 2414.240 1932.850 2414.300 ;
        RECT 1487.250 2414.100 1932.850 2414.240 ;
        RECT 1933.080 2414.240 1933.220 2414.440 ;
        RECT 1934.830 2414.440 1938.830 2414.580 ;
        RECT 1934.830 2414.380 1935.150 2414.440 ;
        RECT 1938.510 2414.380 1938.830 2414.440 ;
        RECT 2269.710 2414.580 2270.030 2414.640 ;
        RECT 2525.930 2414.580 2526.250 2414.640 ;
        RECT 2269.710 2414.440 2526.250 2414.580 ;
        RECT 2269.710 2414.380 2270.030 2414.440 ;
        RECT 2525.930 2414.380 2526.250 2414.440 ;
        RECT 1947.710 2414.240 1948.030 2414.300 ;
        RECT 1933.080 2414.100 1948.030 2414.240 ;
        RECT 1487.250 2414.040 1487.570 2414.100 ;
        RECT 1932.530 2414.040 1932.850 2414.100 ;
        RECT 1947.710 2414.040 1948.030 2414.100 ;
        RECT 2283.510 2414.240 2283.830 2414.300 ;
        RECT 2551.230 2414.240 2551.550 2414.300 ;
        RECT 2283.510 2414.100 2551.550 2414.240 ;
        RECT 2283.510 2414.040 2283.830 2414.100 ;
        RECT 2551.230 2414.040 2551.550 2414.100 ;
        RECT 1487.710 2413.900 1488.030 2413.960 ;
        RECT 1973.470 2413.900 1973.790 2413.960 ;
        RECT 1487.710 2413.760 1973.790 2413.900 ;
        RECT 1487.710 2413.700 1488.030 2413.760 ;
        RECT 1973.470 2413.700 1973.790 2413.760 ;
        RECT 2153.330 2413.900 2153.650 2413.960 ;
        RECT 2190.590 2413.900 2190.910 2413.960 ;
        RECT 2153.330 2413.760 2190.910 2413.900 ;
        RECT 2153.330 2413.700 2153.650 2413.760 ;
        RECT 2190.590 2413.700 2190.910 2413.760 ;
        RECT 2290.410 2413.900 2290.730 2413.960 ;
        RECT 2564.110 2413.900 2564.430 2413.960 ;
        RECT 2290.410 2413.760 2564.430 2413.900 ;
        RECT 2290.410 2413.700 2290.730 2413.760 ;
        RECT 2564.110 2413.700 2564.430 2413.760 ;
        RECT 1421.470 2413.560 1421.790 2413.620 ;
        RECT 1427.910 2413.560 1428.230 2413.620 ;
        RECT 1421.470 2413.420 1428.230 2413.560 ;
        RECT 1421.470 2413.360 1421.790 2413.420 ;
        RECT 1427.910 2413.360 1428.230 2413.420 ;
        RECT 1488.170 2413.560 1488.490 2413.620 ;
        RECT 1986.350 2413.560 1986.670 2413.620 ;
        RECT 1488.170 2413.420 1986.670 2413.560 ;
        RECT 1488.170 2413.360 1488.490 2413.420 ;
        RECT 1986.350 2413.360 1986.670 2413.420 ;
        RECT 2140.450 2413.560 2140.770 2413.620 ;
        RECT 2183.690 2413.560 2184.010 2413.620 ;
        RECT 2140.450 2413.420 2184.010 2413.560 ;
        RECT 2140.450 2413.360 2140.770 2413.420 ;
        RECT 2183.690 2413.360 2184.010 2413.420 ;
        RECT 2297.310 2413.560 2297.630 2413.620 ;
        RECT 2576.990 2413.560 2577.310 2413.620 ;
        RECT 2297.310 2413.420 2577.310 2413.560 ;
        RECT 2297.310 2413.360 2297.630 2413.420 ;
        RECT 2576.990 2413.360 2577.310 2413.420 ;
        RECT 1488.630 2413.220 1488.950 2413.280 ;
        RECT 1999.230 2413.220 1999.550 2413.280 ;
        RECT 1488.630 2413.080 1999.550 2413.220 ;
        RECT 1488.630 2413.020 1488.950 2413.080 ;
        RECT 1999.230 2413.020 1999.550 2413.080 ;
        RECT 2127.570 2413.220 2127.890 2413.280 ;
        RECT 2184.610 2413.220 2184.930 2413.280 ;
        RECT 2127.570 2413.080 2184.930 2413.220 ;
        RECT 2127.570 2413.020 2127.890 2413.080 ;
        RECT 2184.610 2413.020 2184.930 2413.080 ;
        RECT 2304.210 2413.220 2304.530 2413.280 ;
        RECT 2589.870 2413.220 2590.190 2413.280 ;
        RECT 2304.210 2413.080 2590.190 2413.220 ;
        RECT 2304.210 2413.020 2304.530 2413.080 ;
        RECT 2589.870 2413.020 2590.190 2413.080 ;
        RECT 1395.710 2412.880 1396.030 2412.940 ;
        RECT 1400.310 2412.880 1400.630 2412.940 ;
        RECT 1395.710 2412.740 1400.630 2412.880 ;
        RECT 1395.710 2412.680 1396.030 2412.740 ;
        RECT 1400.310 2412.680 1400.630 2412.740 ;
        RECT 1489.090 2412.880 1489.410 2412.940 ;
        RECT 2012.110 2412.880 2012.430 2412.940 ;
        RECT 1489.090 2412.740 2012.430 2412.880 ;
        RECT 1489.090 2412.680 1489.410 2412.740 ;
        RECT 2012.110 2412.680 2012.430 2412.740 ;
        RECT 2063.630 2412.880 2063.950 2412.940 ;
        RECT 2069.610 2412.880 2069.930 2412.940 ;
        RECT 2063.630 2412.740 2069.930 2412.880 ;
        RECT 2063.630 2412.680 2063.950 2412.740 ;
        RECT 2069.610 2412.680 2069.930 2412.740 ;
        RECT 2114.690 2412.880 2115.010 2412.940 ;
        RECT 2176.790 2412.880 2177.110 2412.940 ;
        RECT 2114.690 2412.740 2177.110 2412.880 ;
        RECT 2114.690 2412.680 2115.010 2412.740 ;
        RECT 2176.790 2412.680 2177.110 2412.740 ;
        RECT 2303.750 2412.880 2304.070 2412.940 ;
        RECT 2602.750 2412.880 2603.070 2412.940 ;
        RECT 2303.750 2412.740 2603.070 2412.880 ;
        RECT 2303.750 2412.680 2304.070 2412.740 ;
        RECT 2602.750 2412.680 2603.070 2412.740 ;
        RECT 1489.550 2412.540 1489.870 2412.600 ;
        RECT 2024.990 2412.540 2025.310 2412.600 ;
        RECT 1489.550 2412.400 2025.310 2412.540 ;
        RECT 1489.550 2412.340 1489.870 2412.400 ;
        RECT 2024.990 2412.340 2025.310 2412.400 ;
        RECT 2166.210 2412.540 2166.530 2412.600 ;
        RECT 2294.550 2412.540 2294.870 2412.600 ;
        RECT 2166.210 2412.400 2294.870 2412.540 ;
        RECT 2166.210 2412.340 2166.530 2412.400 ;
        RECT 2294.550 2412.340 2294.870 2412.400 ;
        RECT 2318.010 2412.540 2318.330 2412.600 ;
        RECT 2628.510 2412.540 2628.830 2412.600 ;
        RECT 2318.010 2412.400 2628.830 2412.540 ;
        RECT 2318.010 2412.340 2318.330 2412.400 ;
        RECT 2628.510 2412.340 2628.830 2412.400 ;
        RECT 1490.010 2412.200 1490.330 2412.260 ;
        RECT 2037.870 2412.200 2038.190 2412.260 ;
        RECT 1490.010 2412.060 2038.190 2412.200 ;
        RECT 1490.010 2412.000 1490.330 2412.060 ;
        RECT 2037.870 2412.000 2038.190 2412.060 ;
        RECT 2173.110 2412.200 2173.430 2412.260 ;
        RECT 2307.430 2412.200 2307.750 2412.260 ;
        RECT 2173.110 2412.060 2307.750 2412.200 ;
        RECT 2173.110 2412.000 2173.430 2412.060 ;
        RECT 2307.430 2412.000 2307.750 2412.060 ;
        RECT 2311.110 2412.200 2311.430 2412.260 ;
        RECT 2615.630 2412.200 2615.950 2412.260 ;
        RECT 2311.110 2412.060 2615.950 2412.200 ;
        RECT 2311.110 2412.000 2311.430 2412.060 ;
        RECT 2615.630 2412.000 2615.950 2412.060 ;
        RECT 1486.790 2411.860 1487.110 2411.920 ;
        RECT 2076.510 2411.860 2076.830 2411.920 ;
        RECT 1486.790 2411.720 2076.830 2411.860 ;
        RECT 1486.790 2411.660 1487.110 2411.720 ;
        RECT 2076.510 2411.660 2076.830 2411.720 ;
        RECT 2101.810 2411.860 2102.130 2411.920 ;
        RECT 2168.970 2411.860 2169.290 2411.920 ;
        RECT 2101.810 2411.720 2169.290 2411.860 ;
        RECT 2101.810 2411.660 2102.130 2411.720 ;
        RECT 2168.970 2411.660 2169.290 2411.720 ;
        RECT 2180.010 2411.860 2180.330 2411.920 ;
        RECT 2320.310 2411.860 2320.630 2411.920 ;
        RECT 2180.010 2411.720 2320.630 2411.860 ;
        RECT 2180.010 2411.660 2180.330 2411.720 ;
        RECT 2320.310 2411.660 2320.630 2411.720 ;
        RECT 2324.910 2411.860 2325.230 2411.920 ;
        RECT 2641.390 2411.860 2641.710 2411.920 ;
        RECT 2324.910 2411.720 2641.710 2411.860 ;
        RECT 2324.910 2411.660 2325.230 2411.720 ;
        RECT 2641.390 2411.660 2641.710 2411.720 ;
        RECT 1306.010 2411.520 1306.330 2411.580 ;
        RECT 1883.770 2411.520 1884.090 2411.580 ;
        RECT 1890.210 2411.520 1890.530 2411.580 ;
        RECT 1306.010 2411.380 1870.660 2411.520 ;
        RECT 1306.010 2411.320 1306.330 2411.380 ;
        RECT 1551.650 2411.180 1551.970 2411.240 ;
        RECT 1819.370 2411.180 1819.690 2411.240 ;
        RECT 1551.650 2411.040 1819.690 2411.180 ;
        RECT 1551.650 2410.980 1551.970 2411.040 ;
        RECT 1819.370 2410.980 1819.690 2411.040 ;
        RECT 1551.190 2410.840 1551.510 2410.900 ;
        RECT 1806.490 2410.840 1806.810 2410.900 ;
        RECT 1551.190 2410.700 1806.810 2410.840 ;
        RECT 1551.190 2410.640 1551.510 2410.700 ;
        RECT 1806.490 2410.640 1806.810 2410.700 ;
        RECT 1545.210 2410.500 1545.530 2410.560 ;
        RECT 1793.610 2410.500 1793.930 2410.560 ;
        RECT 1545.210 2410.360 1793.930 2410.500 ;
        RECT 1870.520 2410.500 1870.660 2411.380 ;
        RECT 1883.770 2411.380 1890.530 2411.520 ;
        RECT 1883.770 2411.320 1884.090 2411.380 ;
        RECT 1890.210 2411.320 1890.530 2411.380 ;
        RECT 1932.530 2411.520 1932.850 2411.580 ;
        RECT 1960.590 2411.520 1960.910 2411.580 ;
        RECT 1932.530 2411.380 1960.910 2411.520 ;
        RECT 1932.530 2411.320 1932.850 2411.380 ;
        RECT 1960.590 2411.320 1960.910 2411.380 ;
        RECT 2088.930 2411.520 2089.250 2411.580 ;
        RECT 2162.990 2411.520 2163.310 2411.580 ;
        RECT 2088.930 2411.380 2163.310 2411.520 ;
        RECT 2088.930 2411.320 2089.250 2411.380 ;
        RECT 2162.990 2411.320 2163.310 2411.380 ;
        RECT 2186.910 2411.520 2187.230 2411.580 ;
        RECT 2333.190 2411.520 2333.510 2411.580 ;
        RECT 2186.910 2411.380 2333.510 2411.520 ;
        RECT 2186.910 2411.320 2187.230 2411.380 ;
        RECT 2333.190 2411.320 2333.510 2411.380 ;
        RECT 2338.710 2411.520 2339.030 2411.580 ;
        RECT 2667.150 2411.520 2667.470 2411.580 ;
        RECT 2338.710 2411.380 2667.470 2411.520 ;
        RECT 2338.710 2411.320 2339.030 2411.380 ;
        RECT 2667.150 2411.320 2667.470 2411.380 ;
        RECT 1870.890 2411.180 1871.210 2411.240 ;
        RECT 2087.090 2411.180 2087.410 2411.240 ;
        RECT 1870.890 2411.040 2087.410 2411.180 ;
        RECT 1870.890 2410.980 1871.210 2411.040 ;
        RECT 2087.090 2410.980 2087.410 2411.040 ;
        RECT 2269.250 2411.180 2269.570 2411.240 ;
        RECT 2513.050 2411.180 2513.370 2411.240 ;
        RECT 2269.250 2411.040 2513.370 2411.180 ;
        RECT 2269.250 2410.980 2269.570 2411.040 ;
        RECT 2513.050 2410.980 2513.370 2411.040 ;
        RECT 2179.090 2410.840 2179.410 2410.900 ;
        RECT 2204.390 2410.840 2204.710 2410.900 ;
        RECT 2179.090 2410.700 2204.710 2410.840 ;
        RECT 2179.090 2410.640 2179.410 2410.700 ;
        RECT 2204.390 2410.640 2204.710 2410.700 ;
        RECT 2262.810 2410.840 2263.130 2410.900 ;
        RECT 2500.170 2410.840 2500.490 2410.900 ;
        RECT 2262.810 2410.700 2500.490 2410.840 ;
        RECT 2262.810 2410.640 2263.130 2410.700 ;
        RECT 2500.170 2410.640 2500.490 2410.700 ;
        RECT 1898.950 2410.500 1899.270 2410.560 ;
        RECT 1870.520 2410.360 1899.270 2410.500 ;
        RECT 1545.210 2410.300 1545.530 2410.360 ;
        RECT 1793.610 2410.300 1793.930 2410.360 ;
        RECT 1898.950 2410.300 1899.270 2410.360 ;
        RECT 2255.910 2410.500 2256.230 2410.560 ;
        RECT 2487.290 2410.500 2487.610 2410.560 ;
        RECT 2255.910 2410.360 2487.610 2410.500 ;
        RECT 2255.910 2410.300 2256.230 2410.360 ;
        RECT 2487.290 2410.300 2487.610 2410.360 ;
        RECT 1382.830 2410.160 1383.150 2410.220 ;
        RECT 1386.510 2410.160 1386.830 2410.220 ;
        RECT 1382.830 2410.020 1386.830 2410.160 ;
        RECT 1382.830 2409.960 1383.150 2410.020 ;
        RECT 1386.510 2409.960 1386.830 2410.020 ;
        RECT 1460.110 2410.160 1460.430 2410.220 ;
        RECT 1600.870 2410.160 1601.190 2410.220 ;
        RECT 1460.110 2410.020 1601.190 2410.160 ;
        RECT 1460.110 2409.960 1460.430 2410.020 ;
        RECT 1600.870 2409.960 1601.190 2410.020 ;
        RECT 1601.330 2410.160 1601.650 2410.220 ;
        RECT 1607.310 2410.160 1607.630 2410.220 ;
        RECT 1601.330 2410.020 1607.630 2410.160 ;
        RECT 1601.330 2409.960 1601.650 2410.020 ;
        RECT 1607.310 2409.960 1607.630 2410.020 ;
        RECT 1607.770 2410.160 1608.090 2410.220 ;
        RECT 1622.490 2410.160 1622.810 2410.220 ;
        RECT 1607.770 2410.020 1622.810 2410.160 ;
        RECT 1607.770 2409.960 1608.090 2410.020 ;
        RECT 1622.490 2409.960 1622.810 2410.020 ;
        RECT 1665.270 2410.160 1665.590 2410.220 ;
        RECT 1669.410 2410.160 1669.730 2410.220 ;
        RECT 1665.270 2410.020 1669.730 2410.160 ;
        RECT 1665.270 2409.960 1665.590 2410.020 ;
        RECT 1669.410 2409.960 1669.730 2410.020 ;
        RECT 1691.030 2410.160 1691.350 2410.220 ;
        RECT 1697.010 2410.160 1697.330 2410.220 ;
        RECT 1691.030 2410.020 1697.330 2410.160 ;
        RECT 1691.030 2409.960 1691.350 2410.020 ;
        RECT 1697.010 2409.960 1697.330 2410.020 ;
        RECT 1716.790 2410.160 1717.110 2410.220 ;
        RECT 1721.390 2410.160 1721.710 2410.220 ;
        RECT 1716.790 2410.020 1721.710 2410.160 ;
        RECT 1716.790 2409.960 1717.110 2410.020 ;
        RECT 1721.390 2409.960 1721.710 2410.020 ;
        RECT 1755.430 2410.160 1755.750 2410.220 ;
        RECT 1759.110 2410.160 1759.430 2410.220 ;
        RECT 1755.430 2410.020 1759.430 2410.160 ;
        RECT 1755.430 2409.960 1755.750 2410.020 ;
        RECT 1759.110 2409.960 1759.430 2410.020 ;
        RECT 1768.310 2410.160 1768.630 2410.220 ;
        RECT 1772.910 2410.160 1773.230 2410.220 ;
        RECT 1768.310 2410.020 1773.230 2410.160 ;
        RECT 1768.310 2409.960 1768.630 2410.020 ;
        RECT 1772.910 2409.960 1773.230 2410.020 ;
        RECT 2249.010 2410.160 2249.330 2410.220 ;
        RECT 2474.410 2410.160 2474.730 2410.220 ;
        RECT 2249.010 2410.020 2474.730 2410.160 ;
        RECT 2249.010 2409.960 2249.330 2410.020 ;
        RECT 2474.410 2409.960 2474.730 2410.020 ;
        RECT 1472.530 2409.820 1472.850 2409.880 ;
        RECT 1622.030 2409.820 1622.350 2409.880 ;
        RECT 1472.530 2409.680 1622.350 2409.820 ;
        RECT 1472.530 2409.620 1472.850 2409.680 ;
        RECT 1622.030 2409.620 1622.350 2409.680 ;
        RECT 1628.930 2409.820 1629.250 2409.880 ;
        RECT 2214.510 2409.820 2214.830 2409.880 ;
        RECT 2397.130 2409.820 2397.450 2409.880 ;
        RECT 1628.930 2409.680 1652.620 2409.820 ;
        RECT 1628.930 2409.620 1629.250 2409.680 ;
        RECT 1485.410 2409.480 1485.730 2409.540 ;
        RECT 1628.470 2409.480 1628.790 2409.540 ;
        RECT 1485.410 2409.340 1628.790 2409.480 ;
        RECT 1485.410 2409.280 1485.730 2409.340 ;
        RECT 1628.470 2409.280 1628.790 2409.340 ;
        RECT 1498.290 2409.140 1498.610 2409.200 ;
        RECT 1635.830 2409.140 1636.150 2409.200 ;
        RECT 1498.290 2409.000 1636.150 2409.140 ;
        RECT 1498.290 2408.940 1498.610 2409.000 ;
        RECT 1635.830 2408.940 1636.150 2409.000 ;
        RECT 1511.170 2408.800 1511.490 2408.860 ;
        RECT 1642.270 2408.800 1642.590 2408.860 ;
        RECT 1511.170 2408.660 1642.590 2408.800 ;
        RECT 1652.480 2408.800 1652.620 2409.680 ;
        RECT 2214.510 2409.680 2397.450 2409.820 ;
        RECT 2214.510 2409.620 2214.830 2409.680 ;
        RECT 2397.130 2409.620 2397.450 2409.680 ;
        RECT 2397.590 2409.820 2397.910 2409.880 ;
        RECT 2422.890 2409.820 2423.210 2409.880 ;
        RECT 2397.590 2409.680 2423.210 2409.820 ;
        RECT 2397.590 2409.620 2397.910 2409.680 ;
        RECT 2422.890 2409.620 2423.210 2409.680 ;
        RECT 1780.730 2409.480 1781.050 2409.540 ;
        RECT 1786.710 2409.480 1787.030 2409.540 ;
        RECT 1780.730 2409.340 1787.030 2409.480 ;
        RECT 1780.730 2409.280 1781.050 2409.340 ;
        RECT 1786.710 2409.280 1787.030 2409.340 ;
        RECT 2207.610 2409.480 2207.930 2409.540 ;
        RECT 2384.710 2409.480 2385.030 2409.540 ;
        RECT 2435.770 2409.480 2436.090 2409.540 ;
        RECT 2207.610 2409.340 2385.030 2409.480 ;
        RECT 2207.610 2409.280 2207.930 2409.340 ;
        RECT 2384.710 2409.280 2385.030 2409.340 ;
        RECT 2385.260 2409.340 2436.090 2409.480 ;
        RECT 2200.710 2409.140 2201.030 2409.200 ;
        RECT 2371.830 2409.140 2372.150 2409.200 ;
        RECT 2200.710 2409.000 2372.150 2409.140 ;
        RECT 2200.710 2408.940 2201.030 2409.000 ;
        RECT 2371.830 2408.940 2372.150 2409.000 ;
        RECT 2383.790 2409.140 2384.110 2409.200 ;
        RECT 2385.260 2409.140 2385.400 2409.340 ;
        RECT 2435.770 2409.280 2436.090 2409.340 ;
        RECT 2448.650 2409.140 2448.970 2409.200 ;
        RECT 2383.790 2409.000 2385.400 2409.140 ;
        RECT 2385.720 2409.000 2448.970 2409.140 ;
        RECT 2383.790 2408.940 2384.110 2409.000 ;
        RECT 1676.770 2408.800 1677.090 2408.860 ;
        RECT 1652.480 2408.660 1677.090 2408.800 ;
        RECT 1511.170 2408.600 1511.490 2408.660 ;
        RECT 1642.270 2408.600 1642.590 2408.660 ;
        RECT 1676.770 2408.600 1677.090 2408.660 ;
        RECT 1678.150 2408.800 1678.470 2408.860 ;
        RECT 1686.890 2408.800 1687.210 2408.860 ;
        RECT 1678.150 2408.660 1687.210 2408.800 ;
        RECT 1678.150 2408.600 1678.470 2408.660 ;
        RECT 1686.890 2408.600 1687.210 2408.660 ;
        RECT 2193.810 2408.800 2194.130 2408.860 ;
        RECT 2358.950 2408.800 2359.270 2408.860 ;
        RECT 2193.810 2408.660 2359.270 2408.800 ;
        RECT 2193.810 2408.600 2194.130 2408.660 ;
        RECT 2358.950 2408.600 2359.270 2408.660 ;
        RECT 2369.990 2408.800 2370.310 2408.860 ;
        RECT 2385.720 2408.800 2385.860 2409.000 ;
        RECT 2448.650 2408.940 2448.970 2409.000 ;
        RECT 2369.990 2408.660 2385.860 2408.800 ;
        RECT 2386.090 2408.800 2386.410 2408.860 ;
        RECT 2461.530 2408.800 2461.850 2408.860 ;
        RECT 2386.090 2408.660 2461.850 2408.800 ;
        RECT 2369.990 2408.600 2370.310 2408.660 ;
        RECT 2386.090 2408.600 2386.410 2408.660 ;
        RECT 2461.530 2408.600 2461.850 2408.660 ;
        RECT 1575.570 2408.460 1575.890 2408.520 ;
        RECT 1579.710 2408.460 1580.030 2408.520 ;
        RECT 1575.570 2408.320 1580.030 2408.460 ;
        RECT 1575.570 2408.260 1575.890 2408.320 ;
        RECT 1579.710 2408.260 1580.030 2408.320 ;
        RECT 1588.450 2408.460 1588.770 2408.520 ;
        RECT 1628.470 2408.460 1628.790 2408.520 ;
        RECT 1588.450 2408.320 1628.790 2408.460 ;
        RECT 1588.450 2408.260 1588.770 2408.320 ;
        RECT 1628.470 2408.260 1628.790 2408.320 ;
        RECT 2193.350 2408.460 2193.670 2408.520 ;
        RECT 2346.070 2408.460 2346.390 2408.520 ;
        RECT 2193.350 2408.320 2346.390 2408.460 ;
        RECT 2193.350 2408.260 2193.670 2408.320 ;
        RECT 2346.070 2408.260 2346.390 2408.320 ;
        RECT 2349.290 2408.460 2349.610 2408.520 ;
        RECT 2385.630 2408.460 2385.950 2408.520 ;
        RECT 2349.290 2408.320 2369.300 2408.460 ;
        RECT 2349.290 2408.260 2349.610 2408.320 ;
        RECT 2369.160 2407.780 2369.300 2408.320 ;
        RECT 2370.080 2408.320 2385.950 2408.460 ;
        RECT 2370.080 2407.780 2370.220 2408.320 ;
        RECT 2385.630 2408.260 2385.950 2408.320 ;
        RECT 2386.550 2408.460 2386.870 2408.520 ;
        RECT 2410.010 2408.460 2410.330 2408.520 ;
        RECT 2386.550 2408.320 2410.330 2408.460 ;
        RECT 2386.550 2408.260 2386.870 2408.320 ;
        RECT 2410.010 2408.260 2410.330 2408.320 ;
        RECT 2369.160 2407.640 2370.220 2407.780 ;
      LAYER met1 ;
        RECT 1305.520 1205.820 2694.260 2389.620 ;
      LAYER met1 ;
        RECT 1655.610 1193.640 1655.930 1193.700 ;
        RECT 1703.910 1193.640 1704.230 1193.700 ;
        RECT 1655.610 1193.500 1704.230 1193.640 ;
        RECT 1655.610 1193.440 1655.930 1193.500 ;
        RECT 1703.910 1193.440 1704.230 1193.500 ;
        RECT 2166.210 1193.640 2166.530 1193.700 ;
        RECT 2245.790 1193.640 2246.110 1193.700 ;
        RECT 2166.210 1193.500 2246.110 1193.640 ;
        RECT 2166.210 1193.440 2166.530 1193.500 ;
        RECT 2245.790 1193.440 2246.110 1193.500 ;
        RECT 2320.310 1193.640 2320.630 1193.700 ;
        RECT 2385.170 1193.640 2385.490 1193.700 ;
        RECT 2320.310 1193.500 2385.490 1193.640 ;
        RECT 2320.310 1193.440 2320.630 1193.500 ;
        RECT 2385.170 1193.440 2385.490 1193.500 ;
        RECT 2386.090 1193.640 2386.410 1193.700 ;
        RECT 2487.290 1193.640 2487.610 1193.700 ;
        RECT 2386.090 1193.500 2487.610 1193.640 ;
        RECT 2386.090 1193.440 2386.410 1193.500 ;
        RECT 2487.290 1193.440 2487.610 1193.500 ;
        RECT 1626.630 1193.300 1626.950 1193.360 ;
        RECT 1683.670 1193.300 1683.990 1193.360 ;
        RECT 1626.630 1193.160 1683.990 1193.300 ;
        RECT 1626.630 1193.100 1626.950 1193.160 ;
        RECT 1683.670 1193.100 1683.990 1193.160 ;
        RECT 1955.990 1193.300 1956.310 1193.360 ;
        RECT 2024.990 1193.300 2025.310 1193.360 ;
        RECT 1955.990 1193.160 2025.310 1193.300 ;
        RECT 1955.990 1193.100 1956.310 1193.160 ;
        RECT 2024.990 1193.100 2025.310 1193.160 ;
        RECT 2153.330 1193.300 2153.650 1193.360 ;
        RECT 2252.690 1193.300 2253.010 1193.360 ;
        RECT 2153.330 1193.160 2253.010 1193.300 ;
        RECT 2153.330 1193.100 2153.650 1193.160 ;
        RECT 2252.690 1193.100 2253.010 1193.160 ;
        RECT 2294.550 1193.300 2294.870 1193.360 ;
        RECT 2397.590 1193.300 2397.910 1193.360 ;
        RECT 2294.550 1193.160 2397.910 1193.300 ;
        RECT 2294.550 1193.100 2294.870 1193.160 ;
        RECT 2397.590 1193.100 2397.910 1193.160 ;
        RECT 1318.430 1192.960 1318.750 1193.020 ;
        RECT 1489.090 1192.960 1489.410 1193.020 ;
        RECT 1318.430 1192.820 1489.410 1192.960 ;
        RECT 1318.430 1192.760 1318.750 1192.820 ;
        RECT 1489.090 1192.760 1489.410 1192.820 ;
        RECT 1648.710 1192.960 1649.030 1193.020 ;
        RECT 1716.790 1192.960 1717.110 1193.020 ;
        RECT 1648.710 1192.820 1717.110 1192.960 ;
        RECT 1648.710 1192.760 1649.030 1192.820 ;
        RECT 1716.790 1192.760 1717.110 1192.820 ;
        RECT 1942.190 1192.960 1942.510 1193.020 ;
        RECT 2012.110 1192.960 2012.430 1193.020 ;
        RECT 1942.190 1192.820 2012.430 1192.960 ;
        RECT 1942.190 1192.760 1942.510 1192.820 ;
        RECT 2012.110 1192.760 2012.430 1192.820 ;
        RECT 2140.450 1192.960 2140.770 1193.020 ;
        RECT 2259.590 1192.960 2259.910 1193.020 ;
        RECT 2140.450 1192.820 2259.910 1192.960 ;
        RECT 2140.450 1192.760 2140.770 1192.820 ;
        RECT 2259.590 1192.760 2259.910 1192.820 ;
        RECT 2318.010 1192.960 2318.330 1193.020 ;
        RECT 2525.930 1192.960 2526.250 1193.020 ;
        RECT 2318.010 1192.820 2526.250 1192.960 ;
        RECT 2318.010 1192.760 2318.330 1192.820 ;
        RECT 2525.930 1192.760 2526.250 1192.820 ;
        RECT 1641.810 1192.620 1642.130 1192.680 ;
        RECT 1729.670 1192.620 1729.990 1192.680 ;
        RECT 1641.810 1192.480 1729.990 1192.620 ;
        RECT 1641.810 1192.420 1642.130 1192.480 ;
        RECT 1729.670 1192.420 1729.990 1192.480 ;
        RECT 1901.710 1192.620 1902.030 1192.680 ;
        RECT 1973.470 1192.620 1973.790 1192.680 ;
        RECT 1901.710 1192.480 1973.790 1192.620 ;
        RECT 1901.710 1192.420 1902.030 1192.480 ;
        RECT 1973.470 1192.420 1973.790 1192.480 ;
        RECT 2101.810 1192.620 2102.130 1192.680 ;
        RECT 2281.210 1192.620 2281.530 1192.680 ;
        RECT 2101.810 1192.480 2281.530 1192.620 ;
        RECT 2101.810 1192.420 2102.130 1192.480 ;
        RECT 2281.210 1192.420 2281.530 1192.480 ;
        RECT 2304.210 1192.620 2304.530 1192.680 ;
        RECT 2564.110 1192.620 2564.430 1192.680 ;
        RECT 2304.210 1192.480 2564.430 1192.620 ;
        RECT 2304.210 1192.420 2304.530 1192.480 ;
        RECT 2564.110 1192.420 2564.430 1192.480 ;
        RECT 1485.410 1192.280 1485.730 1192.340 ;
        RECT 1735.190 1192.280 1735.510 1192.340 ;
        RECT 1485.410 1192.140 1735.510 1192.280 ;
        RECT 1485.410 1192.080 1485.730 1192.140 ;
        RECT 1735.190 1192.080 1735.510 1192.140 ;
        RECT 1901.250 1192.280 1901.570 1192.340 ;
        RECT 1986.350 1192.280 1986.670 1192.340 ;
        RECT 1901.250 1192.140 1986.670 1192.280 ;
        RECT 1901.250 1192.080 1901.570 1192.140 ;
        RECT 1986.350 1192.080 1986.670 1192.140 ;
        RECT 2088.930 1192.280 2089.250 1192.340 ;
        RECT 2280.290 1192.280 2280.610 1192.340 ;
        RECT 2088.930 1192.140 2280.610 1192.280 ;
        RECT 2088.930 1192.080 2089.250 1192.140 ;
        RECT 2280.290 1192.080 2280.610 1192.140 ;
        RECT 2290.410 1192.280 2290.730 1192.340 ;
        RECT 2589.870 1192.280 2590.190 1192.340 ;
        RECT 2290.410 1192.140 2590.190 1192.280 ;
        RECT 2290.410 1192.080 2290.730 1192.140 ;
        RECT 2589.870 1192.080 2590.190 1192.140 ;
        RECT 1472.530 1191.940 1472.850 1192.000 ;
        RECT 1721.390 1191.940 1721.710 1192.000 ;
        RECT 1472.530 1191.800 1721.710 1191.940 ;
        RECT 1472.530 1191.740 1472.850 1191.800 ;
        RECT 1721.390 1191.740 1721.710 1191.800 ;
        RECT 1855.710 1191.940 1856.030 1192.000 ;
        RECT 1947.710 1191.940 1948.030 1192.000 ;
        RECT 1855.710 1191.800 1948.030 1191.940 ;
        RECT 1855.710 1191.740 1856.030 1191.800 ;
        RECT 1947.710 1191.740 1948.030 1191.800 ;
        RECT 1969.790 1191.940 1970.110 1192.000 ;
        RECT 2037.870 1191.940 2038.190 1192.000 ;
        RECT 1969.790 1191.800 2038.190 1191.940 ;
        RECT 1969.790 1191.740 1970.110 1191.800 ;
        RECT 2037.870 1191.740 2038.190 1191.800 ;
        RECT 2114.690 1191.940 2115.010 1192.000 ;
        RECT 2273.390 1191.940 2273.710 1192.000 ;
        RECT 2114.690 1191.800 2273.710 1191.940 ;
        RECT 2114.690 1191.740 2115.010 1191.800 ;
        RECT 2273.390 1191.740 2273.710 1191.800 ;
        RECT 2276.150 1191.940 2276.470 1192.000 ;
        RECT 2615.630 1191.940 2615.950 1192.000 ;
        RECT 2276.150 1191.800 2615.950 1191.940 ;
        RECT 2276.150 1191.740 2276.470 1191.800 ;
        RECT 2615.630 1191.740 2615.950 1191.800 ;
        RECT 1447.230 1191.600 1447.550 1191.660 ;
        RECT 1707.590 1191.600 1707.910 1191.660 ;
        RECT 1447.230 1191.460 1707.910 1191.600 ;
        RECT 1447.230 1191.400 1447.550 1191.460 ;
        RECT 1707.590 1191.400 1707.910 1191.460 ;
        RECT 1902.170 1191.600 1902.490 1191.660 ;
        RECT 2076.510 1191.600 2076.830 1191.660 ;
        RECT 1902.170 1191.460 2076.830 1191.600 ;
        RECT 1902.170 1191.400 1902.490 1191.460 ;
        RECT 2076.510 1191.400 2076.830 1191.460 ;
        RECT 2127.570 1191.600 2127.890 1191.660 ;
        RECT 2266.490 1191.600 2266.810 1191.660 ;
        RECT 2127.570 1191.460 2266.810 1191.600 ;
        RECT 2127.570 1191.400 2127.890 1191.460 ;
        RECT 2266.490 1191.400 2266.810 1191.460 ;
        RECT 2269.710 1191.600 2270.030 1191.660 ;
        RECT 2641.390 1191.600 2641.710 1191.660 ;
        RECT 2269.710 1191.460 2641.710 1191.600 ;
        RECT 2269.710 1191.400 2270.030 1191.460 ;
        RECT 2641.390 1191.400 2641.710 1191.460 ;
        RECT 1421.470 1191.260 1421.790 1191.320 ;
        RECT 1693.790 1191.260 1694.110 1191.320 ;
        RECT 1421.470 1191.120 1694.110 1191.260 ;
        RECT 1421.470 1191.060 1421.790 1191.120 ;
        RECT 1693.790 1191.060 1694.110 1191.120 ;
        RECT 1922.410 1191.260 1922.730 1191.320 ;
        RECT 2238.890 1191.260 2239.210 1191.320 ;
        RECT 1922.410 1191.120 2239.210 1191.260 ;
        RECT 1922.410 1191.060 1922.730 1191.120 ;
        RECT 2238.890 1191.060 2239.210 1191.120 ;
        RECT 2255.910 1191.260 2256.230 1191.320 ;
        RECT 2667.150 1191.260 2667.470 1191.320 ;
        RECT 2255.910 1191.120 2667.470 1191.260 ;
        RECT 2255.910 1191.060 2256.230 1191.120 ;
        RECT 2667.150 1191.060 2667.470 1191.120 ;
        RECT 1434.350 1190.920 1434.670 1190.980 ;
        RECT 1700.690 1190.920 1701.010 1190.980 ;
        RECT 1434.350 1190.780 1701.010 1190.920 ;
        RECT 1434.350 1190.720 1434.670 1190.780 ;
        RECT 1700.690 1190.720 1701.010 1190.780 ;
        RECT 1900.790 1190.920 1901.110 1190.980 ;
        RECT 1999.230 1190.920 1999.550 1190.980 ;
        RECT 1900.790 1190.780 1999.550 1190.920 ;
        RECT 1900.790 1190.720 1901.110 1190.780 ;
        RECT 1999.230 1190.720 1999.550 1190.780 ;
        RECT 2063.630 1190.920 2063.950 1190.980 ;
        RECT 2481.770 1190.920 2482.090 1190.980 ;
        RECT 2063.630 1190.780 2482.090 1190.920 ;
        RECT 2063.630 1190.720 2063.950 1190.780 ;
        RECT 2481.770 1190.720 2482.090 1190.780 ;
        RECT 1460.110 1190.580 1460.430 1190.640 ;
        RECT 1728.750 1190.580 1729.070 1190.640 ;
        RECT 1460.110 1190.440 1729.070 1190.580 ;
        RECT 1460.110 1190.380 1460.430 1190.440 ;
        RECT 1728.750 1190.380 1729.070 1190.440 ;
        RECT 1780.730 1190.580 1781.050 1190.640 ;
        RECT 2391.150 1190.580 2391.470 1190.640 ;
        RECT 1780.730 1190.440 2391.470 1190.580 ;
        RECT 1780.730 1190.380 1781.050 1190.440 ;
        RECT 2391.150 1190.380 2391.470 1190.440 ;
        RECT 1331.310 1190.240 1331.630 1190.300 ;
        RECT 1728.290 1190.240 1728.610 1190.300 ;
        RECT 1331.310 1190.100 1728.610 1190.240 ;
        RECT 1331.310 1190.040 1331.630 1190.100 ;
        RECT 1728.290 1190.040 1728.610 1190.100 ;
        RECT 1768.310 1190.240 1768.630 1190.300 ;
        RECT 2385.630 1190.240 2385.950 1190.300 ;
        RECT 1768.310 1190.100 2385.950 1190.240 ;
        RECT 1768.310 1190.040 1768.630 1190.100 ;
        RECT 2385.630 1190.040 2385.950 1190.100 ;
        RECT 2391.610 1190.240 2391.930 1190.300 ;
        RECT 2500.170 1190.240 2500.490 1190.300 ;
        RECT 2391.610 1190.100 2500.490 1190.240 ;
        RECT 2391.610 1190.040 2391.930 1190.100 ;
        RECT 2500.170 1190.040 2500.490 1190.100 ;
        RECT 2179.090 1189.900 2179.410 1189.960 ;
        RECT 2239.350 1189.900 2239.670 1189.960 ;
        RECT 2179.090 1189.760 2239.670 1189.900 ;
        RECT 2179.090 1189.700 2179.410 1189.760 ;
        RECT 2239.350 1189.700 2239.670 1189.760 ;
        RECT 2359.410 1189.900 2359.730 1189.960 ;
        RECT 2435.770 1189.900 2436.090 1189.960 ;
        RECT 2359.410 1189.760 2436.090 1189.900 ;
        RECT 2359.410 1189.700 2359.730 1189.760 ;
        RECT 2435.770 1189.700 2436.090 1189.760 ;
        RECT 2366.310 1189.560 2366.630 1189.620 ;
        RECT 2422.890 1189.560 2423.210 1189.620 ;
        RECT 2366.310 1189.420 2423.210 1189.560 ;
        RECT 2366.310 1189.360 2366.630 1189.420 ;
        RECT 2422.890 1189.360 2423.210 1189.420 ;
        RECT 2333.190 1189.220 2333.510 1189.280 ;
        RECT 2383.790 1189.220 2384.110 1189.280 ;
        RECT 2333.190 1189.080 2384.110 1189.220 ;
        RECT 2333.190 1189.020 2333.510 1189.080 ;
        RECT 2383.790 1189.020 2384.110 1189.080 ;
        RECT 2346.070 1188.880 2346.390 1188.940 ;
        RECT 2390.690 1188.880 2391.010 1188.940 ;
        RECT 2346.070 1188.740 2391.010 1188.880 ;
        RECT 2346.070 1188.680 2346.390 1188.740 ;
        RECT 2390.690 1188.680 2391.010 1188.740 ;
        RECT 2358.950 1188.200 2359.270 1188.260 ;
        RECT 2387.930 1188.200 2388.250 1188.260 ;
        RECT 2358.950 1188.060 2388.250 1188.200 ;
        RECT 2358.950 1188.000 2359.270 1188.060 ;
        RECT 2387.930 1188.000 2388.250 1188.060 ;
        RECT 1662.510 1187.860 1662.830 1187.920 ;
        RECT 1691.030 1187.860 1691.350 1187.920 ;
        RECT 1662.510 1187.720 1691.350 1187.860 ;
        RECT 1662.510 1187.660 1662.830 1187.720 ;
        RECT 1691.030 1187.660 1691.350 1187.720 ;
        RECT 2380.110 1187.860 2380.430 1187.920 ;
        RECT 2397.130 1187.860 2397.450 1187.920 ;
        RECT 2380.110 1187.720 2397.450 1187.860 ;
        RECT 2380.110 1187.660 2380.430 1187.720 ;
        RECT 2397.130 1187.660 2397.450 1187.720 ;
        RECT 1669.410 1187.520 1669.730 1187.580 ;
        RECT 1678.150 1187.520 1678.470 1187.580 ;
        RECT 1669.410 1187.380 1678.470 1187.520 ;
        RECT 1669.410 1187.320 1669.730 1187.380 ;
        RECT 1678.150 1187.320 1678.470 1187.380 ;
        RECT 2384.710 1187.520 2385.030 1187.580 ;
        RECT 2410.010 1187.520 2410.330 1187.580 ;
        RECT 2384.710 1187.380 2410.330 1187.520 ;
        RECT 2384.710 1187.320 2385.030 1187.380 ;
        RECT 2410.010 1187.320 2410.330 1187.380 ;
        RECT 1382.830 1187.180 1383.150 1187.240 ;
        RECT 1386.510 1187.180 1386.830 1187.240 ;
        RECT 1382.830 1187.040 1386.830 1187.180 ;
        RECT 1382.830 1186.980 1383.150 1187.040 ;
        RECT 1386.510 1186.980 1386.830 1187.040 ;
        RECT 1395.710 1187.180 1396.030 1187.240 ;
        RECT 1400.310 1187.180 1400.630 1187.240 ;
        RECT 1395.710 1187.040 1400.630 1187.180 ;
        RECT 1395.710 1186.980 1396.030 1187.040 ;
        RECT 1400.310 1186.980 1400.630 1187.040 ;
        RECT 1408.590 1187.180 1408.910 1187.240 ;
        RECT 1414.110 1187.180 1414.430 1187.240 ;
        RECT 1408.590 1187.040 1414.430 1187.180 ;
        RECT 1408.590 1186.980 1408.910 1187.040 ;
        RECT 1414.110 1186.980 1414.430 1187.040 ;
        RECT 1498.290 1187.180 1498.610 1187.240 ;
        RECT 1503.810 1187.180 1504.130 1187.240 ;
        RECT 1498.290 1187.040 1504.130 1187.180 ;
        RECT 1498.290 1186.980 1498.610 1187.040 ;
        RECT 1503.810 1186.980 1504.130 1187.040 ;
        RECT 1511.170 1187.180 1511.490 1187.240 ;
        RECT 1517.610 1187.180 1517.930 1187.240 ;
        RECT 1511.170 1187.040 1517.930 1187.180 ;
        RECT 1511.170 1186.980 1511.490 1187.040 ;
        RECT 1517.610 1186.980 1517.930 1187.040 ;
        RECT 1575.570 1187.180 1575.890 1187.240 ;
        RECT 1579.710 1187.180 1580.030 1187.240 ;
        RECT 1575.570 1187.040 1580.030 1187.180 ;
        RECT 1575.570 1186.980 1575.890 1187.040 ;
        RECT 1579.710 1186.980 1580.030 1187.040 ;
        RECT 1588.450 1187.180 1588.770 1187.240 ;
        RECT 1593.510 1187.180 1593.830 1187.240 ;
        RECT 1588.450 1187.040 1593.830 1187.180 ;
        RECT 1588.450 1186.980 1588.770 1187.040 ;
        RECT 1593.510 1186.980 1593.830 1187.040 ;
        RECT 1601.330 1187.180 1601.650 1187.240 ;
        RECT 1607.310 1187.180 1607.630 1187.240 ;
        RECT 1601.330 1187.040 1607.630 1187.180 ;
        RECT 1601.330 1186.980 1601.650 1187.040 ;
        RECT 1607.310 1186.980 1607.630 1187.040 ;
        RECT 1665.270 1187.180 1665.590 1187.240 ;
        RECT 1669.870 1187.180 1670.190 1187.240 ;
        RECT 1665.270 1187.040 1670.190 1187.180 ;
        RECT 1665.270 1186.980 1665.590 1187.040 ;
        RECT 1669.870 1186.980 1670.190 1187.040 ;
        RECT 1755.430 1187.180 1755.750 1187.240 ;
        RECT 1759.110 1187.180 1759.430 1187.240 ;
        RECT 1755.430 1187.040 1759.430 1187.180 ;
        RECT 1755.430 1186.980 1755.750 1187.040 ;
        RECT 1759.110 1186.980 1759.430 1187.040 ;
        RECT 1806.490 1187.180 1806.810 1187.240 ;
        RECT 1811.090 1187.180 1811.410 1187.240 ;
        RECT 1806.490 1187.040 1811.410 1187.180 ;
        RECT 1806.490 1186.980 1806.810 1187.040 ;
        RECT 1811.090 1186.980 1811.410 1187.040 ;
        RECT 1858.010 1187.180 1858.330 1187.240 ;
        RECT 1862.610 1187.180 1862.930 1187.240 ;
        RECT 1858.010 1187.040 1862.930 1187.180 ;
        RECT 1858.010 1186.980 1858.330 1187.040 ;
        RECT 1862.610 1186.980 1862.930 1187.040 ;
        RECT 1870.890 1187.180 1871.210 1187.240 ;
        RECT 1876.410 1187.180 1876.730 1187.240 ;
        RECT 1870.890 1187.040 1876.730 1187.180 ;
        RECT 1870.890 1186.980 1871.210 1187.040 ;
        RECT 1876.410 1186.980 1876.730 1187.040 ;
        RECT 1883.770 1187.180 1884.090 1187.240 ;
        RECT 1890.210 1187.180 1890.530 1187.240 ;
        RECT 1883.770 1187.040 1890.530 1187.180 ;
        RECT 1883.770 1186.980 1884.090 1187.040 ;
        RECT 1890.210 1186.980 1890.530 1187.040 ;
        RECT 1934.830 1187.180 1935.150 1187.240 ;
        RECT 1938.510 1187.180 1938.830 1187.240 ;
        RECT 1934.830 1187.040 1938.830 1187.180 ;
        RECT 1934.830 1186.980 1935.150 1187.040 ;
        RECT 1938.510 1186.980 1938.830 1187.040 ;
        RECT 2307.430 1187.180 2307.750 1187.240 ;
        RECT 2311.110 1187.180 2311.430 1187.240 ;
        RECT 2307.430 1187.040 2311.430 1187.180 ;
        RECT 2307.430 1186.980 2307.750 1187.040 ;
        RECT 2311.110 1186.980 2311.430 1187.040 ;
        RECT 2371.830 1187.180 2372.150 1187.240 ;
        RECT 2387.470 1187.180 2387.790 1187.240 ;
        RECT 2371.830 1187.040 2387.790 1187.180 ;
        RECT 2371.830 1186.980 2372.150 1187.040 ;
        RECT 2387.470 1186.980 2387.790 1187.040 ;
        RECT 2352.510 1026.020 2352.830 1026.080 ;
        RECT 2442.670 1026.020 2442.990 1026.080 ;
        RECT 2352.510 1025.880 2442.990 1026.020 ;
        RECT 2352.510 1025.820 2352.830 1025.880 ;
        RECT 2442.670 1025.820 2442.990 1025.880 ;
        RECT 2352.050 1025.340 2352.370 1025.400 ;
        RECT 2456.470 1025.340 2456.790 1025.400 ;
        RECT 2352.050 1025.200 2456.790 1025.340 ;
        RECT 2352.050 1025.140 2352.370 1025.200 ;
        RECT 2456.470 1025.140 2456.790 1025.200 ;
        RECT 2345.610 1025.000 2345.930 1025.060 ;
        RECT 2470.270 1025.000 2470.590 1025.060 ;
        RECT 2345.610 1024.860 2470.590 1025.000 ;
        RECT 2345.610 1024.800 2345.930 1024.860 ;
        RECT 2470.270 1024.800 2470.590 1024.860 ;
        RECT 1848.810 1024.660 1849.130 1024.720 ;
        RECT 2450.950 1024.660 2451.270 1024.720 ;
        RECT 1848.810 1024.520 2451.270 1024.660 ;
        RECT 1848.810 1024.460 1849.130 1024.520 ;
        RECT 2450.950 1024.460 2451.270 1024.520 ;
        RECT 2369.070 1022.280 2369.390 1022.340 ;
        RECT 2386.090 1022.280 2386.410 1022.340 ;
        RECT 2369.070 1022.140 2386.410 1022.280 ;
        RECT 2369.070 1022.080 2369.390 1022.140 ;
        RECT 2386.090 1022.080 2386.410 1022.140 ;
        RECT 1726.910 1021.600 1727.230 1021.660 ;
        RECT 1714.580 1021.460 1727.230 1021.600 ;
        RECT 1655.150 1021.260 1655.470 1021.320 ;
        RECT 1670.330 1021.260 1670.650 1021.320 ;
        RECT 1655.150 1021.120 1670.650 1021.260 ;
        RECT 1655.150 1021.060 1655.470 1021.120 ;
        RECT 1670.330 1021.060 1670.650 1021.120 ;
        RECT 1681.830 1021.260 1682.150 1021.320 ;
        RECT 1710.810 1021.260 1711.130 1021.320 ;
        RECT 1681.830 1021.120 1711.130 1021.260 ;
        RECT 1681.830 1021.060 1682.150 1021.120 ;
        RECT 1710.810 1021.060 1711.130 1021.120 ;
        RECT 1414.110 1020.920 1414.430 1020.980 ;
        RECT 1714.580 1020.920 1714.720 1021.460 ;
        RECT 1726.910 1021.400 1727.230 1021.460 ;
        RECT 1726.450 1021.260 1726.770 1021.320 ;
        RECT 1745.770 1021.260 1746.090 1021.320 ;
        RECT 1726.450 1021.120 1746.090 1021.260 ;
        RECT 1726.450 1021.060 1726.770 1021.120 ;
        RECT 1745.770 1021.060 1746.090 1021.120 ;
        RECT 1821.210 1021.260 1821.530 1021.320 ;
        RECT 1828.570 1021.260 1828.890 1021.320 ;
        RECT 1821.210 1021.120 1828.890 1021.260 ;
        RECT 1821.210 1021.060 1821.530 1021.120 ;
        RECT 1828.570 1021.060 1828.890 1021.120 ;
        RECT 2280.290 1021.260 2280.610 1021.320 ;
        RECT 2283.050 1021.260 2283.370 1021.320 ;
        RECT 2325.370 1021.260 2325.690 1021.320 ;
        RECT 2280.290 1021.120 2325.690 1021.260 ;
        RECT 2280.290 1021.060 2280.610 1021.120 ;
        RECT 2283.050 1021.060 2283.370 1021.120 ;
        RECT 2325.370 1021.060 2325.690 1021.120 ;
        RECT 2385.170 1021.260 2385.490 1021.320 ;
        RECT 2408.170 1021.260 2408.490 1021.320 ;
        RECT 2385.170 1021.120 2408.490 1021.260 ;
        RECT 2385.170 1021.060 2385.490 1021.120 ;
        RECT 2408.170 1021.060 2408.490 1021.120 ;
        RECT 1414.110 1020.780 1714.720 1020.920 ;
        RECT 1726.910 1020.920 1727.230 1020.980 ;
        RECT 1787.170 1020.920 1787.490 1020.980 ;
        RECT 1726.910 1020.780 1787.490 1020.920 ;
        RECT 1414.110 1020.720 1414.430 1020.780 ;
        RECT 1726.910 1020.720 1727.230 1020.780 ;
        RECT 1787.170 1020.720 1787.490 1020.780 ;
        RECT 1811.090 1020.920 1811.410 1020.980 ;
        RECT 1835.470 1020.920 1835.790 1020.980 ;
        RECT 1811.090 1020.780 1835.790 1020.920 ;
        RECT 1811.090 1020.720 1811.410 1020.780 ;
        RECT 1835.470 1020.720 1835.790 1020.780 ;
        RECT 2338.710 1020.920 2339.030 1020.980 ;
        RECT 2369.070 1020.920 2369.390 1020.980 ;
        RECT 2338.710 1020.780 2369.390 1020.920 ;
        RECT 2338.710 1020.720 2339.030 1020.780 ;
        RECT 2369.070 1020.720 2369.390 1020.780 ;
        RECT 2391.150 1020.920 2391.470 1020.980 ;
        RECT 2428.870 1020.920 2429.190 1020.980 ;
        RECT 2391.150 1020.780 2429.190 1020.920 ;
        RECT 2391.150 1020.720 2391.470 1020.780 ;
        RECT 2428.870 1020.720 2429.190 1020.780 ;
        RECT 1503.810 1020.580 1504.130 1020.640 ;
        RECT 1726.450 1020.580 1726.770 1020.640 ;
        RECT 1503.810 1020.440 1726.770 1020.580 ;
        RECT 1503.810 1020.380 1504.130 1020.440 ;
        RECT 1726.450 1020.380 1726.770 1020.440 ;
        RECT 1728.750 1020.580 1729.070 1020.640 ;
        RECT 1759.570 1020.580 1759.890 1020.640 ;
        RECT 1728.750 1020.440 1759.890 1020.580 ;
        RECT 1728.750 1020.380 1729.070 1020.440 ;
        RECT 1759.570 1020.380 1759.890 1020.440 ;
        RECT 2249.010 1020.580 2249.330 1020.640 ;
        RECT 2677.270 1020.580 2677.590 1020.640 ;
        RECT 2249.010 1020.440 2677.590 1020.580 ;
        RECT 2249.010 1020.380 2249.330 1020.440 ;
        RECT 2677.270 1020.380 2677.590 1020.440 ;
        RECT 1517.610 1020.240 1517.930 1020.300 ;
        RECT 1719.090 1020.240 1719.410 1020.300 ;
        RECT 1731.970 1020.240 1732.290 1020.300 ;
        RECT 1517.610 1020.100 1719.410 1020.240 ;
        RECT 1517.610 1020.040 1517.930 1020.100 ;
        RECT 1719.090 1020.040 1719.410 1020.100 ;
        RECT 1719.640 1020.100 1732.290 1020.240 ;
        RECT 1524.510 1019.900 1524.830 1019.960 ;
        RECT 1719.640 1019.900 1719.780 1020.100 ;
        RECT 1731.970 1020.040 1732.290 1020.100 ;
        RECT 1746.230 1020.240 1746.550 1020.300 ;
        RECT 1787.630 1020.240 1787.950 1020.300 ;
        RECT 1746.230 1020.100 1787.950 1020.240 ;
        RECT 1746.230 1020.040 1746.550 1020.100 ;
        RECT 1787.630 1020.040 1787.950 1020.100 ;
        RECT 1800.050 1020.240 1800.370 1020.300 ;
        RECT 2242.570 1020.240 2242.890 1020.300 ;
        RECT 1800.050 1020.100 2242.890 1020.240 ;
        RECT 1800.050 1020.040 1800.370 1020.100 ;
        RECT 2242.570 1020.040 2242.890 1020.100 ;
        RECT 2245.790 1020.240 2246.110 1020.300 ;
        RECT 2295.010 1020.240 2295.330 1020.300 ;
        RECT 2325.830 1020.240 2326.150 1020.300 ;
        RECT 2245.790 1020.100 2326.150 1020.240 ;
        RECT 2245.790 1020.040 2246.110 1020.100 ;
        RECT 2295.010 1020.040 2295.330 1020.100 ;
        RECT 2325.830 1020.040 2326.150 1020.100 ;
        RECT 2332.730 1020.240 2333.050 1020.300 ;
        RECT 2370.910 1020.240 2371.230 1020.300 ;
        RECT 2383.330 1020.240 2383.650 1020.300 ;
        RECT 2332.730 1020.100 2383.650 1020.240 ;
        RECT 2332.730 1020.040 2333.050 1020.100 ;
        RECT 2370.910 1020.040 2371.230 1020.100 ;
        RECT 2383.330 1020.040 2383.650 1020.100 ;
        RECT 2383.790 1020.240 2384.110 1020.300 ;
        RECT 2402.190 1020.240 2402.510 1020.300 ;
        RECT 2383.790 1020.100 2402.510 1020.240 ;
        RECT 2383.790 1020.040 2384.110 1020.100 ;
        RECT 2402.190 1020.040 2402.510 1020.100 ;
        RECT 1524.510 1019.760 1719.780 1019.900 ;
        RECT 1721.390 1019.900 1721.710 1019.960 ;
        RECT 1755.430 1019.900 1755.750 1019.960 ;
        RECT 1721.390 1019.760 1755.750 1019.900 ;
        RECT 1524.510 1019.700 1524.830 1019.760 ;
        RECT 1721.390 1019.700 1721.710 1019.760 ;
        RECT 1755.430 1019.700 1755.750 1019.760 ;
        RECT 1758.650 1019.900 1758.970 1019.960 ;
        RECT 1806.490 1019.900 1806.810 1019.960 ;
        RECT 2228.770 1019.900 2229.090 1019.960 ;
        RECT 1758.650 1019.760 2229.090 1019.900 ;
        RECT 1758.650 1019.700 1758.970 1019.760 ;
        RECT 1806.490 1019.700 1806.810 1019.760 ;
        RECT 2228.770 1019.700 2229.090 1019.760 ;
        RECT 2297.310 1019.900 2297.630 1019.960 ;
        RECT 2573.770 1019.900 2574.090 1019.960 ;
        RECT 2297.310 1019.760 2574.090 1019.900 ;
        RECT 2297.310 1019.700 2297.630 1019.760 ;
        RECT 2573.770 1019.700 2574.090 1019.760 ;
        RECT 1538.310 1019.560 1538.630 1019.620 ;
        RECT 1725.070 1019.560 1725.390 1019.620 ;
        RECT 1538.310 1019.420 1725.390 1019.560 ;
        RECT 1538.310 1019.360 1538.630 1019.420 ;
        RECT 1725.070 1019.360 1725.390 1019.420 ;
        RECT 1728.290 1019.560 1728.610 1019.620 ;
        RECT 1821.670 1019.560 1821.990 1019.620 ;
        RECT 1728.290 1019.420 1821.990 1019.560 ;
        RECT 1728.290 1019.360 1728.610 1019.420 ;
        RECT 1821.670 1019.360 1821.990 1019.420 ;
        RECT 2252.690 1019.560 2253.010 1019.620 ;
        RECT 2302.830 1019.560 2303.150 1019.620 ;
        RECT 2252.690 1019.420 2303.150 1019.560 ;
        RECT 2252.690 1019.360 2253.010 1019.420 ;
        RECT 2302.830 1019.360 2303.150 1019.420 ;
        RECT 2310.650 1019.560 2310.970 1019.620 ;
        RECT 2546.170 1019.560 2546.490 1019.620 ;
        RECT 2310.650 1019.420 2546.490 1019.560 ;
        RECT 2310.650 1019.360 2310.970 1019.420 ;
        RECT 2546.170 1019.360 2546.490 1019.420 ;
        RECT 1552.110 1019.220 1552.430 1019.280 ;
        RECT 1718.170 1019.220 1718.490 1019.280 ;
        RECT 1552.110 1019.080 1718.490 1019.220 ;
        RECT 1552.110 1019.020 1552.430 1019.080 ;
        RECT 1718.170 1019.020 1718.490 1019.080 ;
        RECT 1719.090 1019.220 1719.410 1019.280 ;
        RECT 1738.870 1019.220 1739.190 1019.280 ;
        RECT 1817.530 1019.220 1817.850 1019.280 ;
        RECT 2201.170 1019.220 2201.490 1019.280 ;
        RECT 1719.090 1019.080 1739.190 1019.220 ;
        RECT 1719.090 1019.020 1719.410 1019.080 ;
        RECT 1738.870 1019.020 1739.190 1019.080 ;
        RECT 1774.840 1019.080 2201.490 1019.220 ;
        RECT 1565.910 1018.880 1566.230 1018.940 ;
        RECT 1661.590 1018.880 1661.910 1018.940 ;
        RECT 1565.910 1018.740 1661.910 1018.880 ;
        RECT 1565.910 1018.680 1566.230 1018.740 ;
        RECT 1661.590 1018.680 1661.910 1018.740 ;
        RECT 1662.050 1018.880 1662.370 1018.940 ;
        RECT 1681.830 1018.880 1682.150 1018.940 ;
        RECT 1662.050 1018.740 1682.150 1018.880 ;
        RECT 1662.050 1018.680 1662.370 1018.740 ;
        RECT 1681.830 1018.680 1682.150 1018.740 ;
        RECT 1682.290 1018.880 1682.610 1018.940 ;
        RECT 1700.230 1018.880 1700.550 1018.940 ;
        RECT 1682.290 1018.740 1700.550 1018.880 ;
        RECT 1682.290 1018.680 1682.610 1018.740 ;
        RECT 1700.230 1018.680 1700.550 1018.740 ;
        RECT 1700.690 1018.880 1701.010 1018.940 ;
        RECT 1773.370 1018.880 1773.690 1018.940 ;
        RECT 1700.690 1018.740 1773.690 1018.880 ;
        RECT 1700.690 1018.680 1701.010 1018.740 ;
        RECT 1773.370 1018.680 1773.690 1018.740 ;
        RECT 1703.910 1018.540 1704.230 1018.600 ;
        RECT 1711.270 1018.540 1711.590 1018.600 ;
        RECT 1703.910 1018.400 1711.590 1018.540 ;
        RECT 1703.910 1018.340 1704.230 1018.400 ;
        RECT 1711.270 1018.340 1711.590 1018.400 ;
        RECT 1724.610 1018.540 1724.930 1018.600 ;
        RECT 1771.530 1018.540 1771.850 1018.600 ;
        RECT 1774.840 1018.540 1774.980 1019.080 ;
        RECT 1817.530 1019.020 1817.850 1019.080 ;
        RECT 2201.170 1019.020 2201.490 1019.080 ;
        RECT 2259.590 1019.220 2259.910 1019.280 ;
        RECT 2306.970 1019.220 2307.290 1019.280 ;
        RECT 2259.590 1019.080 2307.290 1019.220 ;
        RECT 2259.590 1019.020 2259.910 1019.080 ;
        RECT 2306.970 1019.020 2307.290 1019.080 ;
        RECT 2317.550 1019.220 2317.870 1019.280 ;
        RECT 2532.370 1019.220 2532.690 1019.280 ;
        RECT 2317.550 1019.080 2532.690 1019.220 ;
        RECT 2317.550 1019.020 2317.870 1019.080 ;
        RECT 2532.370 1019.020 2532.690 1019.080 ;
        RECT 1777.970 1018.880 1778.290 1018.940 ;
        RECT 1823.510 1018.880 1823.830 1018.940 ;
        RECT 2187.370 1018.880 2187.690 1018.940 ;
        RECT 1777.970 1018.740 2187.690 1018.880 ;
        RECT 1777.970 1018.680 1778.290 1018.740 ;
        RECT 1823.510 1018.680 1823.830 1018.740 ;
        RECT 2187.370 1018.680 2187.690 1018.740 ;
        RECT 2239.350 1018.880 2239.670 1018.940 ;
        RECT 2242.110 1018.880 2242.430 1018.940 ;
        RECT 2289.950 1018.880 2290.270 1018.940 ;
        RECT 2239.350 1018.740 2290.270 1018.880 ;
        RECT 2239.350 1018.680 2239.670 1018.740 ;
        RECT 2242.110 1018.680 2242.430 1018.740 ;
        RECT 2289.950 1018.680 2290.270 1018.740 ;
        RECT 2324.910 1018.880 2325.230 1018.940 ;
        RECT 2511.670 1018.880 2511.990 1018.940 ;
        RECT 2324.910 1018.740 2511.990 1018.880 ;
        RECT 2324.910 1018.680 2325.230 1018.740 ;
        RECT 2511.670 1018.680 2511.990 1018.740 ;
        RECT 1724.610 1018.400 1774.980 1018.540 ;
        RECT 2311.110 1018.540 2311.430 1018.600 ;
        RECT 2415.070 1018.540 2415.390 1018.600 ;
        RECT 2311.110 1018.400 2415.390 1018.540 ;
        RECT 1724.610 1018.340 1724.930 1018.400 ;
        RECT 1771.530 1018.340 1771.850 1018.400 ;
        RECT 2311.110 1018.340 2311.430 1018.400 ;
        RECT 2415.070 1018.340 2415.390 1018.400 ;
        RECT 1593.510 1018.200 1593.830 1018.260 ;
        RECT 1704.370 1018.200 1704.690 1018.260 ;
        RECT 1746.230 1018.200 1746.550 1018.260 ;
        RECT 1593.510 1018.060 1704.690 1018.200 ;
        RECT 1593.510 1018.000 1593.830 1018.060 ;
        RECT 1704.370 1018.000 1704.690 1018.060 ;
        RECT 1734.360 1018.060 1746.550 1018.200 ;
        RECT 1607.310 1017.860 1607.630 1017.920 ;
        RECT 1697.010 1017.860 1697.330 1017.920 ;
        RECT 1733.810 1017.860 1734.130 1017.920 ;
        RECT 1607.310 1017.720 1697.330 1017.860 ;
        RECT 1607.310 1017.660 1607.630 1017.720 ;
        RECT 1697.010 1017.660 1697.330 1017.720 ;
        RECT 1697.560 1017.720 1734.130 1017.860 ;
        RECT 1614.210 1017.520 1614.530 1017.580 ;
        RECT 1690.570 1017.520 1690.890 1017.580 ;
        RECT 1614.210 1017.380 1690.890 1017.520 ;
        RECT 1614.210 1017.320 1614.530 1017.380 ;
        RECT 1690.570 1017.320 1690.890 1017.380 ;
        RECT 1691.030 1017.520 1691.350 1017.580 ;
        RECT 1696.090 1017.520 1696.410 1017.580 ;
        RECT 1697.560 1017.520 1697.700 1017.720 ;
        RECT 1733.810 1017.660 1734.130 1017.720 ;
        RECT 1691.030 1017.380 1697.700 1017.520 ;
        RECT 1697.930 1017.520 1698.250 1017.580 ;
        RECT 1734.360 1017.520 1734.500 1018.060 ;
        RECT 1746.230 1018.000 1746.550 1018.060 ;
        RECT 1746.690 1018.200 1747.010 1018.260 ;
        RECT 1754.970 1018.200 1755.290 1018.260 ;
        RECT 1746.690 1018.060 1755.290 1018.200 ;
        RECT 1746.690 1018.000 1747.010 1018.060 ;
        RECT 1754.970 1018.000 1755.290 1018.060 ;
        RECT 1766.010 1018.200 1766.330 1018.260 ;
        RECT 1812.470 1018.200 1812.790 1018.260 ;
        RECT 2214.970 1018.200 2215.290 1018.260 ;
        RECT 1766.010 1018.060 2215.290 1018.200 ;
        RECT 1766.010 1018.000 1766.330 1018.060 ;
        RECT 1812.470 1018.000 1812.790 1018.060 ;
        RECT 2214.970 1018.000 2215.290 1018.060 ;
        RECT 2332.270 1018.200 2332.590 1018.260 ;
        RECT 2391.610 1018.200 2391.930 1018.260 ;
        RECT 2332.270 1018.060 2391.930 1018.200 ;
        RECT 2332.270 1018.000 2332.590 1018.060 ;
        RECT 2391.610 1018.000 2391.930 1018.060 ;
        RECT 2397.590 1018.200 2397.910 1018.260 ;
        RECT 2421.970 1018.200 2422.290 1018.260 ;
        RECT 2397.590 1018.060 2422.290 1018.200 ;
        RECT 2397.590 1018.000 2397.910 1018.060 ;
        RECT 2421.970 1018.000 2422.290 1018.060 ;
        RECT 1734.730 1017.860 1735.050 1017.920 ;
        RECT 1741.630 1017.860 1741.950 1017.920 ;
        RECT 1789.010 1017.860 1789.330 1017.920 ;
        RECT 2263.270 1017.860 2263.590 1017.920 ;
        RECT 1734.730 1017.720 2263.590 1017.860 ;
        RECT 1734.730 1017.660 1735.050 1017.720 ;
        RECT 1741.630 1017.660 1741.950 1017.720 ;
        RECT 1789.010 1017.660 1789.330 1017.720 ;
        RECT 2263.270 1017.660 2263.590 1017.720 ;
        RECT 2306.970 1017.860 2307.290 1017.920 ;
        RECT 2353.430 1017.860 2353.750 1017.920 ;
        RECT 2306.970 1017.720 2353.750 1017.860 ;
        RECT 2306.970 1017.660 2307.290 1017.720 ;
        RECT 2353.430 1017.660 2353.750 1017.720 ;
        RECT 1735.650 1017.520 1735.970 1017.580 ;
        RECT 2346.990 1017.520 2347.310 1017.580 ;
        RECT 2387.930 1017.520 2388.250 1017.580 ;
        RECT 1697.930 1017.380 1734.500 1017.520 ;
        RECT 1734.820 1017.380 1746.460 1017.520 ;
        RECT 1691.030 1017.320 1691.350 1017.380 ;
        RECT 1696.090 1017.320 1696.410 1017.380 ;
        RECT 1697.930 1017.320 1698.250 1017.380 ;
        RECT 1641.810 1017.180 1642.130 1017.240 ;
        RECT 1689.650 1017.180 1689.970 1017.240 ;
        RECT 1734.820 1017.180 1734.960 1017.380 ;
        RECT 1735.650 1017.320 1735.970 1017.380 ;
        RECT 1641.810 1017.040 1734.960 1017.180 ;
        RECT 1735.190 1017.180 1735.510 1017.240 ;
        RECT 1745.770 1017.180 1746.090 1017.240 ;
        RECT 1735.190 1017.040 1746.090 1017.180 ;
        RECT 1746.320 1017.180 1746.460 1017.380 ;
        RECT 2325.460 1017.380 2388.250 1017.520 ;
        RECT 1782.110 1017.180 1782.430 1017.240 ;
        RECT 2277.070 1017.180 2277.390 1017.240 ;
        RECT 1746.320 1017.040 2277.390 1017.180 ;
        RECT 1641.810 1016.980 1642.130 1017.040 ;
        RECT 1689.650 1016.980 1689.970 1017.040 ;
        RECT 1735.190 1016.980 1735.510 1017.040 ;
        RECT 1745.770 1016.980 1746.090 1017.040 ;
        RECT 1782.110 1016.980 1782.430 1017.040 ;
        RECT 2277.070 1016.980 2277.390 1017.040 ;
        RECT 2280.750 1017.180 2281.070 1017.240 ;
        RECT 2302.830 1017.180 2303.150 1017.240 ;
        RECT 2325.460 1017.180 2325.600 1017.380 ;
        RECT 2346.990 1017.320 2347.310 1017.380 ;
        RECT 2387.930 1017.320 2388.250 1017.380 ;
        RECT 2280.750 1017.040 2289.720 1017.180 ;
        RECT 2280.750 1016.980 2281.070 1017.040 ;
        RECT 1641.350 1016.840 1641.670 1016.900 ;
        RECT 1676.770 1016.840 1677.090 1016.900 ;
        RECT 1641.350 1016.700 1677.090 1016.840 ;
        RECT 1641.350 1016.640 1641.670 1016.700 ;
        RECT 1676.770 1016.640 1677.090 1016.700 ;
        RECT 1683.210 1016.840 1683.530 1016.900 ;
        RECT 1729.670 1016.840 1729.990 1016.900 ;
        RECT 1777.970 1016.840 1778.290 1016.900 ;
        RECT 1683.210 1016.700 1778.290 1016.840 ;
        RECT 1683.210 1016.640 1683.530 1016.700 ;
        RECT 1729.670 1016.640 1729.990 1016.700 ;
        RECT 1777.970 1016.640 1778.290 1016.700 ;
        RECT 1793.610 1016.840 1793.930 1016.900 ;
        RECT 1842.370 1016.840 1842.690 1016.900 ;
        RECT 1793.610 1016.700 1842.690 1016.840 ;
        RECT 1793.610 1016.640 1793.930 1016.700 ;
        RECT 1842.370 1016.640 1842.690 1016.700 ;
        RECT 1655.610 1016.500 1655.930 1016.560 ;
        RECT 1669.410 1016.500 1669.730 1016.560 ;
        RECT 1712.190 1016.500 1712.510 1016.560 ;
        RECT 1758.650 1016.500 1758.970 1016.560 ;
        RECT 1655.610 1016.360 1669.180 1016.500 ;
        RECT 1655.610 1016.300 1655.930 1016.360 ;
        RECT 1648.710 1016.160 1649.030 1016.220 ;
        RECT 1669.040 1016.160 1669.180 1016.360 ;
        RECT 1669.410 1016.360 1758.970 1016.500 ;
        RECT 1669.410 1016.300 1669.730 1016.360 ;
        RECT 1712.190 1016.300 1712.510 1016.360 ;
        RECT 1758.650 1016.300 1758.970 1016.360 ;
        RECT 1787.630 1016.500 1787.950 1016.560 ;
        RECT 1793.150 1016.500 1793.470 1016.560 ;
        RECT 2249.470 1016.500 2249.790 1016.560 ;
        RECT 1787.630 1016.360 2249.790 1016.500 ;
        RECT 2289.580 1016.500 2289.720 1017.040 ;
        RECT 2302.830 1017.040 2325.600 1017.180 ;
        RECT 2325.830 1017.180 2326.150 1017.240 ;
        RECT 2342.390 1017.180 2342.710 1017.240 ;
        RECT 2385.630 1017.180 2385.950 1017.240 ;
        RECT 2428.870 1017.180 2429.190 1017.240 ;
        RECT 2325.830 1017.040 2381.260 1017.180 ;
        RECT 2302.830 1016.980 2303.150 1017.040 ;
        RECT 2325.830 1016.980 2326.150 1017.040 ;
        RECT 2342.390 1016.980 2342.710 1017.040 ;
        RECT 2289.950 1016.840 2290.270 1016.900 ;
        RECT 2336.410 1016.840 2336.730 1016.900 ;
        RECT 2380.570 1016.840 2380.890 1016.900 ;
        RECT 2289.950 1016.700 2380.890 1016.840 ;
        RECT 2381.120 1016.840 2381.260 1017.040 ;
        RECT 2385.630 1017.040 2429.190 1017.180 ;
        RECT 2385.630 1016.980 2385.950 1017.040 ;
        RECT 2428.870 1016.980 2429.190 1017.040 ;
        RECT 2387.470 1016.840 2387.790 1016.900 ;
        RECT 2381.120 1016.700 2387.790 1016.840 ;
        RECT 2289.950 1016.640 2290.270 1016.700 ;
        RECT 2336.410 1016.640 2336.730 1016.700 ;
        RECT 2380.570 1016.640 2380.890 1016.700 ;
        RECT 2387.470 1016.640 2387.790 1016.700 ;
        RECT 2388.390 1016.840 2388.710 1016.900 ;
        RECT 2388.390 1016.700 2396.440 1016.840 ;
        RECT 2388.390 1016.640 2388.710 1016.700 ;
        RECT 2323.070 1016.500 2323.390 1016.560 ;
        RECT 2332.270 1016.500 2332.590 1016.560 ;
        RECT 2289.580 1016.360 2332.590 1016.500 ;
        RECT 1787.630 1016.300 1787.950 1016.360 ;
        RECT 1793.150 1016.300 1793.470 1016.360 ;
        RECT 2249.470 1016.300 2249.790 1016.360 ;
        RECT 2323.070 1016.300 2323.390 1016.360 ;
        RECT 2332.270 1016.300 2332.590 1016.360 ;
        RECT 2332.730 1016.500 2333.050 1016.560 ;
        RECT 2377.810 1016.500 2378.130 1016.560 ;
        RECT 2396.300 1016.500 2396.440 1016.700 ;
        RECT 2415.070 1016.500 2415.390 1016.560 ;
        RECT 2332.730 1016.360 2395.980 1016.500 ;
        RECT 2396.300 1016.360 2415.390 1016.500 ;
        RECT 2332.730 1016.300 2333.050 1016.360 ;
        RECT 2377.810 1016.300 2378.130 1016.360 ;
        RECT 1675.850 1016.160 1676.170 1016.220 ;
        RECT 1648.710 1016.020 1668.720 1016.160 ;
        RECT 1669.040 1016.020 1676.170 1016.160 ;
        RECT 1648.710 1015.960 1649.030 1016.020 ;
        RECT 1668.580 1015.820 1668.720 1016.020 ;
        RECT 1675.850 1015.960 1676.170 1016.020 ;
        RECT 1676.310 1016.160 1676.630 1016.220 ;
        RECT 1718.170 1016.160 1718.490 1016.220 ;
        RECT 1766.010 1016.160 1766.330 1016.220 ;
        RECT 2364.470 1016.160 2364.790 1016.220 ;
        RECT 2395.840 1016.160 2395.980 1016.360 ;
        RECT 2415.070 1016.300 2415.390 1016.360 ;
        RECT 2421.970 1016.160 2422.290 1016.220 ;
        RECT 1676.310 1016.020 1766.330 1016.160 ;
        RECT 1676.310 1015.960 1676.630 1016.020 ;
        RECT 1718.170 1015.960 1718.490 1016.020 ;
        RECT 1766.010 1015.960 1766.330 1016.020 ;
        RECT 2358.580 1016.020 2395.520 1016.160 ;
        RECT 2395.840 1016.020 2422.290 1016.160 ;
        RECT 1691.030 1015.820 1691.350 1015.880 ;
        RECT 1668.580 1015.680 1691.350 1015.820 ;
        RECT 1691.030 1015.620 1691.350 1015.680 ;
        RECT 1693.790 1015.820 1694.110 1015.880 ;
        RECT 1780.270 1015.820 1780.590 1015.880 ;
        RECT 1693.790 1015.680 1780.590 1015.820 ;
        RECT 1693.790 1015.620 1694.110 1015.680 ;
        RECT 1780.270 1015.620 1780.590 1015.680 ;
        RECT 2275.230 1015.820 2275.550 1015.880 ;
        RECT 2318.010 1015.820 2318.330 1015.880 ;
        RECT 2358.580 1015.820 2358.720 1016.020 ;
        RECT 2364.470 1015.960 2364.790 1016.020 ;
        RECT 2395.380 1015.820 2395.520 1016.020 ;
        RECT 2421.970 1015.960 2422.290 1016.020 ;
        RECT 2408.170 1015.820 2408.490 1015.880 ;
        RECT 2275.230 1015.680 2358.720 1015.820 ;
        RECT 2359.040 1015.680 2395.060 1015.820 ;
        RECT 2395.380 1015.680 2408.490 1015.820 ;
        RECT 2275.230 1015.620 2275.550 1015.680 ;
        RECT 2318.010 1015.620 2318.330 1015.680 ;
        RECT 2359.040 1015.540 2359.180 1015.680 ;
        RECT 1661.590 1015.480 1661.910 1015.540 ;
        RECT 1682.290 1015.480 1682.610 1015.540 ;
        RECT 1661.590 1015.340 1682.610 1015.480 ;
        RECT 1661.590 1015.280 1661.910 1015.340 ;
        RECT 1682.290 1015.280 1682.610 1015.340 ;
        RECT 1683.210 1015.480 1683.530 1015.540 ;
        RECT 1724.610 1015.480 1724.930 1015.540 ;
        RECT 1683.210 1015.340 1724.930 1015.480 ;
        RECT 1683.210 1015.280 1683.530 1015.340 ;
        RECT 1724.610 1015.280 1724.930 1015.340 ;
        RECT 1754.970 1015.480 1755.290 1015.540 ;
        RECT 1800.050 1015.480 1800.370 1015.540 ;
        RECT 1754.970 1015.340 1800.370 1015.480 ;
        RECT 1754.970 1015.280 1755.290 1015.340 ;
        RECT 1800.050 1015.280 1800.370 1015.340 ;
        RECT 2266.490 1015.480 2266.810 1015.540 ;
        RECT 2312.030 1015.480 2312.350 1015.540 ;
        RECT 2358.950 1015.480 2359.270 1015.540 ;
        RECT 2266.490 1015.340 2359.270 1015.480 ;
        RECT 2266.490 1015.280 2266.810 1015.340 ;
        RECT 2312.030 1015.280 2312.350 1015.340 ;
        RECT 2358.950 1015.280 2359.270 1015.340 ;
        RECT 2359.410 1015.480 2359.730 1015.540 ;
        RECT 2394.370 1015.480 2394.690 1015.540 ;
        RECT 2359.410 1015.340 2394.690 1015.480 ;
        RECT 2394.920 1015.480 2395.060 1015.680 ;
        RECT 2408.170 1015.620 2408.490 1015.680 ;
        RECT 2403.110 1015.480 2403.430 1015.540 ;
        RECT 2394.920 1015.340 2403.430 1015.480 ;
        RECT 2359.410 1015.280 2359.730 1015.340 ;
        RECT 2394.370 1015.280 2394.690 1015.340 ;
        RECT 2403.110 1015.280 2403.430 1015.340 ;
        RECT 1707.590 1015.140 1707.910 1015.200 ;
        RECT 1766.470 1015.140 1766.790 1015.200 ;
        RECT 1707.590 1015.000 1766.790 1015.140 ;
        RECT 1707.590 1014.940 1707.910 1015.000 ;
        RECT 1766.470 1014.940 1766.790 1015.000 ;
        RECT 2276.610 1015.140 2276.930 1015.200 ;
        RECT 2622.070 1015.140 2622.390 1015.200 ;
        RECT 2276.610 1015.000 2622.390 1015.140 ;
        RECT 2276.610 1014.940 2276.930 1015.000 ;
        RECT 2622.070 1014.940 2622.390 1015.000 ;
        RECT 1400.310 1014.800 1400.630 1014.860 ;
        RECT 1787.170 1014.800 1787.490 1014.860 ;
        RECT 1400.310 1014.660 1787.490 1014.800 ;
        RECT 1400.310 1014.600 1400.630 1014.660 ;
        RECT 1787.170 1014.600 1787.490 1014.660 ;
        RECT 2262.810 1014.800 2263.130 1014.860 ;
        RECT 2649.670 1014.800 2649.990 1014.860 ;
        RECT 2262.810 1014.660 2649.990 1014.800 ;
        RECT 2262.810 1014.600 2263.130 1014.660 ;
        RECT 2649.670 1014.600 2649.990 1014.660 ;
        RECT 1579.710 1014.460 1580.030 1014.520 ;
        RECT 1711.270 1014.460 1711.590 1014.520 ;
        RECT 1746.690 1014.460 1747.010 1014.520 ;
        RECT 1579.710 1014.320 1711.590 1014.460 ;
        RECT 1579.710 1014.260 1580.030 1014.320 ;
        RECT 1711.270 1014.260 1711.590 1014.320 ;
        RECT 1711.820 1014.320 1747.010 1014.460 ;
        RECT 1710.810 1014.120 1711.130 1014.180 ;
        RECT 1711.820 1014.120 1711.960 1014.320 ;
        RECT 1746.690 1014.260 1747.010 1014.320 ;
        RECT 2283.050 1014.460 2283.370 1014.520 ;
        RECT 2601.370 1014.460 2601.690 1014.520 ;
        RECT 2283.050 1014.320 2601.690 1014.460 ;
        RECT 2283.050 1014.260 2283.370 1014.320 ;
        RECT 2601.370 1014.260 2601.690 1014.320 ;
        RECT 1710.810 1013.980 1711.960 1014.120 ;
        RECT 2049.370 1014.120 2049.690 1014.180 ;
        RECT 2052.590 1014.120 2052.910 1014.180 ;
        RECT 2049.370 1013.980 2052.910 1014.120 ;
        RECT 1710.810 1013.920 1711.130 1013.980 ;
        RECT 2049.370 1013.920 2049.690 1013.980 ;
        RECT 2052.590 1013.920 2052.910 1013.980 ;
        RECT 1938.510 1011.060 1938.830 1011.120 ;
        RECT 2501.090 1011.060 2501.410 1011.120 ;
        RECT 1938.510 1010.920 2501.410 1011.060 ;
        RECT 1938.510 1010.860 1938.830 1010.920 ;
        RECT 2501.090 1010.860 2501.410 1010.920 ;
        RECT 1910.910 1010.720 1911.230 1010.780 ;
        RECT 2498.790 1010.720 2499.110 1010.780 ;
        RECT 1910.910 1010.580 2499.110 1010.720 ;
        RECT 1910.910 1010.520 1911.230 1010.580 ;
        RECT 2498.790 1010.520 2499.110 1010.580 ;
        RECT 2052.590 1008.000 2052.910 1008.060 ;
        RECT 2501.550 1008.000 2501.870 1008.060 ;
        RECT 2052.590 1007.860 2501.870 1008.000 ;
        RECT 2052.590 1007.800 2052.910 1007.860 ;
        RECT 2501.550 1007.800 2501.870 1007.860 ;
        RECT 2238.890 1005.960 2239.210 1006.020 ;
        RECT 2498.330 1005.960 2498.650 1006.020 ;
        RECT 2238.890 1005.820 2498.650 1005.960 ;
        RECT 2238.890 1005.760 2239.210 1005.820 ;
        RECT 2498.330 1005.760 2498.650 1005.820 ;
        RECT 1897.110 1005.620 1897.430 1005.680 ;
        RECT 2499.250 1005.620 2499.570 1005.680 ;
        RECT 1897.110 1005.480 2499.570 1005.620 ;
        RECT 1897.110 1005.420 1897.430 1005.480 ;
        RECT 2499.250 1005.420 2499.570 1005.480 ;
        RECT 1890.210 1005.280 1890.530 1005.340 ;
        RECT 2499.710 1005.280 2500.030 1005.340 ;
        RECT 1890.210 1005.140 2500.030 1005.280 ;
        RECT 1890.210 1005.080 1890.530 1005.140 ;
        RECT 2499.710 1005.080 2500.030 1005.140 ;
        RECT 1876.410 1004.940 1876.730 1005.000 ;
        RECT 2500.170 1004.940 2500.490 1005.000 ;
        RECT 1876.410 1004.800 2500.490 1004.940 ;
        RECT 1876.410 1004.740 1876.730 1004.800 ;
        RECT 2500.170 1004.740 2500.490 1004.800 ;
        RECT 1862.610 1004.600 1862.930 1004.660 ;
        RECT 2500.630 1004.600 2500.950 1004.660 ;
        RECT 1862.610 1004.460 2500.950 1004.600 ;
        RECT 1862.610 1004.400 1862.930 1004.460 ;
        RECT 2500.630 1004.400 2500.950 1004.460 ;
      LAYER met1 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
      LAYER met1 ;
        RECT 1898.950 917.560 1899.270 917.620 ;
        RECT 2052.590 917.560 2052.910 917.620 ;
        RECT 1898.950 917.420 2052.910 917.560 ;
        RECT 1898.950 917.360 1899.270 917.420 ;
        RECT 2052.590 917.360 2052.910 917.420 ;
        RECT 1900.330 689.760 1900.650 689.820 ;
        RECT 1900.790 689.760 1901.110 689.820 ;
        RECT 1900.330 689.620 1901.110 689.760 ;
        RECT 1900.330 689.560 1900.650 689.620 ;
        RECT 1900.790 689.560 1901.110 689.620 ;
        RECT 1898.950 676.160 1899.270 676.220 ;
        RECT 1900.330 676.160 1900.650 676.220 ;
        RECT 1898.950 676.020 1900.650 676.160 ;
        RECT 1898.950 675.960 1899.270 676.020 ;
        RECT 1900.330 675.960 1900.650 676.020 ;
        RECT 1904.010 620.740 1904.330 620.800 ;
        RECT 1959.670 620.740 1959.990 620.800 ;
        RECT 1904.010 620.600 1959.990 620.740 ;
        RECT 1904.010 620.540 1904.330 620.600 ;
        RECT 1959.670 620.540 1959.990 620.600 ;
        RECT 1904.010 592.180 1904.330 592.240 ;
        RECT 1942.190 592.180 1942.510 592.240 ;
        RECT 1904.010 592.040 1942.510 592.180 ;
        RECT 1904.010 591.980 1904.330 592.040 ;
        RECT 1942.190 591.980 1942.510 592.040 ;
        RECT 1903.550 579.600 1903.870 579.660 ;
        RECT 1969.790 579.600 1970.110 579.660 ;
        RECT 1903.550 579.460 1970.110 579.600 ;
        RECT 1903.550 579.400 1903.870 579.460 ;
        RECT 1969.790 579.400 1970.110 579.460 ;
        RECT 1904.010 579.260 1904.330 579.320 ;
        RECT 1955.990 579.260 1956.310 579.320 ;
        RECT 1904.010 579.120 1956.310 579.260 ;
        RECT 1904.010 579.060 1904.330 579.120 ;
        RECT 1955.990 579.060 1956.310 579.120 ;
      LAYER met1 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met1 ;
        RECT 1503.810 554.780 1504.130 554.840 ;
        RECT 2083.870 554.780 2084.190 554.840 ;
        RECT 1503.810 554.640 2084.190 554.780 ;
        RECT 1503.810 554.580 1504.130 554.640 ;
        RECT 2083.870 554.580 2084.190 554.640 ;
      LAYER via ;
        RECT 2442.700 3066.840 2442.960 3067.100 ;
        RECT 2469.840 3066.840 2470.100 3067.100 ;
        RECT 1868.160 3063.780 1868.420 3064.040 ;
        RECT 1898.060 3063.780 1898.320 3064.040 ;
        RECT 2442.700 3063.780 2442.960 3064.040 ;
        RECT 2469.840 3063.780 2470.100 3064.040 ;
        RECT 2497.900 3063.780 2498.160 3064.040 ;
        RECT 1899.900 3051.880 1900.160 3052.140 ;
        RECT 2482.260 3051.880 2482.520 3052.140 ;
        RECT 1938.540 3029.100 1938.800 3029.360 ;
        RECT 2083.900 3029.100 2084.160 3029.360 ;
        RECT 1924.740 3022.300 1925.000 3022.560 ;
        RECT 2083.900 3022.300 2084.160 3022.560 ;
        RECT 1910.940 3015.500 1911.200 3015.760 ;
        RECT 2083.900 3015.500 2084.160 3015.760 ;
        RECT 1897.140 3008.360 1897.400 3008.620 ;
        RECT 2083.900 3008.360 2084.160 3008.620 ;
        RECT 1890.240 3001.560 1890.500 3001.820 ;
        RECT 2083.900 3001.560 2084.160 3001.820 ;
        RECT 2069.640 2697.940 2069.900 2698.200 ;
        RECT 2084.820 2697.940 2085.080 2698.200 ;
        RECT 1897.600 2691.140 1897.860 2691.400 ;
        RECT 1898.980 2691.140 1899.240 2691.400 ;
        RECT 2052.620 2691.140 2052.880 2691.400 ;
        RECT 2083.900 2691.140 2084.160 2691.400 ;
        RECT 1897.600 2680.260 1897.860 2680.520 ;
        RECT 1898.980 2680.260 1899.240 2680.520 ;
        RECT 2049.400 2607.840 2049.660 2608.100 ;
        RECT 2052.620 2607.840 2052.880 2608.100 ;
        RECT 1486.360 2604.440 1486.620 2604.700 ;
        RECT 2049.400 2604.440 2049.660 2604.700 ;
        RECT 1898.060 2594.580 1898.320 2594.840 ;
        RECT 1898.980 2594.580 1899.240 2594.840 ;
        RECT 1600.440 2594.240 1600.700 2594.500 ;
        RECT 1644.600 2594.240 1644.860 2594.500 ;
        RECT 1648.280 2594.240 1648.540 2594.500 ;
        RECT 1744.880 2594.240 1745.140 2594.500 ;
        RECT 2277.100 2594.240 2277.360 2594.500 ;
        RECT 1448.640 2593.900 1448.900 2594.160 ;
        RECT 1614.700 2593.900 1614.960 2594.160 ;
        RECT 1636.780 2593.900 1637.040 2594.160 ;
        RECT 1684.620 2593.900 1684.880 2594.160 ;
        RECT 1726.480 2593.900 1726.740 2594.160 ;
        RECT 2242.600 2593.900 2242.860 2594.160 ;
        RECT 2243.520 2593.900 2243.780 2594.160 ;
        RECT 2291.820 2593.900 2292.080 2594.160 ;
        RECT 1538.340 2593.560 1538.600 2593.820 ;
        RECT 1656.560 2593.560 1656.820 2593.820 ;
        RECT 1657.020 2593.560 1657.280 2593.820 ;
        RECT 1703.020 2593.560 1703.280 2593.820 ;
        RECT 1732.920 2593.560 1733.180 2593.820 ;
        RECT 2249.500 2593.560 2249.760 2593.820 ;
        RECT 2256.400 2593.560 2256.660 2593.820 ;
        RECT 2297.800 2593.560 2298.060 2593.820 ;
        RECT 1572.840 2593.220 1573.100 2593.480 ;
        RECT 1615.620 2593.220 1615.880 2593.480 ;
        RECT 1662.080 2593.220 1662.340 2593.480 ;
        RECT 1707.620 2593.220 1707.880 2593.480 ;
        RECT 2215.920 2593.220 2216.180 2593.480 ;
        RECT 2262.840 2593.220 2263.100 2593.480 ;
        RECT 1593.540 2592.880 1593.800 2593.140 ;
        RECT 1636.780 2592.880 1637.040 2593.140 ;
        RECT 1648.280 2592.880 1648.540 2593.140 ;
        RECT 1690.600 2592.880 1690.860 2593.140 ;
        RECT 1738.440 2592.880 1738.700 2593.140 ;
        RECT 2263.300 2592.880 2263.560 2593.140 ;
        RECT 1605.500 2592.540 1605.760 2592.800 ;
        RECT 1650.580 2592.540 1650.840 2592.800 ;
        RECT 1697.500 2592.540 1697.760 2592.800 ;
        RECT 1744.880 2592.540 1745.140 2592.800 ;
        RECT 2212.700 2592.540 2212.960 2592.800 ;
        RECT 2256.400 2592.540 2256.660 2592.800 ;
        RECT 2285.380 2593.220 2285.640 2593.480 ;
        RECT 2332.300 2593.220 2332.560 2593.480 ;
        RECT 2305.160 2592.540 2305.420 2592.800 ;
        RECT 1372.740 2592.200 1373.000 2592.460 ;
        RECT 1580.200 2592.200 1580.460 2592.460 ;
        RECT 1586.640 2592.200 1586.900 2592.460 ;
        RECT 1632.180 2592.200 1632.440 2592.460 ;
        RECT 1679.100 2592.200 1679.360 2592.460 ;
        RECT 1726.480 2592.200 1726.740 2592.460 ;
        RECT 2239.840 2592.200 2240.100 2592.460 ;
        RECT 2285.380 2592.200 2285.640 2592.460 ;
        RECT 2291.820 2592.200 2292.080 2592.460 ;
        RECT 2332.300 2592.200 2332.560 2592.460 ;
        RECT 1565.940 2591.860 1566.200 2592.120 ;
        RECT 1358.940 2591.520 1359.200 2591.780 ;
        RECT 1573.300 2591.520 1573.560 2591.780 ;
        RECT 1586.180 2591.860 1586.440 2592.120 ;
        RECT 1627.120 2591.860 1627.380 2592.120 ;
        RECT 1627.580 2591.860 1627.840 2592.120 ;
        RECT 1657.020 2591.860 1657.280 2592.120 ;
        RECT 1668.980 2591.860 1669.240 2592.120 ;
        RECT 1714.980 2591.860 1715.240 2592.120 ;
        RECT 1848.840 2591.860 1849.100 2592.120 ;
        RECT 2132.200 2591.860 2132.460 2592.120 ;
        RECT 2221.440 2591.860 2221.700 2592.120 ;
        RECT 2268.820 2591.860 2269.080 2592.120 ;
        RECT 2311.600 2591.860 2311.860 2592.120 ;
        RECT 1594.000 2591.520 1594.260 2591.780 ;
        RECT 1684.620 2591.520 1684.880 2591.780 ;
        RECT 1732.920 2591.520 1733.180 2591.780 ;
        RECT 1786.740 2591.520 1787.000 2591.780 ;
        RECT 2152.900 2591.520 2153.160 2591.780 ;
        RECT 2179.580 2591.520 2179.840 2591.780 ;
        RECT 2226.960 2591.520 2227.220 2591.780 ;
        RECT 2276.640 2591.520 2276.900 2591.780 ;
        RECT 2318.500 2591.520 2318.760 2591.780 ;
        RECT 1345.140 2591.180 1345.400 2591.440 ;
        RECT 1566.400 2591.180 1566.660 2591.440 ;
        RECT 1579.280 2591.180 1579.540 2591.440 ;
        RECT 1600.900 2591.180 1601.160 2591.440 ;
        RECT 1627.120 2591.180 1627.380 2591.440 ;
        RECT 1673.580 2591.180 1673.840 2591.440 ;
        RECT 1718.660 2591.180 1718.920 2591.440 ;
        RECT 1721.880 2591.180 1722.140 2591.440 ;
        RECT 1772.940 2591.180 1773.200 2591.440 ;
        RECT 2146.460 2591.180 2146.720 2591.440 ;
        RECT 2184.640 2590.840 2184.900 2591.100 ;
        RECT 2232.020 2591.180 2232.280 2591.440 ;
        RECT 2280.320 2591.180 2280.580 2591.440 ;
        RECT 2325.400 2591.180 2325.660 2591.440 ;
        RECT 1434.840 2590.500 1435.100 2590.760 ;
        RECT 1608.720 2590.500 1608.980 2590.760 ;
        RECT 1655.640 2590.500 1655.900 2590.760 ;
        RECT 1704.400 2590.500 1704.660 2590.760 ;
        RECT 1759.140 2590.500 1759.400 2590.760 ;
        RECT 2146.000 2590.500 2146.260 2590.760 ;
        RECT 2204.420 2590.500 2204.680 2590.760 ;
        RECT 2250.880 2590.840 2251.140 2591.100 ;
        RECT 2297.800 2590.840 2298.060 2591.100 ;
        RECT 2339.200 2590.840 2339.460 2591.100 ;
        RECT 1427.940 2590.160 1428.200 2590.420 ;
        RECT 1579.280 2590.160 1579.540 2590.420 ;
        RECT 1579.740 2590.160 1580.000 2590.420 ;
        RECT 1621.600 2590.160 1621.860 2590.420 ;
        RECT 1627.580 2590.160 1627.840 2590.420 ;
        RECT 1628.040 2590.160 1628.300 2590.420 ;
        RECT 1697.500 2590.160 1697.760 2590.420 ;
        RECT 1745.340 2590.160 1745.600 2590.420 ;
        RECT 2126.680 2590.160 2126.940 2590.420 ;
        RECT 2163.020 2590.160 2163.280 2590.420 ;
        RECT 2212.700 2590.160 2212.960 2590.420 ;
        RECT 1414.140 2589.820 1414.400 2590.080 ;
        RECT 1594.000 2589.820 1594.260 2590.080 ;
        RECT 1641.840 2589.820 1642.100 2590.080 ;
        RECT 1697.960 2589.820 1698.220 2590.080 ;
        RECT 1703.020 2589.820 1703.280 2590.080 ;
        RECT 2187.400 2589.820 2187.660 2590.080 ;
        RECT 2197.520 2589.820 2197.780 2590.080 ;
        RECT 2243.520 2589.820 2243.780 2590.080 ;
        RECT 1400.340 2589.480 1400.600 2589.740 ;
        RECT 1587.560 2589.480 1587.820 2589.740 ;
        RECT 1614.240 2589.480 1614.500 2589.740 ;
        RECT 1690.600 2589.480 1690.860 2589.740 ;
        RECT 1707.620 2589.480 1707.880 2589.740 ;
        RECT 2201.200 2589.480 2201.460 2589.740 ;
        RECT 2220.520 2589.480 2220.780 2589.740 ;
        RECT 2349.320 2589.480 2349.580 2589.740 ;
        RECT 1386.540 2589.140 1386.800 2589.400 ;
        RECT 1587.100 2589.140 1587.360 2589.400 ;
        RECT 1607.340 2589.140 1607.600 2589.400 ;
        RECT 1683.700 2589.140 1683.960 2589.400 ;
        RECT 1714.980 2589.140 1715.240 2589.400 ;
        RECT 2215.000 2589.140 2215.260 2589.400 ;
        RECT 2227.880 2589.140 2228.140 2589.400 ;
        RECT 2383.820 2589.140 2384.080 2589.400 ;
        RECT 1579.740 2588.800 1580.000 2589.060 ;
        RECT 1669.900 2588.800 1670.160 2589.060 ;
        RECT 1721.880 2588.800 1722.140 2589.060 ;
        RECT 2228.800 2588.800 2229.060 2589.060 ;
        RECT 1565.940 2588.460 1566.200 2588.720 ;
        RECT 1663.460 2588.460 1663.720 2588.720 ;
        RECT 1669.440 2588.460 1669.700 2588.720 ;
        RECT 1711.300 2588.460 1711.560 2588.720 ;
        RECT 1721.420 2588.460 1721.680 2588.720 ;
        RECT 1739.360 2588.460 1739.620 2588.720 ;
        RECT 2235.240 2588.460 2235.500 2588.720 ;
        RECT 2370.020 2588.460 2370.280 2588.720 ;
        RECT 1524.540 2588.120 1524.800 2588.380 ;
        RECT 1649.200 2588.120 1649.460 2588.380 ;
        RECT 1686.920 2588.120 1687.180 2588.380 ;
        RECT 1718.200 2588.120 1718.460 2588.380 ;
        RECT 2190.620 2588.120 2190.880 2588.380 ;
        RECT 2235.700 2588.120 2235.960 2588.380 ;
        RECT 2241.680 2588.120 2241.940 2588.380 ;
        RECT 2356.220 2588.120 2356.480 2588.380 ;
        RECT 1552.140 2587.780 1552.400 2588.040 ;
        RECT 1663.000 2587.780 1663.260 2588.040 ;
        RECT 1703.940 2587.780 1704.200 2588.040 ;
        RECT 1732.000 2587.780 1732.260 2588.040 ;
        RECT 2183.720 2587.780 2183.980 2588.040 ;
        RECT 2186.480 2587.780 2186.740 2588.040 ;
        RECT 2232.020 2587.780 2232.280 2588.040 ;
        RECT 1331.340 2587.440 1331.600 2587.700 ;
        RECT 1560.880 2587.440 1561.140 2587.700 ;
        RECT 1627.580 2587.440 1627.840 2587.700 ;
        RECT 1668.980 2587.440 1669.240 2587.700 ;
        RECT 1697.040 2587.440 1697.300 2587.700 ;
        RECT 1726.020 2587.440 1726.280 2587.700 ;
        RECT 1731.540 2587.440 1731.800 2587.700 ;
        RECT 1738.900 2587.440 1739.160 2587.700 ;
        RECT 2170.840 2587.440 2171.100 2587.700 ;
        RECT 2215.920 2587.440 2216.180 2587.700 ;
        RECT 2227.420 2587.440 2227.680 2587.700 ;
        RECT 2397.620 2587.440 2397.880 2587.700 ;
        RECT 1898.060 2570.100 1898.320 2570.360 ;
        RECT 1898.980 2570.100 1899.240 2570.360 ;
        RECT 2170.380 2559.900 2170.640 2560.160 ;
        RECT 2170.840 2559.900 2171.100 2560.160 ;
        RECT 1898.060 2497.680 1898.320 2497.940 ;
        RECT 1898.980 2497.680 1899.240 2497.940 ;
        RECT 1898.060 2473.540 1898.320 2473.800 ;
        RECT 1898.980 2473.540 1899.240 2473.800 ;
        RECT 2168.080 2463.000 2168.340 2463.260 ;
        RECT 2169.460 2463.000 2169.720 2463.260 ;
        RECT 1408.620 2414.720 1408.880 2414.980 ;
        RECT 1414.140 2414.720 1414.400 2414.980 ;
        RECT 1559.040 2414.720 1559.300 2414.980 ;
        RECT 1832.280 2414.720 1832.540 2414.980 ;
        RECT 1858.040 2414.720 1858.300 2414.980 ;
        RECT 2087.580 2414.720 2087.840 2414.980 ;
        RECT 2165.780 2414.720 2166.040 2414.980 ;
        RECT 2197.520 2414.720 2197.780 2414.980 ;
        RECT 2276.640 2414.720 2276.900 2414.980 ;
        RECT 2538.840 2414.720 2539.100 2414.980 ;
        RECT 1537.880 2414.380 1538.140 2414.640 ;
        RECT 1487.280 2414.040 1487.540 2414.300 ;
        RECT 1932.560 2414.040 1932.820 2414.300 ;
        RECT 1934.860 2414.380 1935.120 2414.640 ;
        RECT 1938.540 2414.380 1938.800 2414.640 ;
        RECT 2269.740 2414.380 2270.000 2414.640 ;
        RECT 2525.960 2414.380 2526.220 2414.640 ;
        RECT 1947.740 2414.040 1948.000 2414.300 ;
        RECT 2283.540 2414.040 2283.800 2414.300 ;
        RECT 2551.260 2414.040 2551.520 2414.300 ;
        RECT 1487.740 2413.700 1488.000 2413.960 ;
        RECT 1973.500 2413.700 1973.760 2413.960 ;
        RECT 2153.360 2413.700 2153.620 2413.960 ;
        RECT 2190.620 2413.700 2190.880 2413.960 ;
        RECT 2290.440 2413.700 2290.700 2413.960 ;
        RECT 2564.140 2413.700 2564.400 2413.960 ;
        RECT 1421.500 2413.360 1421.760 2413.620 ;
        RECT 1427.940 2413.360 1428.200 2413.620 ;
        RECT 1488.200 2413.360 1488.460 2413.620 ;
        RECT 1986.380 2413.360 1986.640 2413.620 ;
        RECT 2140.480 2413.360 2140.740 2413.620 ;
        RECT 2183.720 2413.360 2183.980 2413.620 ;
        RECT 2297.340 2413.360 2297.600 2413.620 ;
        RECT 2577.020 2413.360 2577.280 2413.620 ;
        RECT 1488.660 2413.020 1488.920 2413.280 ;
        RECT 1999.260 2413.020 1999.520 2413.280 ;
        RECT 2127.600 2413.020 2127.860 2413.280 ;
        RECT 2184.640 2413.020 2184.900 2413.280 ;
        RECT 2304.240 2413.020 2304.500 2413.280 ;
        RECT 2589.900 2413.020 2590.160 2413.280 ;
        RECT 1395.740 2412.680 1396.000 2412.940 ;
        RECT 1400.340 2412.680 1400.600 2412.940 ;
        RECT 1489.120 2412.680 1489.380 2412.940 ;
        RECT 2012.140 2412.680 2012.400 2412.940 ;
        RECT 2063.660 2412.680 2063.920 2412.940 ;
        RECT 2069.640 2412.680 2069.900 2412.940 ;
        RECT 2114.720 2412.680 2114.980 2412.940 ;
        RECT 2176.820 2412.680 2177.080 2412.940 ;
        RECT 2303.780 2412.680 2304.040 2412.940 ;
        RECT 2602.780 2412.680 2603.040 2412.940 ;
        RECT 1489.580 2412.340 1489.840 2412.600 ;
        RECT 2025.020 2412.340 2025.280 2412.600 ;
        RECT 2166.240 2412.340 2166.500 2412.600 ;
        RECT 2294.580 2412.340 2294.840 2412.600 ;
        RECT 2318.040 2412.340 2318.300 2412.600 ;
        RECT 2628.540 2412.340 2628.800 2412.600 ;
        RECT 1490.040 2412.000 1490.300 2412.260 ;
        RECT 2037.900 2412.000 2038.160 2412.260 ;
        RECT 2173.140 2412.000 2173.400 2412.260 ;
        RECT 2307.460 2412.000 2307.720 2412.260 ;
        RECT 2311.140 2412.000 2311.400 2412.260 ;
        RECT 2615.660 2412.000 2615.920 2412.260 ;
        RECT 1486.820 2411.660 1487.080 2411.920 ;
        RECT 2076.540 2411.660 2076.800 2411.920 ;
        RECT 2101.840 2411.660 2102.100 2411.920 ;
        RECT 2169.000 2411.660 2169.260 2411.920 ;
        RECT 2180.040 2411.660 2180.300 2411.920 ;
        RECT 2320.340 2411.660 2320.600 2411.920 ;
        RECT 2324.940 2411.660 2325.200 2411.920 ;
        RECT 2641.420 2411.660 2641.680 2411.920 ;
        RECT 1306.040 2411.320 1306.300 2411.580 ;
        RECT 1551.680 2410.980 1551.940 2411.240 ;
        RECT 1819.400 2410.980 1819.660 2411.240 ;
        RECT 1551.220 2410.640 1551.480 2410.900 ;
        RECT 1806.520 2410.640 1806.780 2410.900 ;
        RECT 1545.240 2410.300 1545.500 2410.560 ;
        RECT 1793.640 2410.300 1793.900 2410.560 ;
        RECT 1883.800 2411.320 1884.060 2411.580 ;
        RECT 1890.240 2411.320 1890.500 2411.580 ;
        RECT 1932.560 2411.320 1932.820 2411.580 ;
        RECT 1960.620 2411.320 1960.880 2411.580 ;
        RECT 2088.960 2411.320 2089.220 2411.580 ;
        RECT 2163.020 2411.320 2163.280 2411.580 ;
        RECT 2186.940 2411.320 2187.200 2411.580 ;
        RECT 2333.220 2411.320 2333.480 2411.580 ;
        RECT 2338.740 2411.320 2339.000 2411.580 ;
        RECT 2667.180 2411.320 2667.440 2411.580 ;
        RECT 1870.920 2410.980 1871.180 2411.240 ;
        RECT 2087.120 2410.980 2087.380 2411.240 ;
        RECT 2269.280 2410.980 2269.540 2411.240 ;
        RECT 2513.080 2410.980 2513.340 2411.240 ;
        RECT 2179.120 2410.640 2179.380 2410.900 ;
        RECT 2204.420 2410.640 2204.680 2410.900 ;
        RECT 2262.840 2410.640 2263.100 2410.900 ;
        RECT 2500.200 2410.640 2500.460 2410.900 ;
        RECT 1898.980 2410.300 1899.240 2410.560 ;
        RECT 2255.940 2410.300 2256.200 2410.560 ;
        RECT 2487.320 2410.300 2487.580 2410.560 ;
        RECT 1382.860 2409.960 1383.120 2410.220 ;
        RECT 1386.540 2409.960 1386.800 2410.220 ;
        RECT 1460.140 2409.960 1460.400 2410.220 ;
        RECT 1600.900 2409.960 1601.160 2410.220 ;
        RECT 1601.360 2409.960 1601.620 2410.220 ;
        RECT 1607.340 2409.960 1607.600 2410.220 ;
        RECT 1607.800 2409.960 1608.060 2410.220 ;
        RECT 1622.520 2409.960 1622.780 2410.220 ;
        RECT 1665.300 2409.960 1665.560 2410.220 ;
        RECT 1669.440 2409.960 1669.700 2410.220 ;
        RECT 1691.060 2409.960 1691.320 2410.220 ;
        RECT 1697.040 2409.960 1697.300 2410.220 ;
        RECT 1716.820 2409.960 1717.080 2410.220 ;
        RECT 1721.420 2409.960 1721.680 2410.220 ;
        RECT 1755.460 2409.960 1755.720 2410.220 ;
        RECT 1759.140 2409.960 1759.400 2410.220 ;
        RECT 1768.340 2409.960 1768.600 2410.220 ;
        RECT 1772.940 2409.960 1773.200 2410.220 ;
        RECT 2249.040 2409.960 2249.300 2410.220 ;
        RECT 2474.440 2409.960 2474.700 2410.220 ;
        RECT 1472.560 2409.620 1472.820 2409.880 ;
        RECT 1622.060 2409.620 1622.320 2409.880 ;
        RECT 1628.960 2409.620 1629.220 2409.880 ;
        RECT 1485.440 2409.280 1485.700 2409.540 ;
        RECT 1628.500 2409.280 1628.760 2409.540 ;
        RECT 1498.320 2408.940 1498.580 2409.200 ;
        RECT 1635.860 2408.940 1636.120 2409.200 ;
        RECT 1511.200 2408.600 1511.460 2408.860 ;
        RECT 1642.300 2408.600 1642.560 2408.860 ;
        RECT 2214.540 2409.620 2214.800 2409.880 ;
        RECT 2397.160 2409.620 2397.420 2409.880 ;
        RECT 2397.620 2409.620 2397.880 2409.880 ;
        RECT 2422.920 2409.620 2423.180 2409.880 ;
        RECT 1780.760 2409.280 1781.020 2409.540 ;
        RECT 1786.740 2409.280 1787.000 2409.540 ;
        RECT 2207.640 2409.280 2207.900 2409.540 ;
        RECT 2384.740 2409.280 2385.000 2409.540 ;
        RECT 2200.740 2408.940 2201.000 2409.200 ;
        RECT 2371.860 2408.940 2372.120 2409.200 ;
        RECT 2383.820 2408.940 2384.080 2409.200 ;
        RECT 2435.800 2409.280 2436.060 2409.540 ;
        RECT 1676.800 2408.600 1677.060 2408.860 ;
        RECT 1678.180 2408.600 1678.440 2408.860 ;
        RECT 1686.920 2408.600 1687.180 2408.860 ;
        RECT 2193.840 2408.600 2194.100 2408.860 ;
        RECT 2358.980 2408.600 2359.240 2408.860 ;
        RECT 2370.020 2408.600 2370.280 2408.860 ;
        RECT 2448.680 2408.940 2448.940 2409.200 ;
        RECT 2386.120 2408.600 2386.380 2408.860 ;
        RECT 2461.560 2408.600 2461.820 2408.860 ;
        RECT 1575.600 2408.260 1575.860 2408.520 ;
        RECT 1579.740 2408.260 1580.000 2408.520 ;
        RECT 1588.480 2408.260 1588.740 2408.520 ;
        RECT 1628.500 2408.260 1628.760 2408.520 ;
        RECT 2193.380 2408.260 2193.640 2408.520 ;
        RECT 2346.100 2408.260 2346.360 2408.520 ;
        RECT 2349.320 2408.260 2349.580 2408.520 ;
        RECT 2385.660 2408.260 2385.920 2408.520 ;
        RECT 2386.580 2408.260 2386.840 2408.520 ;
        RECT 2410.040 2408.260 2410.300 2408.520 ;
        RECT 1655.640 1193.440 1655.900 1193.700 ;
        RECT 1703.940 1193.440 1704.200 1193.700 ;
        RECT 2166.240 1193.440 2166.500 1193.700 ;
        RECT 2245.820 1193.440 2246.080 1193.700 ;
        RECT 2320.340 1193.440 2320.600 1193.700 ;
        RECT 2385.200 1193.440 2385.460 1193.700 ;
        RECT 2386.120 1193.440 2386.380 1193.700 ;
        RECT 2487.320 1193.440 2487.580 1193.700 ;
        RECT 1626.660 1193.100 1626.920 1193.360 ;
        RECT 1683.700 1193.100 1683.960 1193.360 ;
        RECT 1956.020 1193.100 1956.280 1193.360 ;
        RECT 2025.020 1193.100 2025.280 1193.360 ;
        RECT 2153.360 1193.100 2153.620 1193.360 ;
        RECT 2252.720 1193.100 2252.980 1193.360 ;
        RECT 2294.580 1193.100 2294.840 1193.360 ;
        RECT 2397.620 1193.100 2397.880 1193.360 ;
        RECT 1318.460 1192.760 1318.720 1193.020 ;
        RECT 1489.120 1192.760 1489.380 1193.020 ;
        RECT 1648.740 1192.760 1649.000 1193.020 ;
        RECT 1716.820 1192.760 1717.080 1193.020 ;
        RECT 1942.220 1192.760 1942.480 1193.020 ;
        RECT 2012.140 1192.760 2012.400 1193.020 ;
        RECT 2140.480 1192.760 2140.740 1193.020 ;
        RECT 2259.620 1192.760 2259.880 1193.020 ;
        RECT 2318.040 1192.760 2318.300 1193.020 ;
        RECT 2525.960 1192.760 2526.220 1193.020 ;
        RECT 1641.840 1192.420 1642.100 1192.680 ;
        RECT 1729.700 1192.420 1729.960 1192.680 ;
        RECT 1901.740 1192.420 1902.000 1192.680 ;
        RECT 1973.500 1192.420 1973.760 1192.680 ;
        RECT 2101.840 1192.420 2102.100 1192.680 ;
        RECT 2281.240 1192.420 2281.500 1192.680 ;
        RECT 2304.240 1192.420 2304.500 1192.680 ;
        RECT 2564.140 1192.420 2564.400 1192.680 ;
        RECT 1485.440 1192.080 1485.700 1192.340 ;
        RECT 1735.220 1192.080 1735.480 1192.340 ;
        RECT 1901.280 1192.080 1901.540 1192.340 ;
        RECT 1986.380 1192.080 1986.640 1192.340 ;
        RECT 2088.960 1192.080 2089.220 1192.340 ;
        RECT 2280.320 1192.080 2280.580 1192.340 ;
        RECT 2290.440 1192.080 2290.700 1192.340 ;
        RECT 2589.900 1192.080 2590.160 1192.340 ;
        RECT 1472.560 1191.740 1472.820 1192.000 ;
        RECT 1721.420 1191.740 1721.680 1192.000 ;
        RECT 1855.740 1191.740 1856.000 1192.000 ;
        RECT 1947.740 1191.740 1948.000 1192.000 ;
        RECT 1969.820 1191.740 1970.080 1192.000 ;
        RECT 2037.900 1191.740 2038.160 1192.000 ;
        RECT 2114.720 1191.740 2114.980 1192.000 ;
        RECT 2273.420 1191.740 2273.680 1192.000 ;
        RECT 2276.180 1191.740 2276.440 1192.000 ;
        RECT 2615.660 1191.740 2615.920 1192.000 ;
        RECT 1447.260 1191.400 1447.520 1191.660 ;
        RECT 1707.620 1191.400 1707.880 1191.660 ;
        RECT 1902.200 1191.400 1902.460 1191.660 ;
        RECT 2076.540 1191.400 2076.800 1191.660 ;
        RECT 2127.600 1191.400 2127.860 1191.660 ;
        RECT 2266.520 1191.400 2266.780 1191.660 ;
        RECT 2269.740 1191.400 2270.000 1191.660 ;
        RECT 2641.420 1191.400 2641.680 1191.660 ;
        RECT 1421.500 1191.060 1421.760 1191.320 ;
        RECT 1693.820 1191.060 1694.080 1191.320 ;
        RECT 1922.440 1191.060 1922.700 1191.320 ;
        RECT 2238.920 1191.060 2239.180 1191.320 ;
        RECT 2255.940 1191.060 2256.200 1191.320 ;
        RECT 2667.180 1191.060 2667.440 1191.320 ;
        RECT 1434.380 1190.720 1434.640 1190.980 ;
        RECT 1700.720 1190.720 1700.980 1190.980 ;
        RECT 1900.820 1190.720 1901.080 1190.980 ;
        RECT 1999.260 1190.720 1999.520 1190.980 ;
        RECT 2063.660 1190.720 2063.920 1190.980 ;
        RECT 2481.800 1190.720 2482.060 1190.980 ;
        RECT 1460.140 1190.380 1460.400 1190.640 ;
        RECT 1728.780 1190.380 1729.040 1190.640 ;
        RECT 1780.760 1190.380 1781.020 1190.640 ;
        RECT 2391.180 1190.380 2391.440 1190.640 ;
        RECT 1331.340 1190.040 1331.600 1190.300 ;
        RECT 1728.320 1190.040 1728.580 1190.300 ;
        RECT 1768.340 1190.040 1768.600 1190.300 ;
        RECT 2385.660 1190.040 2385.920 1190.300 ;
        RECT 2391.640 1190.040 2391.900 1190.300 ;
        RECT 2500.200 1190.040 2500.460 1190.300 ;
        RECT 2179.120 1189.700 2179.380 1189.960 ;
        RECT 2239.380 1189.700 2239.640 1189.960 ;
        RECT 2359.440 1189.700 2359.700 1189.960 ;
        RECT 2435.800 1189.700 2436.060 1189.960 ;
        RECT 2366.340 1189.360 2366.600 1189.620 ;
        RECT 2422.920 1189.360 2423.180 1189.620 ;
        RECT 2333.220 1189.020 2333.480 1189.280 ;
        RECT 2383.820 1189.020 2384.080 1189.280 ;
        RECT 2346.100 1188.680 2346.360 1188.940 ;
        RECT 2390.720 1188.680 2390.980 1188.940 ;
        RECT 2358.980 1188.000 2359.240 1188.260 ;
        RECT 2387.960 1188.000 2388.220 1188.260 ;
        RECT 1662.540 1187.660 1662.800 1187.920 ;
        RECT 1691.060 1187.660 1691.320 1187.920 ;
        RECT 2380.140 1187.660 2380.400 1187.920 ;
        RECT 2397.160 1187.660 2397.420 1187.920 ;
        RECT 1669.440 1187.320 1669.700 1187.580 ;
        RECT 1678.180 1187.320 1678.440 1187.580 ;
        RECT 2384.740 1187.320 2385.000 1187.580 ;
        RECT 2410.040 1187.320 2410.300 1187.580 ;
        RECT 1382.860 1186.980 1383.120 1187.240 ;
        RECT 1386.540 1186.980 1386.800 1187.240 ;
        RECT 1395.740 1186.980 1396.000 1187.240 ;
        RECT 1400.340 1186.980 1400.600 1187.240 ;
        RECT 1408.620 1186.980 1408.880 1187.240 ;
        RECT 1414.140 1186.980 1414.400 1187.240 ;
        RECT 1498.320 1186.980 1498.580 1187.240 ;
        RECT 1503.840 1186.980 1504.100 1187.240 ;
        RECT 1511.200 1186.980 1511.460 1187.240 ;
        RECT 1517.640 1186.980 1517.900 1187.240 ;
        RECT 1575.600 1186.980 1575.860 1187.240 ;
        RECT 1579.740 1186.980 1580.000 1187.240 ;
        RECT 1588.480 1186.980 1588.740 1187.240 ;
        RECT 1593.540 1186.980 1593.800 1187.240 ;
        RECT 1601.360 1186.980 1601.620 1187.240 ;
        RECT 1607.340 1186.980 1607.600 1187.240 ;
        RECT 1665.300 1186.980 1665.560 1187.240 ;
        RECT 1669.900 1186.980 1670.160 1187.240 ;
        RECT 1755.460 1186.980 1755.720 1187.240 ;
        RECT 1759.140 1186.980 1759.400 1187.240 ;
        RECT 1806.520 1186.980 1806.780 1187.240 ;
        RECT 1811.120 1186.980 1811.380 1187.240 ;
        RECT 1858.040 1186.980 1858.300 1187.240 ;
        RECT 1862.640 1186.980 1862.900 1187.240 ;
        RECT 1870.920 1186.980 1871.180 1187.240 ;
        RECT 1876.440 1186.980 1876.700 1187.240 ;
        RECT 1883.800 1186.980 1884.060 1187.240 ;
        RECT 1890.240 1186.980 1890.500 1187.240 ;
        RECT 1934.860 1186.980 1935.120 1187.240 ;
        RECT 1938.540 1186.980 1938.800 1187.240 ;
        RECT 2307.460 1186.980 2307.720 1187.240 ;
        RECT 2311.140 1186.980 2311.400 1187.240 ;
        RECT 2371.860 1186.980 2372.120 1187.240 ;
        RECT 2387.500 1186.980 2387.760 1187.240 ;
        RECT 2352.540 1025.820 2352.800 1026.080 ;
        RECT 2442.700 1025.820 2442.960 1026.080 ;
        RECT 2352.080 1025.140 2352.340 1025.400 ;
        RECT 2456.500 1025.140 2456.760 1025.400 ;
        RECT 2345.640 1024.800 2345.900 1025.060 ;
        RECT 2470.300 1024.800 2470.560 1025.060 ;
        RECT 1848.840 1024.460 1849.100 1024.720 ;
        RECT 2450.980 1024.460 2451.240 1024.720 ;
        RECT 2369.100 1022.080 2369.360 1022.340 ;
        RECT 2386.120 1022.080 2386.380 1022.340 ;
        RECT 1655.180 1021.060 1655.440 1021.320 ;
        RECT 1670.360 1021.060 1670.620 1021.320 ;
        RECT 1681.860 1021.060 1682.120 1021.320 ;
        RECT 1710.840 1021.060 1711.100 1021.320 ;
        RECT 1414.140 1020.720 1414.400 1020.980 ;
        RECT 1726.940 1021.400 1727.200 1021.660 ;
        RECT 1726.480 1021.060 1726.740 1021.320 ;
        RECT 1745.800 1021.060 1746.060 1021.320 ;
        RECT 1821.240 1021.060 1821.500 1021.320 ;
        RECT 1828.600 1021.060 1828.860 1021.320 ;
        RECT 2280.320 1021.060 2280.580 1021.320 ;
        RECT 2283.080 1021.060 2283.340 1021.320 ;
        RECT 2325.400 1021.060 2325.660 1021.320 ;
        RECT 2385.200 1021.060 2385.460 1021.320 ;
        RECT 2408.200 1021.060 2408.460 1021.320 ;
        RECT 1726.940 1020.720 1727.200 1020.980 ;
        RECT 1787.200 1020.720 1787.460 1020.980 ;
        RECT 1811.120 1020.720 1811.380 1020.980 ;
        RECT 1835.500 1020.720 1835.760 1020.980 ;
        RECT 2338.740 1020.720 2339.000 1020.980 ;
        RECT 2369.100 1020.720 2369.360 1020.980 ;
        RECT 2391.180 1020.720 2391.440 1020.980 ;
        RECT 2428.900 1020.720 2429.160 1020.980 ;
        RECT 1503.840 1020.380 1504.100 1020.640 ;
        RECT 1726.480 1020.380 1726.740 1020.640 ;
        RECT 1728.780 1020.380 1729.040 1020.640 ;
        RECT 1759.600 1020.380 1759.860 1020.640 ;
        RECT 2249.040 1020.380 2249.300 1020.640 ;
        RECT 2677.300 1020.380 2677.560 1020.640 ;
        RECT 1517.640 1020.040 1517.900 1020.300 ;
        RECT 1719.120 1020.040 1719.380 1020.300 ;
        RECT 1524.540 1019.700 1524.800 1019.960 ;
        RECT 1732.000 1020.040 1732.260 1020.300 ;
        RECT 1746.260 1020.040 1746.520 1020.300 ;
        RECT 1787.660 1020.040 1787.920 1020.300 ;
        RECT 1800.080 1020.040 1800.340 1020.300 ;
        RECT 2242.600 1020.040 2242.860 1020.300 ;
        RECT 2245.820 1020.040 2246.080 1020.300 ;
        RECT 2295.040 1020.040 2295.300 1020.300 ;
        RECT 2325.860 1020.040 2326.120 1020.300 ;
        RECT 2332.760 1020.040 2333.020 1020.300 ;
        RECT 2370.940 1020.040 2371.200 1020.300 ;
        RECT 2383.360 1020.040 2383.620 1020.300 ;
        RECT 2383.820 1020.040 2384.080 1020.300 ;
        RECT 2402.220 1020.040 2402.480 1020.300 ;
        RECT 1721.420 1019.700 1721.680 1019.960 ;
        RECT 1755.460 1019.700 1755.720 1019.960 ;
        RECT 1758.680 1019.700 1758.940 1019.960 ;
        RECT 1806.520 1019.700 1806.780 1019.960 ;
        RECT 2228.800 1019.700 2229.060 1019.960 ;
        RECT 2297.340 1019.700 2297.600 1019.960 ;
        RECT 2573.800 1019.700 2574.060 1019.960 ;
        RECT 1538.340 1019.360 1538.600 1019.620 ;
        RECT 1725.100 1019.360 1725.360 1019.620 ;
        RECT 1728.320 1019.360 1728.580 1019.620 ;
        RECT 1821.700 1019.360 1821.960 1019.620 ;
        RECT 2252.720 1019.360 2252.980 1019.620 ;
        RECT 2302.860 1019.360 2303.120 1019.620 ;
        RECT 2310.680 1019.360 2310.940 1019.620 ;
        RECT 2546.200 1019.360 2546.460 1019.620 ;
        RECT 1552.140 1019.020 1552.400 1019.280 ;
        RECT 1718.200 1019.020 1718.460 1019.280 ;
        RECT 1719.120 1019.020 1719.380 1019.280 ;
        RECT 1738.900 1019.020 1739.160 1019.280 ;
        RECT 1565.940 1018.680 1566.200 1018.940 ;
        RECT 1661.620 1018.680 1661.880 1018.940 ;
        RECT 1662.080 1018.680 1662.340 1018.940 ;
        RECT 1681.860 1018.680 1682.120 1018.940 ;
        RECT 1682.320 1018.680 1682.580 1018.940 ;
        RECT 1700.260 1018.680 1700.520 1018.940 ;
        RECT 1700.720 1018.680 1700.980 1018.940 ;
        RECT 1773.400 1018.680 1773.660 1018.940 ;
        RECT 1703.940 1018.340 1704.200 1018.600 ;
        RECT 1711.300 1018.340 1711.560 1018.600 ;
        RECT 1724.640 1018.340 1724.900 1018.600 ;
        RECT 1771.560 1018.340 1771.820 1018.600 ;
        RECT 1817.560 1019.020 1817.820 1019.280 ;
        RECT 2201.200 1019.020 2201.460 1019.280 ;
        RECT 2259.620 1019.020 2259.880 1019.280 ;
        RECT 2307.000 1019.020 2307.260 1019.280 ;
        RECT 2317.580 1019.020 2317.840 1019.280 ;
        RECT 2532.400 1019.020 2532.660 1019.280 ;
        RECT 1778.000 1018.680 1778.260 1018.940 ;
        RECT 1823.540 1018.680 1823.800 1018.940 ;
        RECT 2187.400 1018.680 2187.660 1018.940 ;
        RECT 2239.380 1018.680 2239.640 1018.940 ;
        RECT 2242.140 1018.680 2242.400 1018.940 ;
        RECT 2289.980 1018.680 2290.240 1018.940 ;
        RECT 2324.940 1018.680 2325.200 1018.940 ;
        RECT 2511.700 1018.680 2511.960 1018.940 ;
        RECT 2311.140 1018.340 2311.400 1018.600 ;
        RECT 2415.100 1018.340 2415.360 1018.600 ;
        RECT 1593.540 1018.000 1593.800 1018.260 ;
        RECT 1704.400 1018.000 1704.660 1018.260 ;
        RECT 1607.340 1017.660 1607.600 1017.920 ;
        RECT 1697.040 1017.660 1697.300 1017.920 ;
        RECT 1614.240 1017.320 1614.500 1017.580 ;
        RECT 1690.600 1017.320 1690.860 1017.580 ;
        RECT 1691.060 1017.320 1691.320 1017.580 ;
        RECT 1696.120 1017.320 1696.380 1017.580 ;
        RECT 1733.840 1017.660 1734.100 1017.920 ;
        RECT 1697.960 1017.320 1698.220 1017.580 ;
        RECT 1746.260 1018.000 1746.520 1018.260 ;
        RECT 1746.720 1018.000 1746.980 1018.260 ;
        RECT 1755.000 1018.000 1755.260 1018.260 ;
        RECT 1766.040 1018.000 1766.300 1018.260 ;
        RECT 1812.500 1018.000 1812.760 1018.260 ;
        RECT 2215.000 1018.000 2215.260 1018.260 ;
        RECT 2332.300 1018.000 2332.560 1018.260 ;
        RECT 2391.640 1018.000 2391.900 1018.260 ;
        RECT 2397.620 1018.000 2397.880 1018.260 ;
        RECT 2422.000 1018.000 2422.260 1018.260 ;
        RECT 1734.760 1017.660 1735.020 1017.920 ;
        RECT 1741.660 1017.660 1741.920 1017.920 ;
        RECT 1789.040 1017.660 1789.300 1017.920 ;
        RECT 2263.300 1017.660 2263.560 1017.920 ;
        RECT 2307.000 1017.660 2307.260 1017.920 ;
        RECT 2353.460 1017.660 2353.720 1017.920 ;
        RECT 1641.840 1016.980 1642.100 1017.240 ;
        RECT 1689.680 1016.980 1689.940 1017.240 ;
        RECT 1735.680 1017.320 1735.940 1017.580 ;
        RECT 1735.220 1016.980 1735.480 1017.240 ;
        RECT 1745.800 1016.980 1746.060 1017.240 ;
        RECT 1782.140 1016.980 1782.400 1017.240 ;
        RECT 2277.100 1016.980 2277.360 1017.240 ;
        RECT 2280.780 1016.980 2281.040 1017.240 ;
        RECT 1641.380 1016.640 1641.640 1016.900 ;
        RECT 1676.800 1016.640 1677.060 1016.900 ;
        RECT 1683.240 1016.640 1683.500 1016.900 ;
        RECT 1729.700 1016.640 1729.960 1016.900 ;
        RECT 1778.000 1016.640 1778.260 1016.900 ;
        RECT 1793.640 1016.640 1793.900 1016.900 ;
        RECT 1842.400 1016.640 1842.660 1016.900 ;
        RECT 1655.640 1016.300 1655.900 1016.560 ;
        RECT 1648.740 1015.960 1649.000 1016.220 ;
        RECT 1669.440 1016.300 1669.700 1016.560 ;
        RECT 1712.220 1016.300 1712.480 1016.560 ;
        RECT 1758.680 1016.300 1758.940 1016.560 ;
        RECT 1787.660 1016.300 1787.920 1016.560 ;
        RECT 1793.180 1016.300 1793.440 1016.560 ;
        RECT 2249.500 1016.300 2249.760 1016.560 ;
        RECT 2302.860 1016.980 2303.120 1017.240 ;
        RECT 2347.020 1017.320 2347.280 1017.580 ;
        RECT 2387.960 1017.320 2388.220 1017.580 ;
        RECT 2325.860 1016.980 2326.120 1017.240 ;
        RECT 2342.420 1016.980 2342.680 1017.240 ;
        RECT 2289.980 1016.640 2290.240 1016.900 ;
        RECT 2336.440 1016.640 2336.700 1016.900 ;
        RECT 2380.600 1016.640 2380.860 1016.900 ;
        RECT 2385.660 1016.980 2385.920 1017.240 ;
        RECT 2428.900 1016.980 2429.160 1017.240 ;
        RECT 2387.500 1016.640 2387.760 1016.900 ;
        RECT 2388.420 1016.640 2388.680 1016.900 ;
        RECT 2323.100 1016.300 2323.360 1016.560 ;
        RECT 2332.300 1016.300 2332.560 1016.560 ;
        RECT 2332.760 1016.300 2333.020 1016.560 ;
        RECT 2377.840 1016.300 2378.100 1016.560 ;
        RECT 1675.880 1015.960 1676.140 1016.220 ;
        RECT 1676.340 1015.960 1676.600 1016.220 ;
        RECT 1718.200 1015.960 1718.460 1016.220 ;
        RECT 1766.040 1015.960 1766.300 1016.220 ;
        RECT 1691.060 1015.620 1691.320 1015.880 ;
        RECT 1693.820 1015.620 1694.080 1015.880 ;
        RECT 1780.300 1015.620 1780.560 1015.880 ;
        RECT 2275.260 1015.620 2275.520 1015.880 ;
        RECT 2318.040 1015.620 2318.300 1015.880 ;
        RECT 2364.500 1015.960 2364.760 1016.220 ;
        RECT 2415.100 1016.300 2415.360 1016.560 ;
        RECT 2422.000 1015.960 2422.260 1016.220 ;
        RECT 1661.620 1015.280 1661.880 1015.540 ;
        RECT 1682.320 1015.280 1682.580 1015.540 ;
        RECT 1683.240 1015.280 1683.500 1015.540 ;
        RECT 1724.640 1015.280 1724.900 1015.540 ;
        RECT 1755.000 1015.280 1755.260 1015.540 ;
        RECT 1800.080 1015.280 1800.340 1015.540 ;
        RECT 2266.520 1015.280 2266.780 1015.540 ;
        RECT 2312.060 1015.280 2312.320 1015.540 ;
        RECT 2358.980 1015.280 2359.240 1015.540 ;
        RECT 2359.440 1015.280 2359.700 1015.540 ;
        RECT 2394.400 1015.280 2394.660 1015.540 ;
        RECT 2408.200 1015.620 2408.460 1015.880 ;
        RECT 2403.140 1015.280 2403.400 1015.540 ;
        RECT 1707.620 1014.940 1707.880 1015.200 ;
        RECT 1766.500 1014.940 1766.760 1015.200 ;
        RECT 2276.640 1014.940 2276.900 1015.200 ;
        RECT 2622.100 1014.940 2622.360 1015.200 ;
        RECT 1400.340 1014.600 1400.600 1014.860 ;
        RECT 1787.200 1014.600 1787.460 1014.860 ;
        RECT 2262.840 1014.600 2263.100 1014.860 ;
        RECT 2649.700 1014.600 2649.960 1014.860 ;
        RECT 1579.740 1014.260 1580.000 1014.520 ;
        RECT 1711.300 1014.260 1711.560 1014.520 ;
        RECT 1710.840 1013.920 1711.100 1014.180 ;
        RECT 1746.720 1014.260 1746.980 1014.520 ;
        RECT 2283.080 1014.260 2283.340 1014.520 ;
        RECT 2601.400 1014.260 2601.660 1014.520 ;
        RECT 2049.400 1013.920 2049.660 1014.180 ;
        RECT 2052.620 1013.920 2052.880 1014.180 ;
        RECT 1938.540 1010.860 1938.800 1011.120 ;
        RECT 2501.120 1010.860 2501.380 1011.120 ;
        RECT 1910.940 1010.520 1911.200 1010.780 ;
        RECT 2498.820 1010.520 2499.080 1010.780 ;
        RECT 2052.620 1007.800 2052.880 1008.060 ;
        RECT 2501.580 1007.800 2501.840 1008.060 ;
        RECT 2238.920 1005.760 2239.180 1006.020 ;
        RECT 2498.360 1005.760 2498.620 1006.020 ;
        RECT 1897.140 1005.420 1897.400 1005.680 ;
        RECT 2499.280 1005.420 2499.540 1005.680 ;
        RECT 1890.240 1005.080 1890.500 1005.340 ;
        RECT 2499.740 1005.080 2500.000 1005.340 ;
        RECT 1876.440 1004.740 1876.700 1005.000 ;
        RECT 2500.200 1004.740 2500.460 1005.000 ;
        RECT 1862.640 1004.400 1862.900 1004.660 ;
        RECT 2500.660 1004.400 2500.920 1004.660 ;
        RECT 1898.980 917.360 1899.240 917.620 ;
        RECT 2052.620 917.360 2052.880 917.620 ;
        RECT 1900.360 689.560 1900.620 689.820 ;
        RECT 1900.820 689.560 1901.080 689.820 ;
        RECT 1898.980 675.960 1899.240 676.220 ;
        RECT 1900.360 675.960 1900.620 676.220 ;
        RECT 1904.040 620.540 1904.300 620.800 ;
        RECT 1959.700 620.540 1959.960 620.800 ;
        RECT 1904.040 591.980 1904.300 592.240 ;
        RECT 1942.220 591.980 1942.480 592.240 ;
        RECT 1903.580 579.400 1903.840 579.660 ;
        RECT 1969.820 579.400 1970.080 579.660 ;
        RECT 1904.040 579.060 1904.300 579.320 ;
        RECT 1956.020 579.060 1956.280 579.320 ;
        RECT 1503.840 554.580 1504.100 554.840 ;
        RECT 2083.900 554.580 2084.160 554.840 ;
      LAYER met2 ;
        RECT 2442.700 3066.810 2442.960 3067.130 ;
        RECT 2469.840 3066.810 2470.100 3067.130 ;
        RECT 2442.760 3064.070 2442.900 3066.810 ;
        RECT 2469.900 3064.070 2470.040 3066.810 ;
        RECT 1868.160 3063.925 1868.420 3064.070 ;
        RECT 1868.150 3063.555 1868.430 3063.925 ;
        RECT 1898.060 3063.750 1898.320 3064.070 ;
        RECT 2442.700 3063.925 2442.960 3064.070 ;
        RECT 2469.840 3063.925 2470.100 3064.070 ;
        RECT 1490.030 3032.955 1490.310 3033.325 ;
        RECT 1489.570 3026.835 1489.850 3027.205 ;
        RECT 1489.110 3018.675 1489.390 3019.045 ;
        RECT 1488.650 3012.555 1488.930 3012.925 ;
        RECT 1488.190 3004.395 1488.470 3004.765 ;
        RECT 1487.730 2998.955 1488.010 2999.325 ;
        RECT 1487.270 2990.115 1487.550 2990.485 ;
        RECT 1486.810 2701.115 1487.090 2701.485 ;
        RECT 1486.350 2692.275 1486.630 2692.645 ;
        RECT 1486.420 2604.730 1486.560 2692.275 ;
        RECT 1486.360 2604.410 1486.620 2604.730 ;
        RECT 1448.640 2593.870 1448.900 2594.190 ;
        RECT 1372.740 2592.170 1373.000 2592.490 ;
        RECT 1358.940 2591.490 1359.200 2591.810 ;
        RECT 1345.140 2591.150 1345.400 2591.470 ;
        RECT 1331.340 2587.410 1331.600 2587.730 ;
        RECT 1306.040 2411.290 1306.300 2411.610 ;
        RECT 1306.100 2400.000 1306.240 2411.290 ;
        RECT 1318.450 2410.755 1318.730 2411.125 ;
        RECT 1318.520 2400.000 1318.660 2410.755 ;
        RECT 1331.400 2400.000 1331.540 2587.410 ;
        RECT 1306.070 2396.000 1306.350 2400.000 ;
        RECT 1318.490 2396.000 1318.770 2400.000 ;
        RECT 1331.370 2396.000 1331.650 2400.000 ;
        RECT 1344.250 2399.450 1344.530 2400.000 ;
        RECT 1345.200 2399.450 1345.340 2591.150 ;
        RECT 1344.250 2399.310 1345.340 2399.450 ;
        RECT 1357.130 2399.450 1357.410 2400.000 ;
        RECT 1359.000 2399.450 1359.140 2591.490 ;
        RECT 1357.130 2399.310 1359.140 2399.450 ;
        RECT 1344.250 2396.000 1344.530 2399.310 ;
        RECT 1357.130 2396.000 1357.410 2399.310 ;
        RECT 1370.010 2398.770 1370.290 2400.000 ;
        RECT 1372.800 2398.770 1372.940 2592.170 ;
        RECT 1434.840 2590.470 1435.100 2590.790 ;
        RECT 1427.940 2590.130 1428.200 2590.450 ;
        RECT 1414.140 2589.790 1414.400 2590.110 ;
        RECT 1400.340 2589.450 1400.600 2589.770 ;
        RECT 1386.540 2589.110 1386.800 2589.430 ;
        RECT 1386.600 2410.250 1386.740 2589.110 ;
        RECT 1400.400 2412.970 1400.540 2589.450 ;
        RECT 1414.200 2415.010 1414.340 2589.790 ;
        RECT 1408.620 2414.690 1408.880 2415.010 ;
        RECT 1414.140 2414.690 1414.400 2415.010 ;
        RECT 1395.740 2412.650 1396.000 2412.970 ;
        RECT 1400.340 2412.650 1400.600 2412.970 ;
        RECT 1382.860 2409.930 1383.120 2410.250 ;
        RECT 1386.540 2409.930 1386.800 2410.250 ;
        RECT 1382.920 2400.000 1383.060 2409.930 ;
        RECT 1395.800 2400.000 1395.940 2412.650 ;
        RECT 1408.680 2400.000 1408.820 2414.690 ;
        RECT 1428.000 2413.650 1428.140 2590.130 ;
        RECT 1421.500 2413.330 1421.760 2413.650 ;
        RECT 1427.940 2413.330 1428.200 2413.650 ;
        RECT 1421.560 2400.000 1421.700 2413.330 ;
        RECT 1370.010 2398.630 1372.940 2398.770 ;
        RECT 1370.010 2396.000 1370.290 2398.630 ;
        RECT 1382.890 2396.000 1383.170 2400.000 ;
        RECT 1395.770 2396.000 1396.050 2400.000 ;
        RECT 1408.650 2396.000 1408.930 2400.000 ;
        RECT 1421.530 2396.000 1421.810 2400.000 ;
        RECT 1434.410 2399.450 1434.690 2400.000 ;
        RECT 1434.900 2399.450 1435.040 2590.470 ;
        RECT 1434.410 2399.310 1435.040 2399.450 ;
        RECT 1447.290 2399.450 1447.570 2400.000 ;
        RECT 1448.700 2399.450 1448.840 2593.870 ;
        RECT 1486.880 2411.950 1487.020 2701.115 ;
        RECT 1487.340 2414.330 1487.480 2990.115 ;
        RECT 1487.280 2414.010 1487.540 2414.330 ;
        RECT 1487.800 2413.990 1487.940 2998.955 ;
        RECT 1487.740 2413.670 1488.000 2413.990 ;
        RECT 1488.260 2413.650 1488.400 3004.395 ;
        RECT 1488.200 2413.330 1488.460 2413.650 ;
        RECT 1488.720 2413.310 1488.860 3012.555 ;
        RECT 1488.660 2412.990 1488.920 2413.310 ;
        RECT 1489.180 2412.970 1489.320 3018.675 ;
        RECT 1489.120 2412.650 1489.380 2412.970 ;
        RECT 1489.640 2412.630 1489.780 3026.835 ;
        RECT 1489.580 2412.310 1489.840 2412.630 ;
        RECT 1490.100 2412.290 1490.240 3032.955 ;
      LAYER met2 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
      LAYER met2 ;
        RECT 1897.140 3008.330 1897.400 3008.650 ;
        RECT 1890.240 3001.530 1890.500 3001.850 ;
        RECT 1600.440 2594.210 1600.700 2594.530 ;
        RECT 1600.500 2594.045 1600.640 2594.210 ;
        RECT 1636.840 2594.190 1636.980 2594.345 ;
        RECT 1644.600 2594.210 1644.860 2594.530 ;
        RECT 1648.280 2594.210 1648.540 2594.530 ;
        RECT 1744.880 2594.210 1745.140 2594.530 ;
        RECT 1614.700 2594.045 1614.960 2594.190 ;
        RECT 1636.780 2594.045 1637.040 2594.190 ;
        RECT 1644.660 2594.045 1644.800 2594.210 ;
        RECT 1538.340 2593.530 1538.600 2593.850 ;
        RECT 1572.830 2593.675 1573.110 2594.045 ;
        RECT 1600.430 2593.675 1600.710 2594.045 ;
        RECT 1614.690 2593.675 1614.970 2594.045 ;
        RECT 1621.590 2593.675 1621.870 2594.045 ;
        RECT 1627.110 2593.675 1627.390 2594.045 ;
        RECT 1632.170 2593.675 1632.450 2594.045 ;
        RECT 1636.770 2593.675 1637.050 2594.045 ;
        RECT 1644.590 2593.675 1644.870 2594.045 ;
        RECT 1524.540 2588.090 1524.800 2588.410 ;
        RECT 1490.040 2411.970 1490.300 2412.290 ;
        RECT 1486.820 2411.630 1487.080 2411.950 ;
        RECT 1460.140 2409.930 1460.400 2410.250 ;
        RECT 1460.200 2400.000 1460.340 2409.930 ;
        RECT 1472.560 2409.590 1472.820 2409.910 ;
        RECT 1472.620 2400.000 1472.760 2409.590 ;
        RECT 1485.440 2409.250 1485.700 2409.570 ;
        RECT 1485.500 2400.000 1485.640 2409.250 ;
        RECT 1498.320 2408.910 1498.580 2409.230 ;
        RECT 1498.380 2400.000 1498.520 2408.910 ;
        RECT 1511.200 2408.570 1511.460 2408.890 ;
        RECT 1511.260 2400.000 1511.400 2408.570 ;
        RECT 1447.290 2399.310 1448.840 2399.450 ;
        RECT 1434.410 2396.000 1434.690 2399.310 ;
        RECT 1447.290 2396.000 1447.570 2399.310 ;
        RECT 1460.170 2396.000 1460.450 2400.000 ;
        RECT 1472.590 2396.000 1472.870 2400.000 ;
        RECT 1485.470 2396.000 1485.750 2400.000 ;
        RECT 1498.350 2396.000 1498.630 2400.000 ;
        RECT 1511.230 2396.000 1511.510 2400.000 ;
        RECT 1524.110 2399.450 1524.390 2400.000 ;
        RECT 1524.600 2399.450 1524.740 2588.090 ;
        RECT 1537.870 2587.555 1538.150 2587.925 ;
        RECT 1537.940 2414.670 1538.080 2587.555 ;
        RECT 1537.880 2414.350 1538.140 2414.670 ;
        RECT 1524.110 2399.310 1524.740 2399.450 ;
        RECT 1536.990 2399.450 1537.270 2400.000 ;
        RECT 1538.400 2399.450 1538.540 2593.530 ;
        RECT 1572.900 2593.510 1573.040 2593.675 ;
        RECT 1565.930 2592.995 1566.210 2593.365 ;
        RECT 1572.840 2593.190 1573.100 2593.510 ;
        RECT 1615.620 2593.365 1615.880 2593.510 ;
        RECT 1586.170 2592.995 1586.450 2593.365 ;
        RECT 1593.530 2592.995 1593.810 2593.365 ;
        RECT 1605.490 2592.995 1605.770 2593.365 ;
        RECT 1615.610 2592.995 1615.890 2593.365 ;
        RECT 1566.000 2592.150 1566.140 2592.995 ;
        RECT 1573.290 2592.315 1573.570 2592.685 ;
        RECT 1580.190 2592.315 1580.470 2592.685 ;
        RECT 1565.940 2591.830 1566.200 2592.150 ;
        RECT 1566.390 2591.635 1566.670 2592.005 ;
        RECT 1573.360 2591.810 1573.500 2592.315 ;
        RECT 1580.200 2592.170 1580.460 2592.315 ;
        RECT 1586.240 2592.150 1586.380 2592.995 ;
        RECT 1593.540 2592.850 1593.800 2592.995 ;
        RECT 1605.560 2592.830 1605.700 2592.995 ;
        RECT 1586.630 2592.315 1586.910 2592.685 ;
        RECT 1587.550 2592.315 1587.830 2592.685 ;
        RECT 1605.500 2592.510 1605.760 2592.830 ;
        RECT 1586.640 2592.170 1586.900 2592.315 ;
        RECT 1586.180 2591.830 1586.440 2592.150 ;
        RECT 1566.460 2591.470 1566.600 2591.635 ;
        RECT 1573.300 2591.490 1573.560 2591.810 ;
        RECT 1566.400 2591.150 1566.660 2591.470 ;
        RECT 1579.280 2591.150 1579.540 2591.470 ;
        RECT 1579.340 2590.450 1579.480 2591.150 ;
        RECT 1579.280 2590.130 1579.540 2590.450 ;
        RECT 1579.730 2590.275 1580.010 2590.645 ;
        RECT 1579.740 2590.130 1580.000 2590.275 ;
        RECT 1587.090 2589.595 1587.370 2589.965 ;
        RECT 1587.620 2589.770 1587.760 2592.315 ;
        RECT 1593.990 2591.635 1594.270 2592.005 ;
        RECT 1600.890 2591.635 1601.170 2592.005 ;
        RECT 1594.000 2591.490 1594.260 2591.635 ;
        RECT 1600.960 2591.470 1601.100 2591.635 ;
        RECT 1600.900 2591.150 1601.160 2591.470 ;
        RECT 1608.710 2590.955 1608.990 2591.325 ;
        RECT 1608.780 2590.790 1608.920 2590.955 ;
        RECT 1593.990 2590.275 1594.270 2590.645 ;
        RECT 1608.720 2590.470 1608.980 2590.790 ;
        RECT 1621.660 2590.450 1621.800 2593.675 ;
        RECT 1627.180 2592.150 1627.320 2593.675 ;
        RECT 1627.570 2592.315 1627.850 2592.685 ;
        RECT 1632.240 2592.490 1632.380 2593.675 ;
        RECT 1636.840 2593.170 1636.980 2593.675 ;
        RECT 1648.340 2593.170 1648.480 2594.210 ;
        RECT 1684.620 2594.045 1684.880 2594.190 ;
        RECT 1726.480 2594.045 1726.740 2594.190 ;
        RECT 1744.940 2594.045 1745.080 2594.210 ;
        RECT 1650.570 2593.675 1650.850 2594.045 ;
        RECT 1656.550 2593.675 1656.830 2594.045 ;
        RECT 1636.780 2592.850 1637.040 2593.170 ;
        RECT 1648.280 2592.850 1648.540 2593.170 ;
        RECT 1650.640 2592.830 1650.780 2593.675 ;
        RECT 1656.560 2593.530 1656.820 2593.675 ;
        RECT 1657.020 2593.530 1657.280 2593.850 ;
        RECT 1662.070 2593.675 1662.350 2594.045 ;
        RECT 1668.970 2593.675 1669.250 2594.045 ;
        RECT 1673.570 2593.675 1673.850 2594.045 ;
        RECT 1679.090 2593.675 1679.370 2594.045 ;
        RECT 1684.610 2593.675 1684.890 2594.045 ;
        RECT 1690.590 2593.675 1690.870 2594.045 ;
        RECT 1697.490 2593.675 1697.770 2594.045 ;
        RECT 1703.010 2593.675 1703.290 2594.045 ;
        RECT 1707.610 2593.675 1707.890 2594.045 ;
        RECT 1726.470 2593.675 1726.750 2594.045 ;
        RECT 1732.910 2593.675 1733.190 2594.045 ;
        RECT 1744.870 2593.675 1745.150 2594.045 ;
        RECT 1657.080 2593.365 1657.220 2593.530 ;
        RECT 1662.140 2593.510 1662.280 2593.675 ;
        RECT 1657.010 2592.995 1657.290 2593.365 ;
        RECT 1662.080 2593.190 1662.340 2593.510 ;
        RECT 1627.640 2592.150 1627.780 2592.315 ;
        RECT 1632.180 2592.170 1632.440 2592.490 ;
        RECT 1649.190 2592.315 1649.470 2592.685 ;
        RECT 1650.580 2592.510 1650.840 2592.830 ;
        RECT 1627.120 2591.830 1627.380 2592.150 ;
        RECT 1627.580 2591.830 1627.840 2592.150 ;
        RECT 1627.180 2591.470 1627.320 2591.830 ;
        RECT 1627.120 2591.150 1627.380 2591.470 ;
        RECT 1594.060 2590.110 1594.200 2590.275 ;
        RECT 1621.600 2590.130 1621.860 2590.450 ;
        RECT 1627.580 2590.130 1627.840 2590.450 ;
        RECT 1628.040 2590.130 1628.300 2590.450 ;
        RECT 1594.000 2589.790 1594.260 2590.110 ;
        RECT 1587.160 2589.430 1587.300 2589.595 ;
        RECT 1587.560 2589.450 1587.820 2589.770 ;
        RECT 1614.240 2589.450 1614.500 2589.770 ;
        RECT 1560.870 2588.915 1561.150 2589.285 ;
        RECT 1587.100 2589.110 1587.360 2589.430 ;
        RECT 1607.340 2589.110 1607.600 2589.430 ;
        RECT 1551.210 2588.235 1551.490 2588.605 ;
        RECT 1545.230 2587.555 1545.510 2587.925 ;
        RECT 1545.300 2410.590 1545.440 2587.555 ;
        RECT 1551.280 2410.930 1551.420 2588.235 ;
        RECT 1551.670 2587.555 1551.950 2587.925 ;
        RECT 1552.140 2587.750 1552.400 2588.070 ;
        RECT 1551.740 2411.270 1551.880 2587.555 ;
        RECT 1551.680 2410.950 1551.940 2411.270 ;
        RECT 1551.220 2410.610 1551.480 2410.930 ;
        RECT 1545.240 2410.270 1545.500 2410.590 ;
        RECT 1536.990 2399.310 1538.540 2399.450 ;
        RECT 1549.870 2399.450 1550.150 2400.000 ;
        RECT 1552.200 2399.450 1552.340 2587.750 ;
        RECT 1559.030 2587.555 1559.310 2587.925 ;
        RECT 1560.940 2587.730 1561.080 2588.915 ;
        RECT 1579.740 2588.770 1580.000 2589.090 ;
        RECT 1565.940 2588.430 1566.200 2588.750 ;
        RECT 1559.100 2415.010 1559.240 2587.555 ;
        RECT 1560.880 2587.410 1561.140 2587.730 ;
        RECT 1559.040 2414.690 1559.300 2415.010 ;
        RECT 1549.870 2399.310 1552.340 2399.450 ;
        RECT 1524.110 2396.000 1524.390 2399.310 ;
        RECT 1536.990 2396.000 1537.270 2399.310 ;
        RECT 1549.870 2396.000 1550.150 2399.310 ;
        RECT 1562.750 2398.770 1563.030 2400.000 ;
        RECT 1566.000 2398.770 1566.140 2588.430 ;
        RECT 1579.800 2408.550 1579.940 2588.770 ;
        RECT 1600.890 2410.075 1601.170 2410.445 ;
        RECT 1607.400 2410.250 1607.540 2589.110 ;
        RECT 1600.900 2409.930 1601.160 2410.075 ;
        RECT 1601.360 2409.930 1601.620 2410.250 ;
        RECT 1607.340 2409.930 1607.600 2410.250 ;
        RECT 1607.790 2410.075 1608.070 2410.445 ;
        RECT 1607.800 2409.930 1608.060 2410.075 ;
        RECT 1575.600 2408.230 1575.860 2408.550 ;
        RECT 1579.740 2408.230 1580.000 2408.550 ;
        RECT 1588.480 2408.230 1588.740 2408.550 ;
        RECT 1575.660 2400.000 1575.800 2408.230 ;
        RECT 1588.540 2400.000 1588.680 2408.230 ;
        RECT 1601.420 2400.000 1601.560 2409.930 ;
        RECT 1614.300 2400.000 1614.440 2589.450 ;
        RECT 1622.510 2588.235 1622.790 2588.605 ;
        RECT 1622.050 2587.555 1622.330 2587.925 ;
        RECT 1622.120 2409.910 1622.260 2587.555 ;
        RECT 1622.580 2410.250 1622.720 2588.235 ;
        RECT 1627.640 2587.730 1627.780 2590.130 ;
        RECT 1627.580 2587.410 1627.840 2587.730 ;
        RECT 1622.520 2409.930 1622.780 2410.250 ;
        RECT 1622.060 2409.590 1622.320 2409.910 ;
        RECT 1562.750 2398.630 1566.140 2398.770 ;
        RECT 1562.750 2396.000 1563.030 2398.630 ;
        RECT 1575.630 2396.000 1575.910 2400.000 ;
        RECT 1588.510 2396.000 1588.790 2400.000 ;
        RECT 1601.390 2396.000 1601.670 2400.000 ;
        RECT 1614.270 2396.000 1614.550 2400.000 ;
        RECT 1626.690 2399.450 1626.970 2400.000 ;
        RECT 1628.100 2399.450 1628.240 2590.130 ;
        RECT 1641.840 2589.790 1642.100 2590.110 ;
        RECT 1628.490 2588.235 1628.770 2588.605 ;
        RECT 1635.850 2588.235 1636.130 2588.605 ;
        RECT 1628.560 2409.570 1628.700 2588.235 ;
        RECT 1628.960 2409.590 1629.220 2409.910 ;
        RECT 1628.500 2409.250 1628.760 2409.570 ;
        RECT 1628.500 2408.460 1628.760 2408.550 ;
        RECT 1629.020 2408.460 1629.160 2409.590 ;
        RECT 1635.920 2409.230 1636.060 2588.235 ;
        RECT 1635.860 2408.910 1636.120 2409.230 ;
        RECT 1628.500 2408.320 1629.160 2408.460 ;
        RECT 1628.500 2408.230 1628.760 2408.320 ;
        RECT 1626.690 2399.310 1628.240 2399.450 ;
        RECT 1626.690 2396.000 1626.970 2399.310 ;
        RECT 1639.570 2398.770 1639.850 2400.000 ;
        RECT 1641.900 2398.770 1642.040 2589.790 ;
        RECT 1642.290 2588.235 1642.570 2588.605 ;
        RECT 1649.260 2588.410 1649.400 2592.315 ;
        RECT 1657.080 2592.150 1657.220 2592.995 ;
        RECT 1669.040 2592.150 1669.180 2593.675 ;
        RECT 1657.020 2591.830 1657.280 2592.150 ;
        RECT 1668.980 2591.830 1669.240 2592.150 ;
        RECT 1663.450 2590.955 1663.730 2591.325 ;
        RECT 1655.640 2590.470 1655.900 2590.790 ;
        RECT 1642.360 2408.890 1642.500 2588.235 ;
        RECT 1649.200 2588.090 1649.460 2588.410 ;
        RECT 1642.300 2408.570 1642.560 2408.890 ;
        RECT 1639.570 2398.630 1642.040 2398.770 ;
        RECT 1652.450 2398.770 1652.730 2400.000 ;
        RECT 1655.700 2398.770 1655.840 2590.470 ;
        RECT 1663.520 2588.750 1663.660 2590.955 ;
        RECT 1662.990 2588.235 1663.270 2588.605 ;
        RECT 1663.460 2588.430 1663.720 2588.750 ;
        RECT 1663.060 2588.070 1663.200 2588.235 ;
        RECT 1663.000 2587.750 1663.260 2588.070 ;
        RECT 1669.040 2587.730 1669.180 2591.830 ;
        RECT 1673.640 2591.470 1673.780 2593.675 ;
        RECT 1679.160 2592.490 1679.300 2593.675 ;
        RECT 1679.100 2592.170 1679.360 2592.490 ;
        RECT 1683.690 2591.635 1683.970 2592.005 ;
        RECT 1684.680 2591.810 1684.820 2593.675 ;
        RECT 1690.660 2593.170 1690.800 2593.675 ;
        RECT 1690.600 2592.850 1690.860 2593.170 ;
        RECT 1697.560 2592.830 1697.700 2593.675 ;
        RECT 1703.020 2593.530 1703.280 2593.675 ;
        RECT 1697.950 2592.995 1698.230 2593.365 ;
        RECT 1697.500 2592.510 1697.760 2592.830 ;
        RECT 1673.580 2591.150 1673.840 2591.470 ;
        RECT 1683.760 2589.430 1683.900 2591.635 ;
        RECT 1684.620 2591.490 1684.880 2591.810 ;
        RECT 1690.590 2591.635 1690.870 2592.005 ;
        RECT 1697.490 2591.635 1697.770 2592.005 ;
        RECT 1690.660 2589.770 1690.800 2591.635 ;
        RECT 1697.560 2590.450 1697.700 2591.635 ;
        RECT 1697.500 2590.130 1697.760 2590.450 ;
        RECT 1698.020 2590.110 1698.160 2592.995 ;
        RECT 1703.080 2590.110 1703.220 2593.530 ;
        RECT 1707.680 2593.510 1707.820 2593.675 ;
        RECT 1707.620 2593.190 1707.880 2593.510 ;
        RECT 1704.390 2590.955 1704.670 2591.325 ;
        RECT 1704.460 2590.790 1704.600 2590.955 ;
        RECT 1704.400 2590.470 1704.660 2590.790 ;
        RECT 1697.960 2589.790 1698.220 2590.110 ;
        RECT 1703.020 2589.790 1703.280 2590.110 ;
        RECT 1707.680 2589.770 1707.820 2593.190 ;
        RECT 1714.970 2592.315 1715.250 2592.685 ;
        RECT 1726.540 2592.490 1726.680 2593.675 ;
        RECT 1732.920 2593.530 1733.180 2593.675 ;
        RECT 1715.040 2592.150 1715.180 2592.315 ;
        RECT 1726.480 2592.170 1726.740 2592.490 ;
        RECT 1714.980 2591.830 1715.240 2592.150 ;
        RECT 1690.600 2589.450 1690.860 2589.770 ;
        RECT 1707.620 2589.450 1707.880 2589.770 ;
        RECT 1715.040 2589.430 1715.180 2591.830 ;
        RECT 1718.650 2591.635 1718.930 2592.005 ;
        RECT 1732.980 2591.810 1733.120 2593.530 ;
        RECT 1738.430 2592.995 1738.710 2593.365 ;
        RECT 1738.440 2592.850 1738.700 2592.995 ;
        RECT 1744.940 2592.830 1745.080 2593.675 ;
        RECT 1738.890 2592.315 1739.170 2592.685 ;
        RECT 1744.880 2592.510 1745.140 2592.830 ;
        RECT 1718.720 2591.470 1718.860 2591.635 ;
        RECT 1732.920 2591.490 1733.180 2591.810 ;
        RECT 1718.660 2591.150 1718.920 2591.470 ;
        RECT 1721.880 2591.150 1722.140 2591.470 ;
        RECT 1669.890 2588.915 1670.170 2589.285 ;
        RECT 1683.700 2589.110 1683.960 2589.430 ;
        RECT 1711.290 2588.915 1711.570 2589.285 ;
        RECT 1714.980 2589.110 1715.240 2589.430 ;
        RECT 1721.940 2589.090 1722.080 2591.150 ;
        RECT 1669.900 2588.770 1670.160 2588.915 ;
        RECT 1711.360 2588.750 1711.500 2588.915 ;
        RECT 1721.880 2588.770 1722.140 2589.090 ;
        RECT 1669.440 2588.430 1669.700 2588.750 ;
        RECT 1668.980 2587.410 1669.240 2587.730 ;
        RECT 1669.500 2410.250 1669.640 2588.430 ;
        RECT 1676.790 2588.235 1677.070 2588.605 ;
        RECT 1711.300 2588.430 1711.560 2588.750 ;
        RECT 1665.300 2409.930 1665.560 2410.250 ;
        RECT 1669.440 2409.930 1669.700 2410.250 ;
        RECT 1665.360 2400.000 1665.500 2409.930 ;
        RECT 1676.860 2408.890 1677.000 2588.235 ;
        RECT 1686.920 2588.090 1687.180 2588.410 ;
        RECT 1718.190 2588.235 1718.470 2588.605 ;
        RECT 1721.420 2588.430 1721.680 2588.750 ;
        RECT 1718.200 2588.090 1718.460 2588.235 ;
        RECT 1686.980 2408.890 1687.120 2588.090 ;
        RECT 1703.940 2587.750 1704.200 2588.070 ;
        RECT 1697.040 2587.410 1697.300 2587.730 ;
        RECT 1697.100 2410.250 1697.240 2587.410 ;
        RECT 1691.060 2409.930 1691.320 2410.250 ;
        RECT 1697.040 2409.930 1697.300 2410.250 ;
        RECT 1676.800 2408.570 1677.060 2408.890 ;
        RECT 1678.180 2408.570 1678.440 2408.890 ;
        RECT 1686.920 2408.570 1687.180 2408.890 ;
        RECT 1678.240 2400.000 1678.380 2408.570 ;
        RECT 1691.120 2400.000 1691.260 2409.930 ;
        RECT 1704.000 2400.000 1704.140 2587.750 ;
        RECT 1721.480 2410.250 1721.620 2588.430 ;
        RECT 1726.010 2588.235 1726.290 2588.605 ;
        RECT 1731.990 2588.235 1732.270 2588.605 ;
        RECT 1726.080 2587.730 1726.220 2588.235 ;
        RECT 1732.060 2588.070 1732.200 2588.235 ;
        RECT 1732.000 2587.750 1732.260 2588.070 ;
        RECT 1738.960 2587.730 1739.100 2592.315 ;
        RECT 1848.840 2591.830 1849.100 2592.150 ;
        RECT 1786.740 2591.490 1787.000 2591.810 ;
        RECT 1772.940 2591.150 1773.200 2591.470 ;
        RECT 1759.140 2590.470 1759.400 2590.790 ;
        RECT 1745.340 2590.130 1745.600 2590.450 ;
        RECT 1739.350 2588.915 1739.630 2589.285 ;
        RECT 1739.420 2588.750 1739.560 2588.915 ;
        RECT 1739.360 2588.430 1739.620 2588.750 ;
        RECT 1726.020 2587.410 1726.280 2587.730 ;
        RECT 1731.540 2587.410 1731.800 2587.730 ;
        RECT 1738.900 2587.410 1739.160 2587.730 ;
        RECT 1716.820 2409.930 1717.080 2410.250 ;
        RECT 1721.420 2409.930 1721.680 2410.250 ;
        RECT 1716.880 2400.000 1717.020 2409.930 ;
        RECT 1652.450 2398.630 1655.840 2398.770 ;
        RECT 1639.570 2396.000 1639.850 2398.630 ;
        RECT 1652.450 2396.000 1652.730 2398.630 ;
        RECT 1665.330 2396.000 1665.610 2400.000 ;
        RECT 1678.210 2396.000 1678.490 2400.000 ;
        RECT 1691.090 2396.000 1691.370 2400.000 ;
        RECT 1703.970 2396.000 1704.250 2400.000 ;
        RECT 1716.850 2396.000 1717.130 2400.000 ;
        RECT 1729.730 2399.450 1730.010 2400.000 ;
        RECT 1731.600 2399.450 1731.740 2587.410 ;
        RECT 1729.730 2399.310 1731.740 2399.450 ;
        RECT 1729.730 2396.000 1730.010 2399.310 ;
        RECT 1742.610 2398.770 1742.890 2400.000 ;
        RECT 1745.400 2398.770 1745.540 2590.130 ;
        RECT 1759.200 2410.250 1759.340 2590.470 ;
        RECT 1773.000 2410.250 1773.140 2591.150 ;
        RECT 1755.460 2409.930 1755.720 2410.250 ;
        RECT 1759.140 2409.930 1759.400 2410.250 ;
        RECT 1768.340 2409.930 1768.600 2410.250 ;
        RECT 1772.940 2409.930 1773.200 2410.250 ;
        RECT 1755.520 2400.000 1755.660 2409.930 ;
        RECT 1768.400 2400.000 1768.540 2409.930 ;
        RECT 1786.800 2409.570 1786.940 2591.490 ;
        RECT 1832.280 2414.690 1832.540 2415.010 ;
        RECT 1819.400 2410.950 1819.660 2411.270 ;
        RECT 1806.520 2410.610 1806.780 2410.930 ;
        RECT 1793.640 2410.270 1793.900 2410.590 ;
        RECT 1780.760 2409.250 1781.020 2409.570 ;
        RECT 1786.740 2409.250 1787.000 2409.570 ;
        RECT 1780.820 2400.000 1780.960 2409.250 ;
        RECT 1793.700 2400.000 1793.840 2410.270 ;
        RECT 1806.580 2400.000 1806.720 2410.610 ;
        RECT 1819.460 2400.000 1819.600 2410.950 ;
        RECT 1832.340 2400.000 1832.480 2414.690 ;
        RECT 1742.610 2398.630 1745.540 2398.770 ;
        RECT 1742.610 2396.000 1742.890 2398.630 ;
        RECT 1755.490 2396.000 1755.770 2400.000 ;
        RECT 1768.370 2396.000 1768.650 2400.000 ;
        RECT 1780.790 2396.000 1781.070 2400.000 ;
        RECT 1793.670 2396.000 1793.950 2400.000 ;
        RECT 1806.550 2396.000 1806.830 2400.000 ;
        RECT 1819.430 2396.000 1819.710 2400.000 ;
        RECT 1832.310 2396.000 1832.590 2400.000 ;
        RECT 1845.190 2398.770 1845.470 2400.000 ;
        RECT 1848.900 2398.770 1849.040 2591.830 ;
        RECT 1858.040 2414.690 1858.300 2415.010 ;
        RECT 1858.100 2400.000 1858.240 2414.690 ;
        RECT 1890.300 2411.610 1890.440 3001.530 ;
        RECT 1883.800 2411.290 1884.060 2411.610 ;
        RECT 1890.240 2411.290 1890.500 2411.610 ;
        RECT 1870.920 2410.950 1871.180 2411.270 ;
        RECT 1870.980 2400.000 1871.120 2410.950 ;
        RECT 1883.860 2400.000 1884.000 2411.290 ;
        RECT 1845.190 2398.630 1849.040 2398.770 ;
        RECT 1845.190 2396.000 1845.470 2398.630 ;
        RECT 1858.070 2396.000 1858.350 2400.000 ;
        RECT 1870.950 2396.000 1871.230 2400.000 ;
        RECT 1883.830 2396.000 1884.110 2400.000 ;
        RECT 1896.710 2399.450 1896.990 2400.000 ;
        RECT 1897.200 2399.450 1897.340 3008.330 ;
        RECT 1898.120 2747.045 1898.260 3063.750 ;
        RECT 2442.690 3063.555 2442.970 3063.925 ;
        RECT 2469.830 3063.555 2470.110 3063.925 ;
        RECT 2497.900 3063.750 2498.160 3064.070 ;
        RECT 1899.900 3051.850 1900.160 3052.170 ;
        RECT 2482.260 3051.850 2482.520 3052.170 ;
        RECT 1899.960 3048.285 1900.100 3051.850 ;
        RECT 1898.510 3047.915 1898.790 3048.285 ;
        RECT 1899.890 3047.915 1900.170 3048.285 ;
        RECT 1898.050 2746.675 1898.330 2747.045 ;
        RECT 1897.600 2691.110 1897.860 2691.430 ;
        RECT 1897.660 2680.550 1897.800 2691.110 ;
        RECT 1897.600 2680.230 1897.860 2680.550 ;
        RECT 1898.060 2594.550 1898.320 2594.870 ;
        RECT 1898.120 2570.390 1898.260 2594.550 ;
        RECT 1898.060 2570.070 1898.320 2570.390 ;
        RECT 1898.060 2497.650 1898.320 2497.970 ;
        RECT 1898.120 2473.830 1898.260 2497.650 ;
        RECT 1898.060 2473.510 1898.320 2473.830 ;
        RECT 1898.580 2411.125 1898.720 3047.915 ;
        RECT 2083.890 3030.235 2084.170 3030.605 ;
        RECT 2083.960 3029.390 2084.100 3030.235 ;
        RECT 1938.540 3029.070 1938.800 3029.390 ;
        RECT 2083.900 3029.070 2084.160 3029.390 ;
        RECT 1924.740 3022.270 1925.000 3022.590 ;
        RECT 1910.940 3015.470 1911.200 3015.790 ;
        RECT 1898.970 2704.515 1899.250 2704.885 ;
        RECT 1899.040 2691.430 1899.180 2704.515 ;
        RECT 1898.980 2691.110 1899.240 2691.430 ;
        RECT 1898.980 2680.230 1899.240 2680.550 ;
        RECT 1899.040 2594.870 1899.180 2680.230 ;
        RECT 1898.980 2594.550 1899.240 2594.870 ;
        RECT 1898.980 2570.070 1899.240 2570.390 ;
        RECT 1899.040 2497.970 1899.180 2570.070 ;
        RECT 1898.980 2497.650 1899.240 2497.970 ;
        RECT 1898.980 2473.510 1899.240 2473.830 ;
        RECT 1898.510 2410.755 1898.790 2411.125 ;
        RECT 1899.040 2410.590 1899.180 2473.510 ;
        RECT 1898.980 2410.270 1899.240 2410.590 ;
        RECT 1896.710 2399.310 1897.340 2399.450 ;
        RECT 1909.590 2399.450 1909.870 2400.000 ;
        RECT 1911.000 2399.450 1911.140 3015.470 ;
        RECT 1909.590 2399.310 1911.140 2399.450 ;
        RECT 1922.470 2399.450 1922.750 2400.000 ;
        RECT 1924.800 2399.450 1924.940 3022.270 ;
        RECT 1938.600 2414.670 1938.740 3029.070 ;
        RECT 2083.890 3024.115 2084.170 3024.485 ;
        RECT 2083.960 3022.590 2084.100 3024.115 ;
        RECT 2083.900 3022.270 2084.160 3022.590 ;
        RECT 2083.890 3015.955 2084.170 3016.325 ;
        RECT 2083.960 3015.790 2084.100 3015.955 ;
        RECT 2083.900 3015.470 2084.160 3015.790 ;
        RECT 2083.890 3009.835 2084.170 3010.205 ;
        RECT 2083.960 3008.650 2084.100 3009.835 ;
        RECT 2083.900 3008.330 2084.160 3008.650 ;
        RECT 2083.890 3002.355 2084.170 3002.725 ;
        RECT 2083.960 3001.850 2084.100 3002.355 ;
        RECT 2083.900 3001.530 2084.160 3001.850 ;
        RECT 2087.110 2996.235 2087.390 2996.605 ;
        RECT 2084.810 2698.395 2085.090 2698.765 ;
        RECT 2084.880 2698.230 2085.020 2698.395 ;
        RECT 2069.640 2697.910 2069.900 2698.230 ;
        RECT 2084.820 2697.910 2085.080 2698.230 ;
        RECT 2052.620 2691.110 2052.880 2691.430 ;
        RECT 2052.680 2608.130 2052.820 2691.110 ;
        RECT 2049.400 2607.810 2049.660 2608.130 ;
        RECT 2052.620 2607.810 2052.880 2608.130 ;
        RECT 2049.460 2604.730 2049.600 2607.810 ;
        RECT 2049.400 2604.410 2049.660 2604.730 ;
        RECT 1934.860 2414.350 1935.120 2414.670 ;
        RECT 1938.540 2414.350 1938.800 2414.670 ;
        RECT 1932.560 2414.010 1932.820 2414.330 ;
        RECT 1932.620 2411.610 1932.760 2414.010 ;
        RECT 1932.560 2411.290 1932.820 2411.610 ;
        RECT 1934.920 2400.000 1935.060 2414.350 ;
        RECT 1947.740 2414.010 1948.000 2414.330 ;
        RECT 1947.800 2400.000 1947.940 2414.010 ;
        RECT 1973.500 2413.670 1973.760 2413.990 ;
        RECT 1960.620 2411.290 1960.880 2411.610 ;
        RECT 1960.680 2400.000 1960.820 2411.290 ;
        RECT 1973.560 2400.000 1973.700 2413.670 ;
        RECT 1986.380 2413.330 1986.640 2413.650 ;
        RECT 1986.440 2400.000 1986.580 2413.330 ;
        RECT 1999.260 2412.990 1999.520 2413.310 ;
        RECT 1999.320 2400.000 1999.460 2412.990 ;
        RECT 2012.140 2412.650 2012.400 2412.970 ;
        RECT 2012.200 2400.000 2012.340 2412.650 ;
        RECT 2025.020 2412.310 2025.280 2412.630 ;
        RECT 2025.080 2400.000 2025.220 2412.310 ;
        RECT 2037.900 2411.970 2038.160 2412.290 ;
        RECT 2037.960 2400.000 2038.100 2411.970 ;
        RECT 1922.470 2399.310 1924.940 2399.450 ;
        RECT 1896.710 2396.000 1896.990 2399.310 ;
        RECT 1909.590 2396.000 1909.870 2399.310 ;
        RECT 1922.470 2396.000 1922.750 2399.310 ;
        RECT 1934.890 2396.000 1935.170 2400.000 ;
        RECT 1947.770 2396.000 1948.050 2400.000 ;
        RECT 1960.650 2396.000 1960.930 2400.000 ;
        RECT 1973.530 2396.000 1973.810 2400.000 ;
        RECT 1986.410 2396.000 1986.690 2400.000 ;
        RECT 1999.290 2396.000 1999.570 2400.000 ;
        RECT 2012.170 2396.000 2012.450 2400.000 ;
        RECT 2025.050 2396.000 2025.330 2400.000 ;
        RECT 2037.930 2396.000 2038.210 2400.000 ;
        RECT 2049.460 2399.450 2049.600 2604.410 ;
        RECT 2069.700 2412.970 2069.840 2697.910 ;
        RECT 2083.890 2691.595 2084.170 2691.965 ;
        RECT 2083.960 2691.430 2084.100 2691.595 ;
        RECT 2083.900 2691.110 2084.160 2691.430 ;
        RECT 2063.660 2412.650 2063.920 2412.970 ;
        RECT 2069.640 2412.650 2069.900 2412.970 ;
        RECT 2063.720 2400.000 2063.860 2412.650 ;
        RECT 2076.540 2411.630 2076.800 2411.950 ;
        RECT 2076.600 2400.000 2076.740 2411.630 ;
        RECT 2087.180 2411.270 2087.320 2996.235 ;
        RECT 2087.570 2988.075 2087.850 2988.445 ;
        RECT 2087.640 2415.010 2087.780 2988.075 ;
      LAYER met2 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met2 ;
        RECT 2482.320 3049.645 2482.460 3051.850 ;
        RECT 2482.250 3049.275 2482.530 3049.645 ;
        RECT 2497.960 2747.725 2498.100 3063.750 ;
        RECT 2497.890 2747.355 2498.170 2747.725 ;
        RECT 2497.890 2709.955 2498.170 2710.325 ;
        RECT 2497.960 2704.885 2498.100 2709.955 ;
        RECT 2497.890 2704.515 2498.170 2704.885 ;
        RECT 2126.670 2598.435 2126.950 2598.805 ;
        RECT 2170.830 2598.435 2171.110 2598.805 ;
        RECT 2126.740 2590.450 2126.880 2598.435 ;
        RECT 2146.450 2592.995 2146.730 2593.365 ;
        RECT 2132.190 2592.315 2132.470 2592.685 ;
        RECT 2132.260 2592.150 2132.400 2592.315 ;
        RECT 2132.200 2591.830 2132.460 2592.150 ;
        RECT 2146.520 2591.470 2146.660 2592.995 ;
        RECT 2152.890 2591.635 2153.170 2592.005 ;
        RECT 2152.900 2591.490 2153.160 2591.635 ;
        RECT 2145.990 2590.955 2146.270 2591.325 ;
        RECT 2146.460 2591.150 2146.720 2591.470 ;
        RECT 2146.060 2590.790 2146.200 2590.955 ;
        RECT 2146.000 2590.470 2146.260 2590.790 ;
        RECT 2126.680 2590.130 2126.940 2590.450 ;
        RECT 2163.020 2590.130 2163.280 2590.450 ;
        RECT 2163.080 2589.285 2163.220 2590.130 ;
        RECT 2163.010 2588.915 2163.290 2589.285 ;
        RECT 2087.580 2414.690 2087.840 2415.010 ;
        RECT 2153.360 2413.670 2153.620 2413.990 ;
        RECT 2140.480 2413.330 2140.740 2413.650 ;
        RECT 2127.600 2412.990 2127.860 2413.310 ;
        RECT 2114.720 2412.650 2114.980 2412.970 ;
        RECT 2101.840 2411.630 2102.100 2411.950 ;
        RECT 2088.960 2411.290 2089.220 2411.610 ;
        RECT 2087.120 2410.950 2087.380 2411.270 ;
        RECT 2089.020 2400.000 2089.160 2411.290 ;
        RECT 2101.900 2400.000 2102.040 2411.630 ;
        RECT 2114.780 2400.000 2114.920 2412.650 ;
        RECT 2127.660 2400.000 2127.800 2412.990 ;
        RECT 2140.540 2400.000 2140.680 2413.330 ;
        RECT 2153.420 2400.000 2153.560 2413.670 ;
        RECT 2163.080 2411.610 2163.220 2588.915 ;
        RECT 2166.230 2588.235 2166.510 2588.605 ;
        RECT 2165.780 2414.690 2166.040 2415.010 ;
        RECT 2163.020 2411.290 2163.280 2411.610 ;
        RECT 2050.810 2399.450 2051.090 2400.000 ;
        RECT 2049.460 2399.310 2051.090 2399.450 ;
        RECT 2050.810 2396.000 2051.090 2399.310 ;
        RECT 2063.690 2396.000 2063.970 2400.000 ;
        RECT 2076.570 2396.000 2076.850 2400.000 ;
        RECT 2088.990 2396.000 2089.270 2400.000 ;
        RECT 2101.870 2396.000 2102.150 2400.000 ;
        RECT 2114.750 2396.000 2115.030 2400.000 ;
        RECT 2127.630 2396.000 2127.910 2400.000 ;
        RECT 2140.510 2396.000 2140.790 2400.000 ;
        RECT 2153.390 2396.000 2153.670 2400.000 ;
        RECT 2165.840 2399.450 2165.980 2414.690 ;
        RECT 2166.300 2412.630 2166.440 2588.235 ;
        RECT 2170.900 2587.730 2171.040 2598.435 ;
        RECT 2277.100 2594.210 2277.360 2594.530 ;
        RECT 2215.910 2593.675 2216.190 2594.045 ;
        RECT 2242.600 2593.870 2242.860 2594.190 ;
        RECT 2243.520 2593.870 2243.780 2594.190 ;
        RECT 2215.980 2593.510 2216.120 2593.675 ;
        RECT 2212.690 2592.995 2212.970 2593.365 ;
        RECT 2215.920 2593.190 2216.180 2593.510 ;
        RECT 2212.760 2592.830 2212.900 2592.995 ;
        RECT 2212.700 2592.510 2212.960 2592.830 ;
        RECT 2176.810 2591.635 2177.090 2592.005 ;
        RECT 2179.570 2591.635 2179.850 2592.005 ;
        RECT 2173.130 2588.235 2173.410 2588.605 ;
        RECT 2170.840 2587.410 2171.100 2587.730 ;
        RECT 2170.900 2560.190 2171.040 2587.410 ;
        RECT 2170.380 2559.870 2170.640 2560.190 ;
        RECT 2170.840 2559.870 2171.100 2560.190 ;
        RECT 2170.440 2477.765 2170.580 2559.870 ;
        RECT 2170.370 2477.395 2170.650 2477.765 ;
        RECT 2168.080 2462.970 2168.340 2463.290 ;
        RECT 2169.450 2463.115 2169.730 2463.485 ;
        RECT 2169.460 2462.970 2169.720 2463.115 ;
        RECT 2168.140 2415.205 2168.280 2462.970 ;
        RECT 2168.070 2414.835 2168.350 2415.205 ;
        RECT 2168.990 2414.835 2169.270 2415.205 ;
        RECT 2166.240 2412.310 2166.500 2412.630 ;
        RECT 2169.060 2411.950 2169.200 2414.835 ;
        RECT 2173.200 2412.290 2173.340 2588.235 ;
        RECT 2176.880 2412.970 2177.020 2591.635 ;
        RECT 2179.580 2591.490 2179.840 2591.635 ;
        RECT 2184.630 2590.955 2184.910 2591.325 ;
        RECT 2204.410 2590.955 2204.690 2591.325 ;
        RECT 2184.640 2590.810 2184.900 2590.955 ;
        RECT 2180.030 2588.235 2180.310 2588.605 ;
        RECT 2176.820 2412.650 2177.080 2412.970 ;
        RECT 2173.140 2411.970 2173.400 2412.290 ;
        RECT 2180.100 2411.950 2180.240 2588.235 ;
        RECT 2183.720 2587.750 2183.980 2588.070 ;
        RECT 2183.780 2413.650 2183.920 2587.750 ;
        RECT 2183.720 2413.330 2183.980 2413.650 ;
        RECT 2184.700 2413.310 2184.840 2590.810 ;
        RECT 2204.480 2590.790 2204.620 2590.955 ;
        RECT 2204.420 2590.470 2204.680 2590.790 ;
        RECT 2187.400 2589.790 2187.660 2590.110 ;
        RECT 2197.520 2589.790 2197.780 2590.110 ;
        RECT 2186.470 2588.915 2186.750 2589.285 ;
        RECT 2186.540 2588.070 2186.680 2588.915 ;
        RECT 2186.930 2588.235 2187.210 2588.605 ;
        RECT 2186.480 2587.750 2186.740 2588.070 ;
        RECT 2184.640 2412.990 2184.900 2413.310 ;
        RECT 2169.000 2411.630 2169.260 2411.950 ;
        RECT 2180.040 2411.630 2180.300 2411.950 ;
        RECT 2187.000 2411.610 2187.140 2588.235 ;
        RECT 2186.940 2411.290 2187.200 2411.610 ;
        RECT 2179.120 2410.610 2179.380 2410.930 ;
        RECT 2179.180 2400.000 2179.320 2410.610 ;
        RECT 2187.460 2400.130 2187.600 2589.790 ;
        RECT 2190.620 2588.090 2190.880 2588.410 ;
        RECT 2193.370 2588.235 2193.650 2588.605 ;
        RECT 2190.680 2587.925 2190.820 2588.090 ;
        RECT 2190.610 2587.555 2190.890 2587.925 ;
        RECT 2190.680 2413.990 2190.820 2587.555 ;
        RECT 2190.620 2413.670 2190.880 2413.990 ;
        RECT 2193.440 2408.550 2193.580 2588.235 ;
        RECT 2197.580 2587.925 2197.720 2589.790 ;
        RECT 2201.200 2589.450 2201.460 2589.770 ;
        RECT 2193.830 2587.555 2194.110 2587.925 ;
        RECT 2197.510 2587.555 2197.790 2587.925 ;
        RECT 2200.730 2587.555 2201.010 2587.925 ;
        RECT 2193.900 2408.890 2194.040 2587.555 ;
        RECT 2197.580 2415.010 2197.720 2587.555 ;
        RECT 2197.520 2414.690 2197.780 2415.010 ;
        RECT 2200.800 2409.230 2200.940 2587.555 ;
        RECT 2200.740 2408.910 2201.000 2409.230 ;
        RECT 2193.840 2408.570 2194.100 2408.890 ;
        RECT 2193.380 2408.230 2193.640 2408.550 ;
        RECT 2166.270 2399.450 2166.550 2400.000 ;
        RECT 2165.840 2399.310 2166.550 2399.450 ;
        RECT 2166.270 2396.000 2166.550 2399.310 ;
        RECT 2179.150 2396.000 2179.430 2400.000 ;
        RECT 2187.460 2399.990 2189.900 2400.130 ;
        RECT 2189.760 2398.770 2189.900 2399.990 ;
        RECT 2192.030 2398.770 2192.310 2400.000 ;
        RECT 2201.260 2399.450 2201.400 2589.450 ;
        RECT 2204.480 2410.930 2204.620 2590.470 ;
        RECT 2212.760 2590.450 2212.900 2592.510 ;
        RECT 2212.700 2590.130 2212.960 2590.450 ;
        RECT 2215.000 2589.110 2215.260 2589.430 ;
        RECT 2207.630 2587.555 2207.910 2587.925 ;
        RECT 2214.530 2587.555 2214.810 2587.925 ;
        RECT 2204.420 2410.610 2204.680 2410.930 ;
        RECT 2207.700 2409.570 2207.840 2587.555 ;
        RECT 2214.600 2409.910 2214.740 2587.555 ;
        RECT 2214.540 2409.590 2214.800 2409.910 ;
        RECT 2207.640 2409.250 2207.900 2409.570 ;
        RECT 2201.260 2399.310 2202.780 2399.450 ;
        RECT 2189.760 2398.630 2192.310 2398.770 ;
        RECT 2202.640 2398.770 2202.780 2399.310 ;
        RECT 2204.910 2398.770 2205.190 2400.000 ;
        RECT 2202.640 2398.630 2205.190 2398.770 ;
        RECT 2215.060 2398.770 2215.200 2589.110 ;
        RECT 2215.980 2587.730 2216.120 2593.190 ;
        RECT 2221.430 2592.995 2221.710 2593.365 ;
        RECT 2226.950 2592.995 2227.230 2593.365 ;
        RECT 2232.010 2592.995 2232.290 2593.365 ;
        RECT 2220.510 2592.315 2220.790 2592.685 ;
        RECT 2220.580 2589.770 2220.720 2592.315 ;
        RECT 2221.500 2592.150 2221.640 2592.995 ;
        RECT 2221.440 2591.830 2221.700 2592.150 ;
        RECT 2227.020 2591.810 2227.160 2592.995 ;
        RECT 2227.410 2592.315 2227.690 2592.685 ;
        RECT 2226.960 2591.490 2227.220 2591.810 ;
        RECT 2220.520 2589.450 2220.780 2589.770 ;
        RECT 2227.480 2587.730 2227.620 2592.315 ;
        RECT 2227.870 2591.635 2228.150 2592.005 ;
        RECT 2227.940 2589.430 2228.080 2591.635 ;
        RECT 2232.080 2591.470 2232.220 2592.995 ;
        RECT 2235.690 2592.315 2235.970 2592.685 ;
        RECT 2239.830 2592.315 2240.110 2592.685 ;
        RECT 2235.230 2591.635 2235.510 2592.005 ;
        RECT 2232.020 2591.150 2232.280 2591.470 ;
        RECT 2227.880 2589.110 2228.140 2589.430 ;
        RECT 2228.800 2588.770 2229.060 2589.090 ;
        RECT 2215.920 2587.410 2216.180 2587.730 ;
        RECT 2227.420 2587.410 2227.680 2587.730 ;
        RECT 2217.790 2398.770 2218.070 2400.000 ;
        RECT 2228.860 2399.450 2229.000 2588.770 ;
        RECT 2232.080 2588.070 2232.220 2591.150 ;
        RECT 2235.300 2588.750 2235.440 2591.635 ;
        RECT 2235.240 2588.430 2235.500 2588.750 ;
        RECT 2235.760 2588.410 2235.900 2592.315 ;
        RECT 2239.840 2592.170 2240.100 2592.315 ;
        RECT 2241.670 2590.955 2241.950 2591.325 ;
        RECT 2241.740 2588.410 2241.880 2590.955 ;
        RECT 2235.700 2588.090 2235.960 2588.410 ;
        RECT 2241.680 2588.090 2241.940 2588.410 ;
        RECT 2232.020 2587.750 2232.280 2588.070 ;
        RECT 2230.670 2399.450 2230.950 2400.000 ;
        RECT 2228.860 2399.310 2230.950 2399.450 ;
        RECT 2242.660 2399.450 2242.800 2593.870 ;
        RECT 2243.580 2592.685 2243.720 2593.870 ;
        RECT 2249.500 2593.530 2249.760 2593.850 ;
        RECT 2256.390 2593.675 2256.670 2594.045 ;
        RECT 2262.830 2593.675 2263.110 2594.045 ;
        RECT 2256.400 2593.530 2256.660 2593.675 ;
        RECT 2243.510 2592.315 2243.790 2592.685 ;
        RECT 2243.580 2590.110 2243.720 2592.315 ;
        RECT 2243.520 2589.790 2243.780 2590.110 ;
        RECT 2249.030 2587.555 2249.310 2587.925 ;
        RECT 2249.100 2410.250 2249.240 2587.555 ;
        RECT 2249.040 2409.930 2249.300 2410.250 ;
        RECT 2249.560 2400.130 2249.700 2593.530 ;
        RECT 2256.460 2592.830 2256.600 2593.530 ;
        RECT 2262.900 2593.510 2263.040 2593.675 ;
        RECT 2262.840 2593.190 2263.100 2593.510 ;
        RECT 2263.300 2592.850 2263.560 2593.170 ;
        RECT 2256.400 2592.510 2256.660 2592.830 ;
        RECT 2250.870 2591.635 2251.150 2592.005 ;
        RECT 2250.940 2591.130 2251.080 2591.635 ;
        RECT 2250.880 2590.810 2251.140 2591.130 ;
        RECT 2255.930 2587.555 2256.210 2587.925 ;
        RECT 2262.830 2587.555 2263.110 2587.925 ;
        RECT 2256.000 2410.590 2256.140 2587.555 ;
        RECT 2262.900 2410.930 2263.040 2587.555 ;
        RECT 2262.840 2410.610 2263.100 2410.930 ;
        RECT 2255.940 2410.270 2256.200 2410.590 ;
        RECT 2263.360 2400.130 2263.500 2592.850 ;
        RECT 2268.810 2592.315 2269.090 2592.685 ;
        RECT 2276.630 2592.315 2276.910 2592.685 ;
        RECT 2268.880 2592.150 2269.020 2592.315 ;
        RECT 2268.820 2591.830 2269.080 2592.150 ;
        RECT 2276.700 2591.810 2276.840 2592.315 ;
        RECT 2276.640 2591.490 2276.900 2591.810 ;
        RECT 2269.270 2588.235 2269.550 2588.605 ;
        RECT 2269.340 2411.270 2269.480 2588.235 ;
        RECT 2269.730 2587.555 2270.010 2587.925 ;
        RECT 2276.630 2587.555 2276.910 2587.925 ;
        RECT 2269.800 2414.670 2269.940 2587.555 ;
        RECT 2276.700 2415.010 2276.840 2587.555 ;
        RECT 2276.640 2414.690 2276.900 2415.010 ;
        RECT 2269.740 2414.350 2270.000 2414.670 ;
        RECT 2269.280 2410.950 2269.540 2411.270 ;
        RECT 2277.160 2400.130 2277.300 2594.210 ;
        RECT 2291.820 2594.045 2292.080 2594.190 ;
        RECT 2291.810 2593.675 2292.090 2594.045 ;
        RECT 2297.790 2593.675 2298.070 2594.045 ;
        RECT 2332.290 2593.675 2332.570 2594.045 ;
        RECT 2285.440 2593.510 2285.580 2593.665 ;
        RECT 2285.380 2593.365 2285.640 2593.510 ;
        RECT 2285.370 2592.995 2285.650 2593.365 ;
        RECT 2280.310 2592.315 2280.590 2592.685 ;
        RECT 2285.440 2592.490 2285.580 2592.995 ;
        RECT 2291.880 2592.490 2292.020 2593.675 ;
        RECT 2297.800 2593.530 2298.060 2593.675 ;
        RECT 2332.360 2593.510 2332.500 2593.675 ;
        RECT 2305.150 2592.995 2305.430 2593.365 ;
        RECT 2332.300 2593.190 2332.560 2593.510 ;
        RECT 2305.220 2592.830 2305.360 2592.995 ;
        RECT 2305.160 2592.510 2305.420 2592.830 ;
        RECT 2280.380 2591.470 2280.520 2592.315 ;
        RECT 2285.380 2592.170 2285.640 2592.490 ;
        RECT 2291.820 2592.170 2292.080 2592.490 ;
        RECT 2311.590 2592.315 2311.870 2592.685 ;
        RECT 2318.490 2592.315 2318.770 2592.685 ;
        RECT 2332.290 2592.315 2332.570 2592.685 ;
        RECT 2311.660 2592.150 2311.800 2592.315 ;
        RECT 2297.790 2591.635 2298.070 2592.005 ;
        RECT 2311.600 2591.830 2311.860 2592.150 ;
        RECT 2318.560 2591.810 2318.700 2592.315 ;
        RECT 2332.300 2592.170 2332.560 2592.315 ;
        RECT 2280.320 2591.150 2280.580 2591.470 ;
        RECT 2297.860 2591.130 2298.000 2591.635 ;
        RECT 2318.500 2591.490 2318.760 2591.810 ;
        RECT 2325.390 2591.635 2325.670 2592.005 ;
        RECT 2325.460 2591.470 2325.600 2591.635 ;
        RECT 2325.400 2591.150 2325.660 2591.470 ;
        RECT 2297.800 2590.810 2298.060 2591.130 ;
        RECT 2339.190 2590.955 2339.470 2591.325 ;
        RECT 2339.200 2590.810 2339.460 2590.955 ;
        RECT 2349.320 2589.450 2349.580 2589.770 ;
        RECT 2304.230 2588.235 2304.510 2588.605 ;
        RECT 2345.170 2588.235 2345.450 2588.605 ;
        RECT 2283.530 2587.555 2283.810 2587.925 ;
        RECT 2290.430 2587.555 2290.710 2587.925 ;
        RECT 2297.330 2587.555 2297.610 2587.925 ;
        RECT 2303.770 2587.555 2304.050 2587.925 ;
        RECT 2283.600 2414.330 2283.740 2587.555 ;
        RECT 2283.540 2414.010 2283.800 2414.330 ;
        RECT 2290.500 2413.990 2290.640 2587.555 ;
        RECT 2290.440 2413.670 2290.700 2413.990 ;
        RECT 2297.400 2413.650 2297.540 2587.555 ;
        RECT 2297.340 2413.330 2297.600 2413.650 ;
        RECT 2303.840 2412.970 2303.980 2587.555 ;
        RECT 2304.300 2413.310 2304.440 2588.235 ;
        RECT 2311.130 2587.555 2311.410 2587.925 ;
        RECT 2318.030 2587.555 2318.310 2587.925 ;
        RECT 2324.930 2587.555 2325.210 2587.925 ;
        RECT 2331.830 2587.555 2332.110 2587.925 ;
        RECT 2338.730 2587.555 2339.010 2587.925 ;
        RECT 2304.240 2412.990 2304.500 2413.310 ;
        RECT 2303.780 2412.650 2304.040 2412.970 ;
        RECT 2294.580 2412.310 2294.840 2412.630 ;
        RECT 2243.090 2399.450 2243.370 2400.000 ;
        RECT 2249.560 2399.990 2253.380 2400.130 ;
        RECT 2242.660 2399.310 2243.370 2399.450 ;
        RECT 2215.060 2398.630 2218.070 2398.770 ;
        RECT 2192.030 2396.000 2192.310 2398.630 ;
        RECT 2204.910 2396.000 2205.190 2398.630 ;
        RECT 2217.790 2396.000 2218.070 2398.630 ;
        RECT 2230.670 2396.000 2230.950 2399.310 ;
        RECT 2243.090 2396.000 2243.370 2399.310 ;
        RECT 2253.240 2398.770 2253.380 2399.990 ;
        RECT 2255.970 2398.770 2256.250 2400.000 ;
        RECT 2263.360 2399.990 2266.260 2400.130 ;
        RECT 2253.240 2398.630 2256.250 2398.770 ;
        RECT 2266.120 2398.770 2266.260 2399.990 ;
        RECT 2268.850 2398.770 2269.130 2400.000 ;
        RECT 2277.160 2399.990 2279.140 2400.130 ;
        RECT 2294.640 2400.000 2294.780 2412.310 ;
        RECT 2311.200 2412.290 2311.340 2587.555 ;
        RECT 2318.100 2412.630 2318.240 2587.555 ;
        RECT 2318.040 2412.310 2318.300 2412.630 ;
        RECT 2307.460 2411.970 2307.720 2412.290 ;
        RECT 2311.140 2411.970 2311.400 2412.290 ;
        RECT 2307.520 2400.000 2307.660 2411.970 ;
        RECT 2325.000 2411.950 2325.140 2587.555 ;
        RECT 2331.900 2412.485 2332.040 2587.555 ;
        RECT 2331.830 2412.115 2332.110 2412.485 ;
        RECT 2320.340 2411.630 2320.600 2411.950 ;
        RECT 2324.940 2411.630 2325.200 2411.950 ;
        RECT 2320.400 2400.000 2320.540 2411.630 ;
        RECT 2338.800 2411.610 2338.940 2587.555 ;
        RECT 2345.240 2411.805 2345.380 2588.235 ;
        RECT 2345.630 2587.555 2345.910 2587.925 ;
        RECT 2333.220 2411.290 2333.480 2411.610 ;
        RECT 2338.740 2411.290 2339.000 2411.610 ;
        RECT 2345.170 2411.435 2345.450 2411.805 ;
        RECT 2333.280 2400.000 2333.420 2411.290 ;
        RECT 2345.700 2411.125 2345.840 2587.555 ;
        RECT 2345.630 2410.755 2345.910 2411.125 ;
        RECT 2349.380 2408.550 2349.520 2589.450 ;
        RECT 2383.820 2589.110 2384.080 2589.430 ;
        RECT 2370.020 2588.430 2370.280 2588.750 ;
        RECT 2356.220 2588.090 2356.480 2588.410 ;
        RECT 2356.280 2409.085 2356.420 2588.090 ;
        RECT 2356.210 2408.715 2356.490 2409.085 ;
        RECT 2370.080 2408.890 2370.220 2588.430 ;
        RECT 2383.880 2409.230 2384.020 2589.110 ;
        RECT 2397.620 2587.410 2397.880 2587.730 ;
        RECT 2397.680 2409.910 2397.820 2587.410 ;
        RECT 2538.840 2414.690 2539.100 2415.010 ;
        RECT 2525.960 2414.350 2526.220 2414.670 ;
        RECT 2513.080 2410.950 2513.340 2411.270 ;
        RECT 2500.200 2410.610 2500.460 2410.930 ;
        RECT 2487.320 2410.270 2487.580 2410.590 ;
        RECT 2474.440 2409.930 2474.700 2410.250 ;
        RECT 2397.160 2409.590 2397.420 2409.910 ;
        RECT 2397.620 2409.590 2397.880 2409.910 ;
        RECT 2422.920 2409.590 2423.180 2409.910 ;
        RECT 2384.740 2409.250 2385.000 2409.570 ;
        RECT 2371.860 2408.910 2372.120 2409.230 ;
        RECT 2383.820 2408.910 2384.080 2409.230 ;
        RECT 2358.980 2408.570 2359.240 2408.890 ;
        RECT 2370.020 2408.570 2370.280 2408.890 ;
        RECT 2346.100 2408.230 2346.360 2408.550 ;
        RECT 2349.320 2408.230 2349.580 2408.550 ;
        RECT 2346.160 2400.000 2346.300 2408.230 ;
        RECT 2359.040 2400.000 2359.180 2408.570 ;
        RECT 2371.920 2400.000 2372.060 2408.910 ;
        RECT 2384.800 2400.000 2384.940 2409.250 ;
        RECT 2386.110 2408.715 2386.390 2409.085 ;
        RECT 2386.120 2408.570 2386.380 2408.715 ;
        RECT 2385.660 2408.290 2385.920 2408.550 ;
        RECT 2386.580 2408.290 2386.840 2408.550 ;
        RECT 2385.660 2408.230 2386.840 2408.290 ;
        RECT 2385.720 2408.150 2386.780 2408.230 ;
        RECT 2397.220 2400.000 2397.360 2409.590 ;
        RECT 2410.040 2408.230 2410.300 2408.550 ;
        RECT 2410.100 2400.000 2410.240 2408.230 ;
        RECT 2422.980 2400.000 2423.120 2409.590 ;
        RECT 2435.800 2409.250 2436.060 2409.570 ;
        RECT 2435.860 2400.000 2436.000 2409.250 ;
        RECT 2448.680 2408.910 2448.940 2409.230 ;
        RECT 2448.740 2400.000 2448.880 2408.910 ;
        RECT 2461.560 2408.570 2461.820 2408.890 ;
        RECT 2461.620 2400.000 2461.760 2408.570 ;
        RECT 2474.500 2400.000 2474.640 2409.930 ;
        RECT 2487.380 2400.000 2487.520 2410.270 ;
        RECT 2500.260 2400.000 2500.400 2410.610 ;
        RECT 2513.140 2400.000 2513.280 2410.950 ;
        RECT 2526.020 2400.000 2526.160 2414.350 ;
        RECT 2538.900 2400.000 2539.040 2414.690 ;
        RECT 2551.260 2414.010 2551.520 2414.330 ;
        RECT 2551.320 2400.000 2551.460 2414.010 ;
        RECT 2564.140 2413.670 2564.400 2413.990 ;
        RECT 2564.200 2400.000 2564.340 2413.670 ;
        RECT 2577.020 2413.330 2577.280 2413.650 ;
        RECT 2577.080 2400.000 2577.220 2413.330 ;
        RECT 2589.900 2412.990 2590.160 2413.310 ;
        RECT 2589.960 2400.000 2590.100 2412.990 ;
        RECT 2602.780 2412.650 2603.040 2412.970 ;
        RECT 2602.840 2400.000 2602.980 2412.650 ;
        RECT 2628.540 2412.310 2628.800 2412.630 ;
        RECT 2615.660 2411.970 2615.920 2412.290 ;
        RECT 2615.720 2400.000 2615.860 2411.970 ;
        RECT 2628.600 2400.000 2628.740 2412.310 ;
        RECT 2654.290 2412.115 2654.570 2412.485 ;
        RECT 2641.420 2411.630 2641.680 2411.950 ;
        RECT 2641.480 2400.000 2641.620 2411.630 ;
        RECT 2654.360 2400.000 2654.500 2412.115 ;
        RECT 2667.180 2411.290 2667.440 2411.610 ;
        RECT 2680.050 2411.435 2680.330 2411.805 ;
        RECT 2667.240 2400.000 2667.380 2411.290 ;
        RECT 2680.120 2400.000 2680.260 2411.435 ;
        RECT 2692.930 2410.755 2693.210 2411.125 ;
        RECT 2693.000 2400.000 2693.140 2410.755 ;
        RECT 2266.120 2398.630 2269.130 2398.770 ;
        RECT 2279.000 2398.770 2279.140 2399.990 ;
        RECT 2281.730 2398.770 2282.010 2400.000 ;
        RECT 2279.000 2398.630 2282.010 2398.770 ;
        RECT 2255.970 2396.000 2256.250 2398.630 ;
        RECT 2268.850 2396.000 2269.130 2398.630 ;
        RECT 2281.730 2396.000 2282.010 2398.630 ;
        RECT 2294.610 2396.000 2294.890 2400.000 ;
        RECT 2307.490 2396.000 2307.770 2400.000 ;
        RECT 2320.370 2396.000 2320.650 2400.000 ;
        RECT 2333.250 2396.000 2333.530 2400.000 ;
        RECT 2346.130 2396.000 2346.410 2400.000 ;
        RECT 2359.010 2396.000 2359.290 2400.000 ;
        RECT 2371.890 2396.000 2372.170 2400.000 ;
        RECT 2384.770 2396.000 2385.050 2400.000 ;
        RECT 2397.190 2396.000 2397.470 2400.000 ;
        RECT 2410.070 2396.000 2410.350 2400.000 ;
        RECT 2422.950 2396.000 2423.230 2400.000 ;
        RECT 2435.830 2396.000 2436.110 2400.000 ;
        RECT 2448.710 2396.000 2448.990 2400.000 ;
        RECT 2461.590 2396.000 2461.870 2400.000 ;
        RECT 2474.470 2396.000 2474.750 2400.000 ;
        RECT 2487.350 2396.000 2487.630 2400.000 ;
        RECT 2500.230 2396.000 2500.510 2400.000 ;
        RECT 2513.110 2396.000 2513.390 2400.000 ;
        RECT 2525.990 2396.000 2526.270 2400.000 ;
        RECT 2538.870 2396.000 2539.150 2400.000 ;
        RECT 2551.290 2396.000 2551.570 2400.000 ;
        RECT 2564.170 2396.000 2564.450 2400.000 ;
        RECT 2577.050 2396.000 2577.330 2400.000 ;
        RECT 2589.930 2396.000 2590.210 2400.000 ;
        RECT 2602.810 2396.000 2603.090 2400.000 ;
        RECT 2615.690 2396.000 2615.970 2400.000 ;
        RECT 2628.570 2396.000 2628.850 2400.000 ;
        RECT 2641.450 2396.000 2641.730 2400.000 ;
        RECT 2654.330 2396.000 2654.610 2400.000 ;
        RECT 2667.210 2396.000 2667.490 2400.000 ;
        RECT 2680.090 2396.000 2680.370 2400.000 ;
        RECT 2692.970 2396.000 2693.250 2400.000 ;
      LAYER met2 ;
        RECT 1306.630 2395.720 1318.210 2396.000 ;
        RECT 1319.050 2395.720 1331.090 2396.000 ;
        RECT 1331.930 2395.720 1343.970 2396.000 ;
        RECT 1344.810 2395.720 1356.850 2396.000 ;
        RECT 1357.690 2395.720 1369.730 2396.000 ;
        RECT 1370.570 2395.720 1382.610 2396.000 ;
        RECT 1383.450 2395.720 1395.490 2396.000 ;
        RECT 1396.330 2395.720 1408.370 2396.000 ;
        RECT 1409.210 2395.720 1421.250 2396.000 ;
        RECT 1422.090 2395.720 1434.130 2396.000 ;
        RECT 1434.970 2395.720 1447.010 2396.000 ;
        RECT 1447.850 2395.720 1459.890 2396.000 ;
        RECT 1460.730 2395.720 1472.310 2396.000 ;
        RECT 1473.150 2395.720 1485.190 2396.000 ;
        RECT 1486.030 2395.720 1498.070 2396.000 ;
        RECT 1498.910 2395.720 1510.950 2396.000 ;
        RECT 1511.790 2395.720 1523.830 2396.000 ;
        RECT 1524.670 2395.720 1536.710 2396.000 ;
        RECT 1537.550 2395.720 1549.590 2396.000 ;
        RECT 1550.430 2395.720 1562.470 2396.000 ;
        RECT 1563.310 2395.720 1575.350 2396.000 ;
        RECT 1576.190 2395.720 1588.230 2396.000 ;
        RECT 1589.070 2395.720 1601.110 2396.000 ;
        RECT 1601.950 2395.720 1613.990 2396.000 ;
        RECT 1614.830 2395.720 1626.410 2396.000 ;
        RECT 1627.250 2395.720 1639.290 2396.000 ;
        RECT 1640.130 2395.720 1652.170 2396.000 ;
        RECT 1653.010 2395.720 1665.050 2396.000 ;
        RECT 1665.890 2395.720 1677.930 2396.000 ;
        RECT 1678.770 2395.720 1690.810 2396.000 ;
        RECT 1691.650 2395.720 1703.690 2396.000 ;
        RECT 1704.530 2395.720 1716.570 2396.000 ;
        RECT 1717.410 2395.720 1729.450 2396.000 ;
        RECT 1730.290 2395.720 1742.330 2396.000 ;
        RECT 1743.170 2395.720 1755.210 2396.000 ;
        RECT 1756.050 2395.720 1768.090 2396.000 ;
        RECT 1768.930 2395.720 1780.510 2396.000 ;
        RECT 1781.350 2395.720 1793.390 2396.000 ;
        RECT 1794.230 2395.720 1806.270 2396.000 ;
        RECT 1807.110 2395.720 1819.150 2396.000 ;
        RECT 1819.990 2395.720 1832.030 2396.000 ;
        RECT 1832.870 2395.720 1844.910 2396.000 ;
        RECT 1845.750 2395.720 1857.790 2396.000 ;
        RECT 1858.630 2395.720 1870.670 2396.000 ;
        RECT 1871.510 2395.720 1883.550 2396.000 ;
        RECT 1884.390 2395.720 1896.430 2396.000 ;
        RECT 1897.270 2395.720 1909.310 2396.000 ;
        RECT 1910.150 2395.720 1922.190 2396.000 ;
        RECT 1923.030 2395.720 1934.610 2396.000 ;
        RECT 1935.450 2395.720 1947.490 2396.000 ;
        RECT 1948.330 2395.720 1960.370 2396.000 ;
        RECT 1961.210 2395.720 1973.250 2396.000 ;
        RECT 1974.090 2395.720 1986.130 2396.000 ;
        RECT 1986.970 2395.720 1999.010 2396.000 ;
        RECT 1999.850 2395.720 2011.890 2396.000 ;
        RECT 2012.730 2395.720 2024.770 2396.000 ;
        RECT 2025.610 2395.720 2037.650 2396.000 ;
        RECT 2038.490 2395.720 2050.530 2396.000 ;
        RECT 2051.370 2395.720 2063.410 2396.000 ;
        RECT 2064.250 2395.720 2076.290 2396.000 ;
        RECT 2077.130 2395.720 2088.710 2396.000 ;
        RECT 2089.550 2395.720 2101.590 2396.000 ;
        RECT 2102.430 2395.720 2114.470 2396.000 ;
        RECT 2115.310 2395.720 2127.350 2396.000 ;
        RECT 2128.190 2395.720 2140.230 2396.000 ;
        RECT 2141.070 2395.720 2153.110 2396.000 ;
        RECT 2153.950 2395.720 2165.990 2396.000 ;
        RECT 2166.830 2395.720 2178.870 2396.000 ;
        RECT 2179.710 2395.720 2191.750 2396.000 ;
        RECT 2192.590 2395.720 2204.630 2396.000 ;
        RECT 2205.470 2395.720 2217.510 2396.000 ;
        RECT 2218.350 2395.720 2230.390 2396.000 ;
        RECT 2231.230 2395.720 2242.810 2396.000 ;
        RECT 2243.650 2395.720 2255.690 2396.000 ;
        RECT 2256.530 2395.720 2268.570 2396.000 ;
        RECT 2269.410 2395.720 2281.450 2396.000 ;
        RECT 2282.290 2395.720 2294.330 2396.000 ;
        RECT 2295.170 2395.720 2307.210 2396.000 ;
        RECT 2308.050 2395.720 2320.090 2396.000 ;
        RECT 2320.930 2395.720 2332.970 2396.000 ;
        RECT 2333.810 2395.720 2345.850 2396.000 ;
        RECT 2346.690 2395.720 2358.730 2396.000 ;
        RECT 2359.570 2395.720 2371.610 2396.000 ;
        RECT 2372.450 2395.720 2384.490 2396.000 ;
        RECT 2385.330 2395.720 2396.910 2396.000 ;
        RECT 2397.750 2395.720 2409.790 2396.000 ;
        RECT 2410.630 2395.720 2422.670 2396.000 ;
        RECT 2423.510 2395.720 2435.550 2396.000 ;
        RECT 2436.390 2395.720 2448.430 2396.000 ;
        RECT 2449.270 2395.720 2461.310 2396.000 ;
        RECT 2462.150 2395.720 2474.190 2396.000 ;
        RECT 2475.030 2395.720 2487.070 2396.000 ;
        RECT 2487.910 2395.720 2499.950 2396.000 ;
        RECT 2500.790 2395.720 2512.830 2396.000 ;
        RECT 2513.670 2395.720 2525.710 2396.000 ;
        RECT 2526.550 2395.720 2538.590 2396.000 ;
        RECT 2539.430 2395.720 2551.010 2396.000 ;
        RECT 2551.850 2395.720 2563.890 2396.000 ;
        RECT 2564.730 2395.720 2576.770 2396.000 ;
        RECT 2577.610 2395.720 2589.650 2396.000 ;
        RECT 2590.490 2395.720 2602.530 2396.000 ;
        RECT 2603.370 2395.720 2615.410 2396.000 ;
        RECT 2616.250 2395.720 2628.290 2396.000 ;
        RECT 2629.130 2395.720 2641.170 2396.000 ;
        RECT 2642.010 2395.720 2654.050 2396.000 ;
        RECT 2654.890 2395.720 2666.930 2396.000 ;
        RECT 2667.770 2395.720 2679.810 2396.000 ;
        RECT 2680.650 2395.720 2692.690 2396.000 ;
        RECT 2693.530 2395.720 2695.550 2396.000 ;
        RECT 1306.080 1204.280 2695.550 2395.720 ;
        RECT 1306.630 1204.000 1318.210 1204.280 ;
        RECT 1319.050 1204.000 1331.090 1204.280 ;
        RECT 1331.930 1204.000 1343.970 1204.280 ;
        RECT 1344.810 1204.000 1356.850 1204.280 ;
        RECT 1357.690 1204.000 1369.730 1204.280 ;
        RECT 1370.570 1204.000 1382.610 1204.280 ;
        RECT 1383.450 1204.000 1395.490 1204.280 ;
        RECT 1396.330 1204.000 1408.370 1204.280 ;
        RECT 1409.210 1204.000 1421.250 1204.280 ;
        RECT 1422.090 1204.000 1434.130 1204.280 ;
        RECT 1434.970 1204.000 1447.010 1204.280 ;
        RECT 1447.850 1204.000 1459.890 1204.280 ;
        RECT 1460.730 1204.000 1472.310 1204.280 ;
        RECT 1473.150 1204.000 1485.190 1204.280 ;
        RECT 1486.030 1204.000 1498.070 1204.280 ;
        RECT 1498.910 1204.000 1510.950 1204.280 ;
        RECT 1511.790 1204.000 1523.830 1204.280 ;
        RECT 1524.670 1204.000 1536.710 1204.280 ;
        RECT 1537.550 1204.000 1549.590 1204.280 ;
        RECT 1550.430 1204.000 1562.470 1204.280 ;
        RECT 1563.310 1204.000 1575.350 1204.280 ;
        RECT 1576.190 1204.000 1588.230 1204.280 ;
        RECT 1589.070 1204.000 1601.110 1204.280 ;
        RECT 1601.950 1204.000 1613.990 1204.280 ;
        RECT 1614.830 1204.000 1626.410 1204.280 ;
        RECT 1627.250 1204.000 1639.290 1204.280 ;
        RECT 1640.130 1204.000 1652.170 1204.280 ;
        RECT 1653.010 1204.000 1665.050 1204.280 ;
        RECT 1665.890 1204.000 1677.930 1204.280 ;
        RECT 1678.770 1204.000 1690.810 1204.280 ;
        RECT 1691.650 1204.000 1703.690 1204.280 ;
        RECT 1704.530 1204.000 1716.570 1204.280 ;
        RECT 1717.410 1204.000 1729.450 1204.280 ;
        RECT 1730.290 1204.000 1742.330 1204.280 ;
        RECT 1743.170 1204.000 1755.210 1204.280 ;
        RECT 1756.050 1204.000 1768.090 1204.280 ;
        RECT 1768.930 1204.000 1780.510 1204.280 ;
        RECT 1781.350 1204.000 1793.390 1204.280 ;
        RECT 1794.230 1204.000 1806.270 1204.280 ;
        RECT 1807.110 1204.000 1819.150 1204.280 ;
        RECT 1819.990 1204.000 1832.030 1204.280 ;
        RECT 1832.870 1204.000 1844.910 1204.280 ;
        RECT 1845.750 1204.000 1857.790 1204.280 ;
        RECT 1858.630 1204.000 1870.670 1204.280 ;
        RECT 1871.510 1204.000 1883.550 1204.280 ;
        RECT 1884.390 1204.000 1896.430 1204.280 ;
        RECT 1897.270 1204.000 1909.310 1204.280 ;
        RECT 1910.150 1204.000 1922.190 1204.280 ;
        RECT 1923.030 1204.000 1934.610 1204.280 ;
        RECT 1935.450 1204.000 1947.490 1204.280 ;
        RECT 1948.330 1204.000 1960.370 1204.280 ;
        RECT 1961.210 1204.000 1973.250 1204.280 ;
        RECT 1974.090 1204.000 1986.130 1204.280 ;
        RECT 1986.970 1204.000 1999.010 1204.280 ;
        RECT 1999.850 1204.000 2011.890 1204.280 ;
        RECT 2012.730 1204.000 2024.770 1204.280 ;
        RECT 2025.610 1204.000 2037.650 1204.280 ;
        RECT 2038.490 1204.000 2050.530 1204.280 ;
        RECT 2051.370 1204.000 2063.410 1204.280 ;
        RECT 2064.250 1204.000 2076.290 1204.280 ;
        RECT 2077.130 1204.000 2088.710 1204.280 ;
        RECT 2089.550 1204.000 2101.590 1204.280 ;
        RECT 2102.430 1204.000 2114.470 1204.280 ;
        RECT 2115.310 1204.000 2127.350 1204.280 ;
        RECT 2128.190 1204.000 2140.230 1204.280 ;
        RECT 2141.070 1204.000 2153.110 1204.280 ;
        RECT 2153.950 1204.000 2165.990 1204.280 ;
        RECT 2166.830 1204.000 2178.870 1204.280 ;
        RECT 2179.710 1204.000 2191.750 1204.280 ;
        RECT 2192.590 1204.000 2204.630 1204.280 ;
        RECT 2205.470 1204.000 2217.510 1204.280 ;
        RECT 2218.350 1204.000 2230.390 1204.280 ;
        RECT 2231.230 1204.000 2242.810 1204.280 ;
        RECT 2243.650 1204.000 2255.690 1204.280 ;
        RECT 2256.530 1204.000 2268.570 1204.280 ;
        RECT 2269.410 1204.000 2281.450 1204.280 ;
        RECT 2282.290 1204.000 2294.330 1204.280 ;
        RECT 2295.170 1204.000 2307.210 1204.280 ;
        RECT 2308.050 1204.000 2320.090 1204.280 ;
        RECT 2320.930 1204.000 2332.970 1204.280 ;
        RECT 2333.810 1204.000 2345.850 1204.280 ;
        RECT 2346.690 1204.000 2358.730 1204.280 ;
        RECT 2359.570 1204.000 2371.610 1204.280 ;
        RECT 2372.450 1204.000 2384.490 1204.280 ;
        RECT 2385.330 1204.000 2396.910 1204.280 ;
        RECT 2397.750 1204.000 2409.790 1204.280 ;
        RECT 2410.630 1204.000 2422.670 1204.280 ;
        RECT 2423.510 1204.000 2435.550 1204.280 ;
        RECT 2436.390 1204.000 2448.430 1204.280 ;
        RECT 2449.270 1204.000 2461.310 1204.280 ;
        RECT 2462.150 1204.000 2474.190 1204.280 ;
        RECT 2475.030 1204.000 2487.070 1204.280 ;
        RECT 2487.910 1204.000 2499.950 1204.280 ;
        RECT 2500.790 1204.000 2512.830 1204.280 ;
        RECT 2513.670 1204.000 2525.710 1204.280 ;
        RECT 2526.550 1204.000 2538.590 1204.280 ;
        RECT 2539.430 1204.000 2551.010 1204.280 ;
        RECT 2551.850 1204.000 2563.890 1204.280 ;
        RECT 2564.730 1204.000 2576.770 1204.280 ;
        RECT 2577.610 1204.000 2589.650 1204.280 ;
        RECT 2590.490 1204.000 2602.530 1204.280 ;
        RECT 2603.370 1204.000 2615.410 1204.280 ;
        RECT 2616.250 1204.000 2628.290 1204.280 ;
        RECT 2629.130 1204.000 2641.170 1204.280 ;
        RECT 2642.010 1204.000 2654.050 1204.280 ;
        RECT 2654.890 1204.000 2666.930 1204.280 ;
        RECT 2667.770 1204.000 2679.810 1204.280 ;
        RECT 2680.650 1204.000 2692.690 1204.280 ;
        RECT 2693.530 1204.000 2695.550 1204.280 ;
      LAYER met2 ;
        RECT 1318.490 1200.000 1318.770 1204.000 ;
        RECT 1331.370 1200.000 1331.650 1204.000 ;
        RECT 1344.250 1200.610 1344.530 1204.000 ;
        RECT 1357.130 1200.610 1357.410 1204.000 ;
        RECT 1370.010 1200.610 1370.290 1204.000 ;
        RECT 1344.250 1200.470 1345.340 1200.610 ;
        RECT 1344.250 1200.000 1344.530 1200.470 ;
        RECT 1318.520 1193.050 1318.660 1200.000 ;
        RECT 1318.460 1192.730 1318.720 1193.050 ;
        RECT 1331.400 1190.330 1331.540 1200.000 ;
        RECT 1331.340 1190.010 1331.600 1190.330 ;
        RECT 1345.200 1019.165 1345.340 1200.470 ;
        RECT 1357.130 1200.470 1359.140 1200.610 ;
        RECT 1357.130 1200.000 1357.410 1200.470 ;
        RECT 1359.000 1019.845 1359.140 1200.470 ;
        RECT 1370.010 1200.470 1372.940 1200.610 ;
        RECT 1370.010 1200.000 1370.290 1200.470 ;
        RECT 1372.800 1020.525 1372.940 1200.470 ;
        RECT 1382.890 1200.000 1383.170 1204.000 ;
        RECT 1395.770 1200.000 1396.050 1204.000 ;
        RECT 1408.650 1200.000 1408.930 1204.000 ;
        RECT 1421.530 1200.000 1421.810 1204.000 ;
        RECT 1434.410 1200.000 1434.690 1204.000 ;
        RECT 1447.290 1200.000 1447.570 1204.000 ;
        RECT 1460.170 1200.000 1460.450 1204.000 ;
        RECT 1472.590 1200.000 1472.870 1204.000 ;
        RECT 1485.470 1200.000 1485.750 1204.000 ;
        RECT 1498.350 1200.000 1498.630 1204.000 ;
        RECT 1511.230 1200.000 1511.510 1204.000 ;
        RECT 1524.110 1200.610 1524.390 1204.000 ;
        RECT 1536.990 1200.610 1537.270 1204.000 ;
        RECT 1549.870 1200.610 1550.150 1204.000 ;
        RECT 1562.750 1200.610 1563.030 1204.000 ;
        RECT 1524.110 1200.470 1524.740 1200.610 ;
        RECT 1524.110 1200.000 1524.390 1200.470 ;
        RECT 1382.920 1187.270 1383.060 1200.000 ;
        RECT 1395.800 1187.270 1395.940 1200.000 ;
        RECT 1408.680 1187.270 1408.820 1200.000 ;
        RECT 1421.560 1191.350 1421.700 1200.000 ;
        RECT 1421.500 1191.030 1421.760 1191.350 ;
        RECT 1434.440 1191.010 1434.580 1200.000 ;
        RECT 1447.320 1191.690 1447.460 1200.000 ;
        RECT 1447.260 1191.370 1447.520 1191.690 ;
        RECT 1434.380 1190.690 1434.640 1191.010 ;
        RECT 1460.200 1190.670 1460.340 1200.000 ;
        RECT 1472.620 1192.030 1472.760 1200.000 ;
        RECT 1485.500 1192.370 1485.640 1200.000 ;
        RECT 1489.120 1192.730 1489.380 1193.050 ;
        RECT 1485.440 1192.050 1485.700 1192.370 ;
        RECT 1472.560 1191.710 1472.820 1192.030 ;
        RECT 1460.140 1190.350 1460.400 1190.670 ;
        RECT 1382.860 1186.950 1383.120 1187.270 ;
        RECT 1386.540 1186.950 1386.800 1187.270 ;
        RECT 1395.740 1186.950 1396.000 1187.270 ;
        RECT 1400.340 1186.950 1400.600 1187.270 ;
        RECT 1408.620 1186.950 1408.880 1187.270 ;
        RECT 1414.140 1186.950 1414.400 1187.270 ;
        RECT 1386.600 1021.205 1386.740 1186.950 ;
        RECT 1386.530 1020.835 1386.810 1021.205 ;
        RECT 1372.730 1020.155 1373.010 1020.525 ;
        RECT 1358.930 1019.475 1359.210 1019.845 ;
        RECT 1345.130 1018.795 1345.410 1019.165 ;
        RECT 1400.400 1014.890 1400.540 1186.950 ;
        RECT 1414.200 1021.010 1414.340 1186.950 ;
        RECT 1414.140 1020.690 1414.400 1021.010 ;
        RECT 1400.340 1014.570 1400.600 1014.890 ;
        RECT 1489.180 558.805 1489.320 1192.730 ;
        RECT 1498.380 1187.270 1498.520 1200.000 ;
        RECT 1511.260 1187.270 1511.400 1200.000 ;
        RECT 1498.320 1186.950 1498.580 1187.270 ;
        RECT 1503.840 1186.950 1504.100 1187.270 ;
        RECT 1511.200 1186.950 1511.460 1187.270 ;
        RECT 1517.640 1186.950 1517.900 1187.270 ;
        RECT 1503.900 1020.670 1504.040 1186.950 ;
        RECT 1503.840 1020.350 1504.100 1020.670 ;
        RECT 1517.700 1020.330 1517.840 1186.950 ;
        RECT 1517.640 1020.010 1517.900 1020.330 ;
        RECT 1524.600 1019.990 1524.740 1200.470 ;
        RECT 1536.990 1200.470 1538.540 1200.610 ;
        RECT 1536.990 1200.000 1537.270 1200.470 ;
        RECT 1524.540 1019.670 1524.800 1019.990 ;
        RECT 1538.400 1019.650 1538.540 1200.470 ;
        RECT 1549.870 1200.470 1552.340 1200.610 ;
        RECT 1549.870 1200.000 1550.150 1200.470 ;
        RECT 1538.340 1019.330 1538.600 1019.650 ;
        RECT 1552.200 1019.310 1552.340 1200.470 ;
        RECT 1562.750 1200.470 1566.140 1200.610 ;
        RECT 1562.750 1200.000 1563.030 1200.470 ;
        RECT 1552.140 1018.990 1552.400 1019.310 ;
        RECT 1566.000 1018.970 1566.140 1200.470 ;
        RECT 1575.630 1200.000 1575.910 1204.000 ;
        RECT 1588.510 1200.000 1588.790 1204.000 ;
        RECT 1601.390 1200.000 1601.670 1204.000 ;
        RECT 1614.270 1200.000 1614.550 1204.000 ;
        RECT 1626.690 1200.000 1626.970 1204.000 ;
        RECT 1639.570 1200.610 1639.850 1204.000 ;
        RECT 1652.450 1200.610 1652.730 1204.000 ;
        RECT 1639.570 1200.470 1641.580 1200.610 ;
        RECT 1639.570 1200.000 1639.850 1200.470 ;
        RECT 1575.660 1187.270 1575.800 1200.000 ;
        RECT 1588.540 1187.270 1588.680 1200.000 ;
        RECT 1601.420 1187.270 1601.560 1200.000 ;
        RECT 1575.600 1186.950 1575.860 1187.270 ;
        RECT 1579.740 1186.950 1580.000 1187.270 ;
        RECT 1588.480 1186.950 1588.740 1187.270 ;
        RECT 1593.540 1186.950 1593.800 1187.270 ;
        RECT 1601.360 1186.950 1601.620 1187.270 ;
        RECT 1607.340 1186.950 1607.600 1187.270 ;
        RECT 1565.940 1018.650 1566.200 1018.970 ;
        RECT 1579.800 1014.550 1579.940 1186.950 ;
        RECT 1593.600 1018.290 1593.740 1186.950 ;
        RECT 1593.540 1017.970 1593.800 1018.290 ;
        RECT 1607.400 1017.950 1607.540 1186.950 ;
        RECT 1607.340 1017.630 1607.600 1017.950 ;
        RECT 1614.300 1017.610 1614.440 1200.000 ;
        RECT 1626.720 1193.390 1626.860 1200.000 ;
        RECT 1626.660 1193.070 1626.920 1193.390 ;
        RECT 1614.240 1017.290 1614.500 1017.610 ;
        RECT 1641.440 1016.930 1641.580 1200.470 ;
        RECT 1652.450 1200.470 1655.380 1200.610 ;
        RECT 1652.450 1200.000 1652.730 1200.470 ;
        RECT 1648.740 1192.730 1649.000 1193.050 ;
        RECT 1641.840 1192.390 1642.100 1192.710 ;
        RECT 1641.900 1018.485 1642.040 1192.390 ;
        RECT 1648.800 1018.485 1648.940 1192.730 ;
        RECT 1655.240 1021.350 1655.380 1200.470 ;
        RECT 1665.330 1200.000 1665.610 1204.000 ;
        RECT 1678.210 1200.000 1678.490 1204.000 ;
        RECT 1691.090 1200.000 1691.370 1204.000 ;
        RECT 1703.970 1200.000 1704.250 1204.000 ;
        RECT 1716.850 1200.000 1717.130 1204.000 ;
        RECT 1729.730 1200.000 1730.010 1204.000 ;
        RECT 1742.610 1200.610 1742.890 1204.000 ;
        RECT 1742.610 1200.470 1745.540 1200.610 ;
        RECT 1742.610 1200.000 1742.890 1200.470 ;
        RECT 1655.640 1193.410 1655.900 1193.730 ;
        RECT 1655.180 1021.030 1655.440 1021.350 ;
        RECT 1655.700 1018.485 1655.840 1193.410 ;
        RECT 1662.540 1187.630 1662.800 1187.950 ;
        RECT 1661.620 1018.650 1661.880 1018.970 ;
        RECT 1662.080 1018.650 1662.340 1018.970 ;
        RECT 1641.830 1018.115 1642.110 1018.485 ;
        RECT 1648.730 1018.115 1649.010 1018.485 ;
        RECT 1655.630 1018.115 1655.910 1018.485 ;
        RECT 1641.840 1017.125 1642.100 1017.270 ;
        RECT 1641.380 1016.610 1641.640 1016.930 ;
        RECT 1641.830 1016.755 1642.110 1017.125 ;
        RECT 1655.640 1016.445 1655.900 1016.590 ;
        RECT 1648.740 1015.930 1649.000 1016.250 ;
        RECT 1655.630 1016.075 1655.910 1016.445 ;
        RECT 1648.800 1015.765 1648.940 1015.930 ;
        RECT 1648.730 1015.395 1649.010 1015.765 ;
        RECT 1661.680 1015.570 1661.820 1018.650 ;
        RECT 1662.140 1017.125 1662.280 1018.650 ;
        RECT 1662.070 1016.755 1662.350 1017.125 ;
        RECT 1662.600 1016.445 1662.740 1187.630 ;
        RECT 1665.360 1187.270 1665.500 1200.000 ;
        RECT 1678.240 1187.610 1678.380 1200.000 ;
        RECT 1683.700 1193.070 1683.960 1193.390 ;
        RECT 1669.440 1187.290 1669.700 1187.610 ;
        RECT 1678.180 1187.290 1678.440 1187.610 ;
        RECT 1665.300 1186.950 1665.560 1187.270 ;
        RECT 1669.500 1017.125 1669.640 1187.290 ;
        RECT 1669.900 1186.950 1670.160 1187.270 ;
        RECT 1669.430 1016.755 1669.710 1017.125 ;
        RECT 1662.530 1016.075 1662.810 1016.445 ;
        RECT 1669.440 1016.270 1669.700 1016.590 ;
        RECT 1669.960 1016.445 1670.100 1186.950 ;
        RECT 1670.360 1021.030 1670.620 1021.350 ;
        RECT 1681.860 1021.030 1682.120 1021.350 ;
        RECT 1670.420 1018.485 1670.560 1021.030 ;
        RECT 1681.920 1018.970 1682.060 1021.030 ;
        RECT 1681.860 1018.650 1682.120 1018.970 ;
        RECT 1682.320 1018.650 1682.580 1018.970 ;
        RECT 1670.350 1018.115 1670.630 1018.485 ;
        RECT 1675.870 1017.435 1676.150 1017.805 ;
        RECT 1669.500 1015.765 1669.640 1016.270 ;
        RECT 1669.890 1016.075 1670.170 1016.445 ;
        RECT 1675.940 1016.250 1676.080 1017.435 ;
        RECT 1676.800 1016.610 1677.060 1016.930 ;
        RECT 1676.860 1016.445 1677.000 1016.610 ;
        RECT 1675.880 1015.930 1676.140 1016.250 ;
        RECT 1676.340 1015.930 1676.600 1016.250 ;
        RECT 1676.790 1016.075 1677.070 1016.445 ;
        RECT 1676.400 1015.765 1676.540 1015.930 ;
        RECT 1661.620 1015.250 1661.880 1015.570 ;
        RECT 1669.430 1015.395 1669.710 1015.765 ;
        RECT 1676.330 1015.395 1676.610 1015.765 ;
        RECT 1682.380 1015.570 1682.520 1018.650 ;
        RECT 1683.230 1016.755 1683.510 1017.125 ;
        RECT 1683.240 1016.610 1683.500 1016.755 ;
        RECT 1683.760 1016.445 1683.900 1193.070 ;
        RECT 1691.120 1187.950 1691.260 1200.000 ;
        RECT 1704.000 1193.730 1704.140 1200.000 ;
        RECT 1703.940 1193.410 1704.200 1193.730 ;
        RECT 1716.880 1193.050 1717.020 1200.000 ;
        RECT 1716.820 1192.730 1717.080 1193.050 ;
        RECT 1729.760 1192.710 1729.900 1200.000 ;
        RECT 1729.700 1192.390 1729.960 1192.710 ;
        RECT 1735.220 1192.050 1735.480 1192.370 ;
        RECT 1721.420 1191.710 1721.680 1192.030 ;
        RECT 1707.620 1191.370 1707.880 1191.690 ;
        RECT 1693.820 1191.030 1694.080 1191.350 ;
        RECT 1691.060 1187.630 1691.320 1187.950 ;
        RECT 1690.600 1017.290 1690.860 1017.610 ;
        RECT 1691.060 1017.290 1691.320 1017.610 ;
        RECT 1689.680 1016.950 1689.940 1017.270 ;
        RECT 1690.660 1017.125 1690.800 1017.290 ;
        RECT 1683.690 1016.075 1683.970 1016.445 ;
        RECT 1682.320 1015.250 1682.580 1015.570 ;
        RECT 1683.240 1015.250 1683.500 1015.570 ;
        RECT 1683.300 1015.085 1683.440 1015.250 ;
        RECT 1689.740 1015.085 1689.880 1016.950 ;
        RECT 1690.590 1016.755 1690.870 1017.125 ;
        RECT 1691.120 1015.910 1691.260 1017.290 ;
        RECT 1693.880 1015.910 1694.020 1191.030 ;
        RECT 1700.720 1190.690 1700.980 1191.010 ;
        RECT 1700.780 1018.970 1700.920 1190.690 ;
        RECT 1700.260 1018.650 1700.520 1018.970 ;
        RECT 1700.720 1018.650 1700.980 1018.970 ;
        RECT 1700.320 1018.370 1700.460 1018.650 ;
        RECT 1703.940 1018.370 1704.200 1018.630 ;
        RECT 1700.320 1018.310 1704.200 1018.370 ;
        RECT 1700.320 1018.230 1704.140 1018.310 ;
        RECT 1704.400 1017.970 1704.660 1018.290 ;
        RECT 1697.040 1017.690 1697.300 1017.950 ;
        RECT 1704.460 1017.805 1704.600 1017.970 ;
        RECT 1697.040 1017.630 1697.700 1017.690 ;
        RECT 1696.120 1017.290 1696.380 1017.610 ;
        RECT 1697.100 1017.550 1697.700 1017.630 ;
        RECT 1691.060 1015.590 1691.320 1015.910 ;
        RECT 1693.820 1015.590 1694.080 1015.910 ;
        RECT 1696.180 1015.085 1696.320 1017.290 ;
        RECT 1697.560 1016.445 1697.700 1017.550 ;
        RECT 1697.950 1017.435 1698.230 1017.805 ;
        RECT 1704.390 1017.435 1704.670 1017.805 ;
        RECT 1697.960 1017.290 1698.220 1017.435 ;
        RECT 1697.490 1016.075 1697.770 1016.445 ;
        RECT 1707.680 1015.230 1707.820 1191.370 ;
        RECT 1710.840 1021.030 1711.100 1021.350 ;
        RECT 1710.900 1015.765 1711.040 1021.030 ;
        RECT 1719.120 1020.010 1719.380 1020.330 ;
        RECT 1719.180 1019.310 1719.320 1020.010 ;
        RECT 1721.480 1019.990 1721.620 1191.710 ;
        RECT 1728.780 1190.350 1729.040 1190.670 ;
        RECT 1728.320 1190.010 1728.580 1190.330 ;
        RECT 1726.940 1021.370 1727.200 1021.690 ;
        RECT 1726.480 1021.030 1726.740 1021.350 ;
        RECT 1726.540 1020.670 1726.680 1021.030 ;
        RECT 1727.000 1021.010 1727.140 1021.370 ;
        RECT 1726.940 1020.690 1727.200 1021.010 ;
        RECT 1726.480 1020.350 1726.740 1020.670 ;
        RECT 1721.420 1019.670 1721.680 1019.990 ;
        RECT 1728.380 1019.650 1728.520 1190.010 ;
        RECT 1728.840 1020.670 1728.980 1190.350 ;
        RECT 1728.780 1020.350 1729.040 1020.670 ;
        RECT 1732.000 1020.010 1732.260 1020.330 ;
        RECT 1725.100 1019.330 1725.360 1019.650 ;
        RECT 1728.320 1019.330 1728.580 1019.650 ;
        RECT 1718.200 1018.990 1718.460 1019.310 ;
        RECT 1719.120 1018.990 1719.380 1019.310 ;
        RECT 1711.300 1018.485 1711.560 1018.630 ;
        RECT 1718.260 1018.485 1718.400 1018.990 ;
        RECT 1711.290 1018.115 1711.570 1018.485 ;
        RECT 1718.190 1018.115 1718.470 1018.485 ;
        RECT 1724.640 1018.310 1724.900 1018.630 ;
        RECT 1712.220 1016.270 1712.480 1016.590 ;
        RECT 1710.830 1015.395 1711.110 1015.765 ;
        RECT 1683.230 1014.715 1683.510 1015.085 ;
        RECT 1689.670 1014.715 1689.950 1015.085 ;
        RECT 1696.110 1014.715 1696.390 1015.085 ;
        RECT 1707.620 1014.910 1707.880 1015.230 ;
        RECT 1579.740 1014.230 1580.000 1014.550 ;
        RECT 1710.900 1014.210 1711.040 1015.395 ;
        RECT 1712.280 1015.085 1712.420 1016.270 ;
        RECT 1718.200 1015.930 1718.460 1016.250 ;
        RECT 1718.260 1015.085 1718.400 1015.930 ;
        RECT 1724.700 1015.570 1724.840 1018.310 ;
        RECT 1725.160 1016.445 1725.300 1019.330 ;
        RECT 1729.700 1016.610 1729.960 1016.930 ;
        RECT 1725.090 1016.075 1725.370 1016.445 ;
        RECT 1724.640 1015.250 1724.900 1015.570 ;
        RECT 1724.700 1015.085 1724.840 1015.250 ;
        RECT 1729.760 1015.085 1729.900 1016.610 ;
        RECT 1732.060 1015.765 1732.200 1020.010 ;
        RECT 1733.840 1017.690 1734.100 1017.950 ;
        RECT 1734.760 1017.690 1735.020 1017.950 ;
        RECT 1733.840 1017.630 1735.020 1017.690 ;
        RECT 1733.900 1017.550 1734.960 1017.630 ;
        RECT 1735.280 1017.270 1735.420 1192.050 ;
        RECT 1738.900 1018.990 1739.160 1019.310 ;
        RECT 1735.680 1017.290 1735.940 1017.610 ;
        RECT 1735.220 1016.950 1735.480 1017.270 ;
        RECT 1731.990 1015.395 1732.270 1015.765 ;
        RECT 1735.740 1015.085 1735.880 1017.290 ;
        RECT 1738.960 1015.765 1739.100 1018.990 ;
        RECT 1741.660 1017.630 1741.920 1017.950 ;
        RECT 1745.400 1017.805 1745.540 1200.470 ;
        RECT 1755.490 1200.000 1755.770 1204.000 ;
        RECT 1768.370 1200.000 1768.650 1204.000 ;
        RECT 1780.790 1200.000 1781.070 1204.000 ;
        RECT 1793.670 1200.000 1793.950 1204.000 ;
        RECT 1806.550 1200.000 1806.830 1204.000 ;
        RECT 1819.430 1200.610 1819.710 1204.000 ;
        RECT 1832.310 1200.610 1832.590 1204.000 ;
        RECT 1819.430 1200.470 1821.440 1200.610 ;
        RECT 1819.430 1200.000 1819.710 1200.470 ;
        RECT 1755.520 1187.270 1755.660 1200.000 ;
        RECT 1768.400 1190.330 1768.540 1200.000 ;
        RECT 1780.820 1190.670 1780.960 1200.000 ;
        RECT 1780.760 1190.350 1781.020 1190.670 ;
        RECT 1768.340 1190.010 1768.600 1190.330 ;
        RECT 1755.460 1186.950 1755.720 1187.270 ;
        RECT 1759.140 1186.950 1759.400 1187.270 ;
        RECT 1745.800 1021.030 1746.060 1021.350 ;
        RECT 1745.860 1018.485 1746.000 1021.030 ;
        RECT 1746.260 1020.010 1746.520 1020.330 ;
        RECT 1745.790 1018.115 1746.070 1018.485 ;
        RECT 1746.320 1018.290 1746.460 1020.010 ;
        RECT 1755.460 1019.670 1755.720 1019.990 ;
        RECT 1758.680 1019.670 1758.940 1019.990 ;
        RECT 1755.520 1018.485 1755.660 1019.670 ;
        RECT 1746.260 1017.970 1746.520 1018.290 ;
        RECT 1746.720 1017.970 1746.980 1018.290 ;
        RECT 1755.000 1017.970 1755.260 1018.290 ;
        RECT 1755.450 1018.115 1755.730 1018.485 ;
        RECT 1738.890 1015.395 1739.170 1015.765 ;
        RECT 1741.720 1015.085 1741.860 1017.630 ;
        RECT 1745.330 1017.435 1745.610 1017.805 ;
        RECT 1745.800 1016.950 1746.060 1017.270 ;
        RECT 1745.860 1016.445 1746.000 1016.950 ;
        RECT 1745.790 1016.075 1746.070 1016.445 ;
        RECT 1746.320 1015.085 1746.460 1017.970 ;
        RECT 1711.290 1014.715 1711.570 1015.085 ;
        RECT 1712.210 1014.715 1712.490 1015.085 ;
        RECT 1718.190 1014.715 1718.470 1015.085 ;
        RECT 1724.630 1014.715 1724.910 1015.085 ;
        RECT 1729.690 1014.715 1729.970 1015.085 ;
        RECT 1735.670 1014.715 1735.950 1015.085 ;
        RECT 1741.650 1014.715 1741.930 1015.085 ;
        RECT 1746.250 1014.715 1746.530 1015.085 ;
        RECT 1711.360 1014.550 1711.500 1014.715 ;
        RECT 1746.780 1014.550 1746.920 1017.970 ;
        RECT 1755.060 1015.570 1755.200 1017.970 ;
        RECT 1758.740 1016.590 1758.880 1019.670 ;
        RECT 1759.200 1018.485 1759.340 1186.950 ;
        RECT 1787.200 1020.690 1787.460 1021.010 ;
        RECT 1759.600 1020.350 1759.860 1020.670 ;
        RECT 1759.130 1018.115 1759.410 1018.485 ;
        RECT 1758.680 1016.270 1758.940 1016.590 ;
        RECT 1755.000 1015.250 1755.260 1015.570 ;
        RECT 1755.060 1015.085 1755.200 1015.250 ;
        RECT 1758.740 1015.085 1758.880 1016.270 ;
        RECT 1759.660 1015.765 1759.800 1020.350 ;
        RECT 1773.400 1018.650 1773.660 1018.970 ;
        RECT 1778.000 1018.650 1778.260 1018.970 ;
        RECT 1771.560 1018.310 1771.820 1018.630 ;
        RECT 1766.040 1017.970 1766.300 1018.290 ;
        RECT 1766.100 1016.250 1766.240 1017.970 ;
        RECT 1766.040 1015.930 1766.300 1016.250 ;
        RECT 1766.100 1015.765 1766.240 1015.930 ;
        RECT 1759.590 1015.395 1759.870 1015.765 ;
        RECT 1766.030 1015.395 1766.310 1015.765 ;
        RECT 1766.500 1015.085 1766.760 1015.230 ;
        RECT 1771.620 1015.085 1771.760 1018.310 ;
        RECT 1773.460 1015.765 1773.600 1018.650 ;
        RECT 1778.060 1016.930 1778.200 1018.650 ;
        RECT 1782.140 1016.950 1782.400 1017.270 ;
        RECT 1787.260 1017.125 1787.400 1020.690 ;
        RECT 1787.660 1020.010 1787.920 1020.330 ;
        RECT 1778.000 1016.610 1778.260 1016.930 ;
        RECT 1773.390 1015.395 1773.670 1015.765 ;
        RECT 1778.060 1015.085 1778.200 1016.610 ;
        RECT 1780.300 1015.765 1780.560 1015.910 ;
        RECT 1780.290 1015.395 1780.570 1015.765 ;
        RECT 1782.200 1015.085 1782.340 1016.950 ;
        RECT 1787.190 1016.755 1787.470 1017.125 ;
        RECT 1787.720 1016.590 1787.860 1020.010 ;
        RECT 1789.040 1017.630 1789.300 1017.950 ;
        RECT 1787.660 1016.270 1787.920 1016.590 ;
        RECT 1789.100 1015.765 1789.240 1017.630 ;
        RECT 1793.700 1016.930 1793.840 1200.000 ;
        RECT 1806.580 1187.270 1806.720 1200.000 ;
        RECT 1806.520 1186.950 1806.780 1187.270 ;
        RECT 1811.120 1186.950 1811.380 1187.270 ;
        RECT 1811.180 1021.010 1811.320 1186.950 ;
        RECT 1821.300 1021.350 1821.440 1200.470 ;
        RECT 1831.880 1200.470 1832.590 1200.610 ;
        RECT 1821.240 1021.030 1821.500 1021.350 ;
        RECT 1828.600 1021.030 1828.860 1021.350 ;
        RECT 1831.880 1021.205 1832.020 1200.470 ;
        RECT 1832.310 1200.000 1832.590 1200.470 ;
        RECT 1845.190 1200.610 1845.470 1204.000 ;
        RECT 1845.190 1200.470 1849.040 1200.610 ;
        RECT 1845.190 1200.000 1845.470 1200.470 ;
        RECT 1848.900 1024.750 1849.040 1200.470 ;
        RECT 1858.070 1200.000 1858.350 1204.000 ;
        RECT 1870.950 1200.000 1871.230 1204.000 ;
        RECT 1883.830 1200.000 1884.110 1204.000 ;
        RECT 1896.710 1200.610 1896.990 1204.000 ;
        RECT 1909.590 1200.610 1909.870 1204.000 ;
        RECT 1896.710 1200.470 1897.340 1200.610 ;
        RECT 1896.710 1200.000 1896.990 1200.470 ;
        RECT 1855.740 1191.710 1856.000 1192.030 ;
        RECT 1848.840 1024.430 1849.100 1024.750 ;
        RECT 1855.800 1021.205 1855.940 1191.710 ;
        RECT 1858.100 1187.270 1858.240 1200.000 ;
        RECT 1870.980 1187.270 1871.120 1200.000 ;
        RECT 1883.860 1187.270 1884.000 1200.000 ;
        RECT 1858.040 1186.950 1858.300 1187.270 ;
        RECT 1862.640 1186.950 1862.900 1187.270 ;
        RECT 1870.920 1186.950 1871.180 1187.270 ;
        RECT 1876.440 1186.950 1876.700 1187.270 ;
        RECT 1883.800 1186.950 1884.060 1187.270 ;
        RECT 1890.240 1186.950 1890.500 1187.270 ;
        RECT 1811.120 1020.690 1811.380 1021.010 ;
        RECT 1800.080 1020.010 1800.340 1020.330 ;
        RECT 1793.640 1016.610 1793.900 1016.930 ;
        RECT 1793.180 1016.270 1793.440 1016.590 ;
        RECT 1789.030 1015.395 1789.310 1015.765 ;
        RECT 1793.240 1015.085 1793.380 1016.270 ;
        RECT 1800.140 1015.570 1800.280 1020.010 ;
        RECT 1806.520 1019.670 1806.780 1019.990 ;
        RECT 1828.660 1019.845 1828.800 1021.030 ;
        RECT 1831.810 1020.835 1832.090 1021.205 ;
        RECT 1835.500 1020.690 1835.760 1021.010 ;
        RECT 1855.730 1020.835 1856.010 1021.205 ;
        RECT 1835.560 1020.525 1835.700 1020.690 ;
        RECT 1835.490 1020.155 1835.770 1020.525 ;
        RECT 1800.080 1015.250 1800.340 1015.570 ;
        RECT 1800.140 1015.085 1800.280 1015.250 ;
        RECT 1806.580 1015.085 1806.720 1019.670 ;
        RECT 1821.700 1019.330 1821.960 1019.650 ;
        RECT 1828.590 1019.475 1828.870 1019.845 ;
        RECT 1817.560 1018.990 1817.820 1019.310 ;
        RECT 1821.760 1019.165 1821.900 1019.330 ;
        RECT 1812.500 1017.970 1812.760 1018.290 ;
        RECT 1812.560 1015.085 1812.700 1017.970 ;
        RECT 1817.620 1015.085 1817.760 1018.990 ;
        RECT 1821.690 1018.795 1821.970 1019.165 ;
        RECT 1823.540 1018.650 1823.800 1018.970 ;
        RECT 1823.600 1015.085 1823.740 1018.650 ;
        RECT 1842.400 1016.610 1842.660 1016.930 ;
        RECT 1842.460 1016.445 1842.600 1016.610 ;
        RECT 1842.390 1016.075 1842.670 1016.445 ;
        RECT 1754.990 1014.715 1755.270 1015.085 ;
        RECT 1758.670 1014.715 1758.950 1015.085 ;
        RECT 1766.490 1014.715 1766.770 1015.085 ;
        RECT 1771.550 1014.715 1771.830 1015.085 ;
        RECT 1777.990 1014.715 1778.270 1015.085 ;
        RECT 1782.130 1014.715 1782.410 1015.085 ;
        RECT 1787.190 1014.715 1787.470 1015.085 ;
        RECT 1793.170 1014.715 1793.450 1015.085 ;
        RECT 1800.070 1014.715 1800.350 1015.085 ;
        RECT 1806.510 1014.715 1806.790 1015.085 ;
        RECT 1812.490 1014.715 1812.770 1015.085 ;
        RECT 1817.550 1014.715 1817.830 1015.085 ;
        RECT 1823.530 1014.715 1823.810 1015.085 ;
        RECT 1787.200 1014.570 1787.460 1014.715 ;
        RECT 1711.300 1014.230 1711.560 1014.550 ;
        RECT 1746.720 1014.230 1746.980 1014.550 ;
        RECT 1710.840 1013.890 1711.100 1014.210 ;
        RECT 1862.700 1004.690 1862.840 1186.950 ;
        RECT 1876.500 1005.030 1876.640 1186.950 ;
        RECT 1890.300 1005.370 1890.440 1186.950 ;
        RECT 1897.200 1005.710 1897.340 1200.470 ;
        RECT 1909.590 1200.470 1911.140 1200.610 ;
        RECT 1909.590 1200.000 1909.870 1200.470 ;
        RECT 1901.740 1192.390 1902.000 1192.710 ;
        RECT 1901.280 1192.050 1901.540 1192.370 ;
        RECT 1900.820 1190.690 1901.080 1191.010 ;
        RECT 1897.140 1005.390 1897.400 1005.710 ;
        RECT 1890.240 1005.050 1890.500 1005.370 ;
        RECT 1876.440 1004.710 1876.700 1005.030 ;
        RECT 1862.640 1004.370 1862.900 1004.690 ;
        RECT 1489.110 558.435 1489.390 558.805 ;
        RECT 1503.830 556.395 1504.110 556.765 ;
        RECT 1503.900 554.870 1504.040 556.395 ;
      LAYER met2 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
      LAYER met2 ;
        RECT 1898.980 917.330 1899.240 917.650 ;
        RECT 1899.040 913.765 1899.180 917.330 ;
        RECT 1898.970 913.395 1899.250 913.765 ;
        RECT 1900.880 689.850 1901.020 1190.690 ;
        RECT 1900.360 689.530 1900.620 689.850 ;
        RECT 1900.820 689.530 1901.080 689.850 ;
        RECT 1900.420 676.250 1900.560 689.530 ;
        RECT 1898.980 675.930 1899.240 676.250 ;
        RECT 1900.360 675.930 1900.620 676.250 ;
        RECT 1899.040 628.165 1899.180 675.930 ;
        RECT 1898.970 627.795 1899.250 628.165 ;
        RECT 1899.890 627.795 1900.170 628.165 ;
        RECT 1899.960 596.205 1900.100 627.795 ;
        RECT 1901.340 601.645 1901.480 1192.050 ;
        RECT 1901.800 610.485 1901.940 1192.390 ;
        RECT 1902.200 1191.370 1902.460 1191.690 ;
        RECT 1902.260 904.925 1902.400 1191.370 ;
        RECT 1911.000 1010.810 1911.140 1200.470 ;
        RECT 1922.470 1200.000 1922.750 1204.000 ;
        RECT 1934.890 1200.000 1935.170 1204.000 ;
        RECT 1947.770 1200.000 1948.050 1204.000 ;
        RECT 1960.650 1200.610 1960.930 1204.000 ;
        RECT 1959.760 1200.470 1960.930 1200.610 ;
        RECT 1922.500 1191.350 1922.640 1200.000 ;
        RECT 1922.440 1191.030 1922.700 1191.350 ;
        RECT 1934.920 1187.270 1935.060 1200.000 ;
        RECT 1942.220 1192.730 1942.480 1193.050 ;
        RECT 1934.860 1186.950 1935.120 1187.270 ;
        RECT 1938.540 1186.950 1938.800 1187.270 ;
        RECT 1938.600 1011.150 1938.740 1186.950 ;
        RECT 1938.540 1010.830 1938.800 1011.150 ;
        RECT 1910.940 1010.490 1911.200 1010.810 ;
        RECT 1902.190 904.555 1902.470 904.925 ;
        RECT 1904.040 620.510 1904.300 620.830 ;
        RECT 1904.100 615.925 1904.240 620.510 ;
        RECT 1904.030 615.555 1904.310 615.925 ;
        RECT 1901.730 610.115 1902.010 610.485 ;
        RECT 1901.270 601.275 1901.550 601.645 ;
        RECT 1899.890 595.835 1900.170 596.205 ;
        RECT 1942.280 592.270 1942.420 1192.730 ;
        RECT 1947.800 1192.030 1947.940 1200.000 ;
        RECT 1956.020 1193.070 1956.280 1193.390 ;
        RECT 1947.740 1191.710 1948.000 1192.030 ;
        RECT 1904.040 591.950 1904.300 592.270 ;
        RECT 1942.220 591.950 1942.480 592.270 ;
        RECT 1904.100 590.765 1904.240 591.950 ;
        RECT 1904.030 590.395 1904.310 590.765 ;
        RECT 1903.580 579.370 1903.840 579.690 ;
        RECT 1903.640 573.765 1903.780 579.370 ;
        RECT 1956.080 579.350 1956.220 1193.070 ;
        RECT 1959.760 620.830 1959.900 1200.470 ;
        RECT 1960.650 1200.000 1960.930 1200.470 ;
        RECT 1973.530 1200.000 1973.810 1204.000 ;
        RECT 1986.410 1200.000 1986.690 1204.000 ;
        RECT 1999.290 1200.000 1999.570 1204.000 ;
        RECT 2012.170 1200.000 2012.450 1204.000 ;
        RECT 2025.050 1200.000 2025.330 1204.000 ;
        RECT 2037.930 1200.000 2038.210 1204.000 ;
        RECT 2050.810 1200.610 2051.090 1204.000 ;
        RECT 2049.460 1200.470 2051.090 1200.610 ;
        RECT 1973.560 1192.710 1973.700 1200.000 ;
        RECT 1973.500 1192.390 1973.760 1192.710 ;
        RECT 1986.440 1192.370 1986.580 1200.000 ;
        RECT 1986.380 1192.050 1986.640 1192.370 ;
        RECT 1969.820 1191.710 1970.080 1192.030 ;
        RECT 1959.700 620.510 1959.960 620.830 ;
        RECT 1969.880 579.690 1970.020 1191.710 ;
        RECT 1999.320 1191.010 1999.460 1200.000 ;
        RECT 2012.200 1193.050 2012.340 1200.000 ;
        RECT 2025.080 1193.390 2025.220 1200.000 ;
        RECT 2025.020 1193.070 2025.280 1193.390 ;
        RECT 2012.140 1192.730 2012.400 1193.050 ;
        RECT 2037.960 1192.030 2038.100 1200.000 ;
        RECT 2037.900 1191.710 2038.160 1192.030 ;
        RECT 1999.260 1190.690 1999.520 1191.010 ;
        RECT 2049.460 1014.210 2049.600 1200.470 ;
        RECT 2050.810 1200.000 2051.090 1200.470 ;
        RECT 2063.690 1200.000 2063.970 1204.000 ;
        RECT 2076.570 1200.000 2076.850 1204.000 ;
        RECT 2088.990 1200.000 2089.270 1204.000 ;
        RECT 2101.870 1200.000 2102.150 1204.000 ;
        RECT 2114.750 1200.000 2115.030 1204.000 ;
        RECT 2127.630 1200.000 2127.910 1204.000 ;
        RECT 2140.510 1200.000 2140.790 1204.000 ;
        RECT 2153.390 1200.000 2153.670 1204.000 ;
        RECT 2166.270 1200.000 2166.550 1204.000 ;
        RECT 2179.150 1200.000 2179.430 1204.000 ;
        RECT 2192.030 1200.610 2192.310 1204.000 ;
        RECT 2204.910 1200.610 2205.190 1204.000 ;
        RECT 2217.790 1200.610 2218.070 1204.000 ;
        RECT 2230.670 1200.610 2230.950 1204.000 ;
        RECT 2243.090 1200.610 2243.370 1204.000 ;
        RECT 2255.970 1200.610 2256.250 1204.000 ;
        RECT 2268.850 1200.610 2269.130 1204.000 ;
        RECT 2281.730 1200.610 2282.010 1204.000 ;
        RECT 2187.460 1200.470 2192.310 1200.610 ;
        RECT 2063.720 1191.010 2063.860 1200.000 ;
        RECT 2076.600 1191.690 2076.740 1200.000 ;
        RECT 2089.020 1192.370 2089.160 1200.000 ;
        RECT 2101.900 1192.710 2102.040 1200.000 ;
        RECT 2101.840 1192.390 2102.100 1192.710 ;
        RECT 2088.960 1192.050 2089.220 1192.370 ;
        RECT 2114.780 1192.030 2114.920 1200.000 ;
        RECT 2114.720 1191.710 2114.980 1192.030 ;
        RECT 2127.660 1191.690 2127.800 1200.000 ;
        RECT 2140.540 1193.050 2140.680 1200.000 ;
        RECT 2153.420 1193.390 2153.560 1200.000 ;
        RECT 2166.300 1193.730 2166.440 1200.000 ;
        RECT 2166.240 1193.410 2166.500 1193.730 ;
        RECT 2153.360 1193.070 2153.620 1193.390 ;
        RECT 2140.480 1192.730 2140.740 1193.050 ;
        RECT 2076.540 1191.370 2076.800 1191.690 ;
        RECT 2127.600 1191.370 2127.860 1191.690 ;
        RECT 2063.660 1190.690 2063.920 1191.010 ;
        RECT 2179.180 1189.990 2179.320 1200.000 ;
        RECT 2179.120 1189.670 2179.380 1189.990 ;
        RECT 2187.460 1018.970 2187.600 1200.470 ;
        RECT 2192.030 1200.000 2192.310 1200.470 ;
        RECT 2201.260 1200.470 2205.190 1200.610 ;
        RECT 2201.260 1019.310 2201.400 1200.470 ;
        RECT 2204.910 1200.000 2205.190 1200.470 ;
        RECT 2215.060 1200.470 2218.070 1200.610 ;
        RECT 2201.200 1018.990 2201.460 1019.310 ;
        RECT 2187.400 1018.650 2187.660 1018.970 ;
        RECT 2215.060 1018.290 2215.200 1200.470 ;
        RECT 2217.790 1200.000 2218.070 1200.470 ;
        RECT 2228.860 1200.470 2230.950 1200.610 ;
        RECT 2228.860 1019.990 2229.000 1200.470 ;
        RECT 2230.670 1200.000 2230.950 1200.470 ;
        RECT 2242.660 1200.470 2243.370 1200.610 ;
        RECT 2238.920 1191.030 2239.180 1191.350 ;
        RECT 2228.800 1019.670 2229.060 1019.990 ;
        RECT 2215.000 1017.970 2215.260 1018.290 ;
        RECT 2049.400 1013.890 2049.660 1014.210 ;
        RECT 2052.620 1013.890 2052.880 1014.210 ;
        RECT 2052.680 1008.090 2052.820 1013.890 ;
        RECT 2052.620 1007.770 2052.880 1008.090 ;
        RECT 2052.680 917.650 2052.820 1007.770 ;
        RECT 2238.980 1006.050 2239.120 1191.030 ;
        RECT 2239.380 1189.670 2239.640 1189.990 ;
        RECT 2239.440 1018.970 2239.580 1189.670 ;
        RECT 2242.660 1020.330 2242.800 1200.470 ;
        RECT 2243.090 1200.000 2243.370 1200.470 ;
        RECT 2249.560 1200.470 2256.250 1200.610 ;
        RECT 2245.820 1193.410 2246.080 1193.730 ;
        RECT 2245.880 1020.330 2246.020 1193.410 ;
        RECT 2249.040 1020.525 2249.300 1020.670 ;
        RECT 2242.600 1020.010 2242.860 1020.330 ;
        RECT 2245.820 1020.010 2246.080 1020.330 ;
        RECT 2249.030 1020.155 2249.310 1020.525 ;
        RECT 2239.380 1018.650 2239.640 1018.970 ;
        RECT 2242.140 1018.650 2242.400 1018.970 ;
        RECT 2242.200 1007.605 2242.340 1018.650 ;
        RECT 2245.880 1017.125 2246.020 1020.010 ;
        RECT 2245.810 1016.755 2246.090 1017.125 ;
        RECT 2249.560 1016.590 2249.700 1200.470 ;
        RECT 2255.970 1200.000 2256.250 1200.470 ;
        RECT 2263.360 1200.470 2269.130 1200.610 ;
        RECT 2252.720 1193.070 2252.980 1193.390 ;
        RECT 2252.780 1019.650 2252.920 1193.070 ;
        RECT 2259.620 1192.730 2259.880 1193.050 ;
        RECT 2255.940 1191.030 2256.200 1191.350 ;
        RECT 2252.720 1019.330 2252.980 1019.650 ;
        RECT 2252.780 1017.125 2252.920 1019.330 ;
        RECT 2252.710 1016.755 2252.990 1017.125 ;
        RECT 2249.500 1016.270 2249.760 1016.590 ;
        RECT 2256.000 1016.445 2256.140 1191.030 ;
        RECT 2259.680 1019.310 2259.820 1192.730 ;
        RECT 2259.620 1018.990 2259.880 1019.310 ;
        RECT 2259.680 1017.125 2259.820 1018.990 ;
        RECT 2263.360 1017.950 2263.500 1200.470 ;
        RECT 2268.850 1200.000 2269.130 1200.470 ;
        RECT 2277.160 1200.470 2282.010 1200.610 ;
        RECT 2273.420 1191.710 2273.680 1192.030 ;
        RECT 2276.180 1191.710 2276.440 1192.030 ;
        RECT 2266.520 1191.370 2266.780 1191.690 ;
        RECT 2269.740 1191.370 2270.000 1191.690 ;
        RECT 2263.300 1017.630 2263.560 1017.950 ;
        RECT 2266.580 1017.125 2266.720 1191.370 ;
        RECT 2259.610 1016.755 2259.890 1017.125 ;
        RECT 2266.510 1016.755 2266.790 1017.125 ;
        RECT 2255.930 1016.075 2256.210 1016.445 ;
        RECT 2266.580 1015.570 2266.720 1016.755 ;
        RECT 2269.800 1016.445 2269.940 1191.370 ;
        RECT 2273.480 1016.445 2273.620 1191.710 ;
        RECT 2276.240 1016.445 2276.380 1191.710 ;
        RECT 2277.160 1017.270 2277.300 1200.470 ;
        RECT 2281.730 1200.000 2282.010 1200.470 ;
        RECT 2294.610 1200.000 2294.890 1204.000 ;
        RECT 2307.490 1200.000 2307.770 1204.000 ;
        RECT 2320.370 1200.000 2320.650 1204.000 ;
        RECT 2333.250 1200.000 2333.530 1204.000 ;
        RECT 2346.130 1200.000 2346.410 1204.000 ;
        RECT 2359.010 1200.000 2359.290 1204.000 ;
        RECT 2371.890 1200.000 2372.170 1204.000 ;
        RECT 2384.770 1200.610 2385.050 1204.000 ;
        RECT 2384.340 1200.470 2385.050 1200.610 ;
        RECT 2294.640 1193.390 2294.780 1200.000 ;
        RECT 2294.580 1193.070 2294.840 1193.390 ;
        RECT 2281.240 1192.390 2281.500 1192.710 ;
        RECT 2304.240 1192.390 2304.500 1192.710 ;
        RECT 2280.320 1192.050 2280.580 1192.370 ;
        RECT 2280.380 1021.350 2280.520 1192.050 ;
        RECT 2280.320 1021.030 2280.580 1021.350 ;
        RECT 2281.300 1017.690 2281.440 1192.390 ;
        RECT 2290.440 1192.050 2290.700 1192.370 ;
        RECT 2283.080 1021.205 2283.340 1021.350 ;
        RECT 2283.070 1020.835 2283.350 1021.205 ;
        RECT 2289.980 1018.650 2290.240 1018.970 ;
        RECT 2280.840 1017.550 2281.440 1017.690 ;
        RECT 2280.840 1017.270 2280.980 1017.550 ;
        RECT 2277.100 1016.950 2277.360 1017.270 ;
        RECT 2280.780 1017.125 2281.040 1017.270 ;
        RECT 2280.770 1016.755 2281.050 1017.125 ;
        RECT 2290.040 1016.930 2290.180 1018.650 ;
        RECT 2289.980 1016.610 2290.240 1016.930 ;
        RECT 2269.730 1016.075 2270.010 1016.445 ;
        RECT 2273.410 1016.075 2273.690 1016.445 ;
        RECT 2275.250 1016.075 2275.530 1016.445 ;
        RECT 2276.170 1016.075 2276.450 1016.445 ;
        RECT 2275.320 1015.910 2275.460 1016.075 ;
        RECT 2275.260 1015.590 2275.520 1015.910 ;
        RECT 2266.520 1015.250 2266.780 1015.570 ;
        RECT 2276.640 1015.085 2276.900 1015.230 ;
        RECT 2290.040 1015.085 2290.180 1016.610 ;
        RECT 2290.500 1016.445 2290.640 1192.050 ;
        RECT 2295.040 1020.010 2295.300 1020.330 ;
        RECT 2290.430 1016.075 2290.710 1016.445 ;
        RECT 2295.100 1015.085 2295.240 1020.010 ;
        RECT 2297.340 1019.670 2297.600 1019.990 ;
        RECT 2297.400 1017.125 2297.540 1019.670 ;
        RECT 2302.860 1019.330 2303.120 1019.650 ;
        RECT 2302.920 1017.270 2303.060 1019.330 ;
        RECT 2297.330 1016.755 2297.610 1017.125 ;
        RECT 2302.860 1016.950 2303.120 1017.270 ;
        RECT 2302.920 1015.085 2303.060 1016.950 ;
        RECT 2304.300 1016.445 2304.440 1192.390 ;
        RECT 2307.520 1187.270 2307.660 1200.000 ;
        RECT 2320.400 1193.730 2320.540 1200.000 ;
        RECT 2320.340 1193.410 2320.600 1193.730 ;
        RECT 2318.040 1192.730 2318.300 1193.050 ;
        RECT 2307.460 1186.950 2307.720 1187.270 ;
        RECT 2311.140 1186.950 2311.400 1187.270 ;
        RECT 2310.680 1019.330 2310.940 1019.650 ;
        RECT 2307.000 1018.990 2307.260 1019.310 ;
        RECT 2307.060 1017.950 2307.200 1018.990 ;
        RECT 2307.000 1017.630 2307.260 1017.950 ;
        RECT 2304.230 1016.075 2304.510 1016.445 ;
        RECT 2307.060 1015.085 2307.200 1017.630 ;
        RECT 2310.740 1017.125 2310.880 1019.330 ;
        RECT 2311.200 1018.630 2311.340 1186.950 ;
        RECT 2317.580 1018.990 2317.840 1019.310 ;
        RECT 2311.140 1018.310 2311.400 1018.630 ;
        RECT 2317.640 1017.125 2317.780 1018.990 ;
        RECT 2310.670 1016.755 2310.950 1017.125 ;
        RECT 2317.570 1016.755 2317.850 1017.125 ;
        RECT 2318.100 1016.445 2318.240 1192.730 ;
        RECT 2333.280 1189.310 2333.420 1200.000 ;
        RECT 2333.220 1188.990 2333.480 1189.310 ;
        RECT 2346.160 1188.970 2346.300 1200.000 ;
        RECT 2346.100 1188.650 2346.360 1188.970 ;
        RECT 2359.040 1188.290 2359.180 1200.000 ;
        RECT 2359.440 1189.670 2359.700 1189.990 ;
        RECT 2358.980 1187.970 2359.240 1188.290 ;
        RECT 2352.540 1025.790 2352.800 1026.110 ;
        RECT 2352.080 1025.110 2352.340 1025.430 ;
        RECT 2345.640 1024.770 2345.900 1025.090 ;
        RECT 2325.400 1021.030 2325.660 1021.350 ;
        RECT 2345.700 1021.205 2345.840 1024.770 ;
        RECT 2324.940 1018.650 2325.200 1018.970 ;
        RECT 2323.100 1016.445 2323.360 1016.590 ;
        RECT 2318.030 1016.075 2318.310 1016.445 ;
        RECT 2323.090 1016.075 2323.370 1016.445 ;
        RECT 2318.040 1015.590 2318.300 1015.910 ;
        RECT 2312.060 1015.250 2312.320 1015.570 ;
        RECT 2312.120 1015.085 2312.260 1015.250 ;
        RECT 2318.100 1015.085 2318.240 1015.590 ;
        RECT 2325.000 1015.085 2325.140 1018.650 ;
        RECT 2325.460 1016.445 2325.600 1021.030 ;
        RECT 2338.740 1020.690 2339.000 1021.010 ;
        RECT 2345.630 1020.835 2345.910 1021.205 ;
        RECT 2338.800 1020.525 2338.940 1020.690 ;
        RECT 2352.140 1020.525 2352.280 1025.110 ;
        RECT 2352.600 1021.205 2352.740 1025.790 ;
        RECT 2352.530 1020.835 2352.810 1021.205 ;
        RECT 2325.860 1020.010 2326.120 1020.330 ;
        RECT 2332.760 1020.010 2333.020 1020.330 ;
        RECT 2338.730 1020.155 2339.010 1020.525 ;
        RECT 2352.070 1020.155 2352.350 1020.525 ;
        RECT 2325.920 1017.270 2326.060 1020.010 ;
        RECT 2331.900 1018.290 2332.500 1018.370 ;
        RECT 2331.900 1018.230 2332.560 1018.290 ;
        RECT 2325.860 1016.950 2326.120 1017.270 ;
        RECT 2325.390 1016.075 2325.670 1016.445 ;
        RECT 2331.900 1015.085 2332.040 1018.230 ;
        RECT 2332.300 1017.970 2332.560 1018.230 ;
        RECT 2332.820 1017.690 2332.960 1020.010 ;
        RECT 2332.360 1017.550 2332.960 1017.690 ;
        RECT 2353.460 1017.630 2353.720 1017.950 ;
        RECT 2332.360 1016.590 2332.500 1017.550 ;
        RECT 2347.020 1017.290 2347.280 1017.610 ;
        RECT 2342.420 1016.950 2342.680 1017.270 ;
        RECT 2336.440 1016.610 2336.700 1016.930 ;
        RECT 2332.300 1016.270 2332.560 1016.590 ;
        RECT 2332.760 1016.445 2333.020 1016.590 ;
        RECT 2332.750 1016.075 2333.030 1016.445 ;
        RECT 2336.500 1015.085 2336.640 1016.610 ;
        RECT 2342.480 1015.085 2342.620 1016.950 ;
        RECT 2347.080 1015.085 2347.220 1017.290 ;
        RECT 2353.520 1015.085 2353.660 1017.630 ;
        RECT 2359.500 1016.445 2359.640 1189.670 ;
        RECT 2366.340 1189.330 2366.600 1189.650 ;
        RECT 2366.400 1016.445 2366.540 1189.330 ;
        RECT 2371.920 1187.270 2372.060 1200.000 ;
        RECT 2383.820 1188.990 2384.080 1189.310 ;
        RECT 2380.140 1187.630 2380.400 1187.950 ;
        RECT 2371.860 1186.950 2372.120 1187.270 ;
        RECT 2369.100 1022.050 2369.360 1022.370 ;
        RECT 2369.160 1021.010 2369.300 1022.050 ;
        RECT 2369.100 1020.690 2369.360 1021.010 ;
        RECT 2370.940 1020.010 2371.200 1020.330 ;
        RECT 2359.430 1016.075 2359.710 1016.445 ;
        RECT 2364.500 1015.930 2364.760 1016.250 ;
        RECT 2366.330 1016.075 2366.610 1016.445 ;
        RECT 2358.980 1015.250 2359.240 1015.570 ;
        RECT 2359.440 1015.250 2359.700 1015.570 ;
        RECT 2359.040 1015.085 2359.180 1015.250 ;
        RECT 2262.830 1014.715 2263.110 1015.085 ;
        RECT 2276.630 1014.715 2276.910 1015.085 ;
        RECT 2283.070 1014.715 2283.350 1015.085 ;
        RECT 2289.970 1014.715 2290.250 1015.085 ;
        RECT 2295.030 1014.715 2295.310 1015.085 ;
        RECT 2302.850 1014.715 2303.130 1015.085 ;
        RECT 2306.990 1014.715 2307.270 1015.085 ;
        RECT 2312.050 1014.715 2312.330 1015.085 ;
        RECT 2318.030 1014.715 2318.310 1015.085 ;
        RECT 2324.930 1014.715 2325.210 1015.085 ;
        RECT 2331.830 1014.715 2332.110 1015.085 ;
        RECT 2336.430 1014.715 2336.710 1015.085 ;
        RECT 2342.410 1014.715 2342.690 1015.085 ;
        RECT 2347.010 1014.715 2347.290 1015.085 ;
        RECT 2353.450 1014.715 2353.730 1015.085 ;
        RECT 2358.050 1014.970 2358.330 1015.085 ;
        RECT 2358.050 1014.830 2358.720 1014.970 ;
        RECT 2358.050 1014.715 2358.330 1014.830 ;
        RECT 2262.840 1014.570 2263.100 1014.715 ;
        RECT 2283.140 1014.550 2283.280 1014.715 ;
        RECT 2283.080 1014.230 2283.340 1014.550 ;
        RECT 2358.580 1014.290 2358.720 1014.830 ;
        RECT 2358.970 1014.715 2359.250 1015.085 ;
        RECT 2359.500 1014.290 2359.640 1015.250 ;
        RECT 2364.560 1015.085 2364.700 1015.930 ;
        RECT 2371.000 1015.085 2371.140 1020.010 ;
        RECT 2377.840 1016.270 2378.100 1016.590 ;
        RECT 2380.200 1016.445 2380.340 1187.630 ;
        RECT 2383.880 1020.330 2384.020 1188.990 ;
        RECT 2384.340 1020.525 2384.480 1200.470 ;
        RECT 2384.770 1200.000 2385.050 1200.470 ;
        RECT 2397.190 1200.000 2397.470 1204.000 ;
        RECT 2410.070 1200.000 2410.350 1204.000 ;
        RECT 2422.950 1200.000 2423.230 1204.000 ;
        RECT 2435.830 1200.000 2436.110 1204.000 ;
        RECT 2448.710 1200.610 2448.990 1204.000 ;
        RECT 2461.590 1200.610 2461.870 1204.000 ;
        RECT 2474.470 1200.610 2474.750 1204.000 ;
        RECT 2442.760 1200.470 2448.990 1200.610 ;
        RECT 2385.200 1193.410 2385.460 1193.730 ;
        RECT 2386.120 1193.410 2386.380 1193.730 ;
        RECT 2384.740 1187.290 2385.000 1187.610 ;
        RECT 2384.800 1038.885 2384.940 1187.290 ;
        RECT 2384.730 1038.515 2385.010 1038.885 ;
        RECT 2385.260 1021.350 2385.400 1193.410 ;
        RECT 2385.660 1190.010 2385.920 1190.330 ;
        RECT 2385.200 1021.030 2385.460 1021.350 ;
        RECT 2383.360 1020.010 2383.620 1020.330 ;
        RECT 2383.820 1020.010 2384.080 1020.330 ;
        RECT 2384.270 1020.155 2384.550 1020.525 ;
        RECT 2383.420 1019.845 2383.560 1020.010 ;
        RECT 2383.350 1019.475 2383.630 1019.845 ;
        RECT 2385.720 1017.270 2385.860 1190.010 ;
        RECT 2386.180 1022.370 2386.320 1193.410 ;
        RECT 2391.180 1190.350 2391.440 1190.670 ;
        RECT 2390.720 1188.650 2390.980 1188.970 ;
        RECT 2387.960 1187.970 2388.220 1188.290 ;
        RECT 2387.500 1186.950 2387.760 1187.270 ;
        RECT 2386.120 1022.050 2386.380 1022.370 ;
        RECT 2387.560 1021.205 2387.700 1186.950 ;
        RECT 2387.490 1020.835 2387.770 1021.205 ;
        RECT 2388.020 1020.525 2388.160 1187.970 ;
        RECT 2390.780 1021.205 2390.920 1188.650 ;
        RECT 2390.710 1020.835 2390.990 1021.205 ;
        RECT 2391.240 1021.010 2391.380 1190.350 ;
        RECT 2391.640 1190.010 2391.900 1190.330 ;
        RECT 2391.180 1020.690 2391.440 1021.010 ;
        RECT 2387.950 1020.155 2388.230 1020.525 ;
        RECT 2388.410 1019.475 2388.690 1019.845 ;
        RECT 2387.960 1017.290 2388.220 1017.610 ;
        RECT 2385.660 1016.950 2385.920 1017.270 ;
        RECT 2388.020 1017.125 2388.160 1017.290 ;
        RECT 2380.600 1016.610 2380.860 1016.930 ;
        RECT 2387.500 1016.610 2387.760 1016.930 ;
        RECT 2387.950 1016.755 2388.230 1017.125 ;
        RECT 2388.480 1016.930 2388.620 1019.475 ;
        RECT 2391.700 1018.290 2391.840 1190.010 ;
        RECT 2397.220 1187.950 2397.360 1200.000 ;
        RECT 2397.620 1193.070 2397.880 1193.390 ;
        RECT 2397.160 1187.630 2397.420 1187.950 ;
        RECT 2397.680 1018.290 2397.820 1193.070 ;
        RECT 2410.100 1187.610 2410.240 1200.000 ;
        RECT 2422.980 1189.650 2423.120 1200.000 ;
        RECT 2435.860 1189.990 2436.000 1200.000 ;
        RECT 2435.800 1189.670 2436.060 1189.990 ;
        RECT 2422.920 1189.330 2423.180 1189.650 ;
        RECT 2410.040 1187.290 2410.300 1187.610 ;
        RECT 2442.760 1026.110 2442.900 1200.470 ;
        RECT 2448.710 1200.000 2448.990 1200.470 ;
        RECT 2456.560 1200.470 2461.870 1200.610 ;
        RECT 2442.700 1025.790 2442.960 1026.110 ;
        RECT 2456.560 1025.430 2456.700 1200.470 ;
        RECT 2461.590 1200.000 2461.870 1200.470 ;
        RECT 2470.360 1200.470 2474.750 1200.610 ;
        RECT 2456.500 1025.110 2456.760 1025.430 ;
        RECT 2470.360 1025.090 2470.500 1200.470 ;
        RECT 2474.470 1200.000 2474.750 1200.470 ;
        RECT 2487.350 1200.000 2487.630 1204.000 ;
        RECT 2500.230 1200.000 2500.510 1204.000 ;
        RECT 2513.110 1200.610 2513.390 1204.000 ;
        RECT 2511.760 1200.470 2513.390 1200.610 ;
        RECT 2487.380 1193.730 2487.520 1200.000 ;
        RECT 2487.320 1193.410 2487.580 1193.730 ;
        RECT 2481.800 1190.690 2482.060 1191.010 ;
        RECT 2470.300 1024.770 2470.560 1025.090 ;
        RECT 2450.980 1024.430 2451.240 1024.750 ;
        RECT 2408.200 1021.205 2408.460 1021.350 ;
        RECT 2451.040 1021.205 2451.180 1024.430 ;
        RECT 2408.190 1020.835 2408.470 1021.205 ;
        RECT 2428.900 1020.690 2429.160 1021.010 ;
        RECT 2450.970 1020.835 2451.250 1021.205 ;
        RECT 2428.960 1020.525 2429.100 1020.690 ;
        RECT 2402.220 1020.010 2402.480 1020.330 ;
        RECT 2428.890 1020.155 2429.170 1020.525 ;
        RECT 2402.280 1019.845 2402.420 1020.010 ;
        RECT 2402.210 1019.475 2402.490 1019.845 ;
        RECT 2415.100 1018.485 2415.360 1018.630 ;
        RECT 2391.640 1017.970 2391.900 1018.290 ;
        RECT 2397.620 1017.970 2397.880 1018.290 ;
        RECT 2415.090 1018.115 2415.370 1018.485 ;
        RECT 2422.000 1017.970 2422.260 1018.290 ;
        RECT 2422.060 1017.805 2422.200 1017.970 ;
        RECT 2421.990 1017.435 2422.270 1017.805 ;
        RECT 2428.900 1016.950 2429.160 1017.270 ;
        RECT 2388.420 1016.610 2388.680 1016.930 ;
        RECT 2377.900 1015.085 2378.040 1016.270 ;
        RECT 2380.130 1016.075 2380.410 1016.445 ;
        RECT 2380.660 1015.085 2380.800 1016.610 ;
        RECT 2387.560 1016.445 2387.700 1016.610 ;
        RECT 2387.490 1016.075 2387.770 1016.445 ;
        RECT 2415.100 1016.270 2415.360 1016.590 ;
        RECT 2428.960 1016.445 2429.100 1016.950 ;
        RECT 2408.200 1015.590 2408.460 1015.910 ;
        RECT 2394.400 1015.250 2394.660 1015.570 ;
        RECT 2403.140 1015.250 2403.400 1015.570 ;
        RECT 2394.460 1015.085 2394.600 1015.250 ;
        RECT 2403.200 1015.085 2403.340 1015.250 ;
        RECT 2408.260 1015.085 2408.400 1015.590 ;
        RECT 2415.160 1015.085 2415.300 1016.270 ;
        RECT 2422.000 1015.930 2422.260 1016.250 ;
        RECT 2428.890 1016.075 2429.170 1016.445 ;
        RECT 2422.060 1015.085 2422.200 1015.930 ;
        RECT 2364.490 1014.715 2364.770 1015.085 ;
        RECT 2370.930 1014.715 2371.210 1015.085 ;
        RECT 2377.830 1014.715 2378.110 1015.085 ;
        RECT 2380.590 1014.715 2380.870 1015.085 ;
        RECT 2394.390 1014.715 2394.670 1015.085 ;
        RECT 2403.130 1014.715 2403.410 1015.085 ;
        RECT 2408.190 1014.715 2408.470 1015.085 ;
        RECT 2415.090 1014.715 2415.370 1015.085 ;
        RECT 2421.990 1014.715 2422.270 1015.085 ;
        RECT 2358.580 1014.150 2359.640 1014.290 ;
        RECT 2242.130 1007.235 2242.410 1007.605 ;
        RECT 2238.920 1005.730 2239.180 1006.050 ;
        RECT 2052.620 917.330 2052.880 917.650 ;
        RECT 1969.820 579.370 1970.080 579.690 ;
        RECT 1904.040 579.205 1904.300 579.350 ;
        RECT 1904.030 578.835 1904.310 579.205 ;
        RECT 1956.020 579.030 1956.280 579.350 ;
        RECT 1903.570 573.395 1903.850 573.765 ;
        RECT 2083.890 556.395 2084.170 556.765 ;
        RECT 2083.960 554.870 2084.100 556.395 ;
      LAYER met2 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met2 ;
        RECT 2481.860 906.850 2482.000 1190.690 ;
        RECT 2500.260 1190.330 2500.400 1200.000 ;
        RECT 2500.200 1190.010 2500.460 1190.330 ;
        RECT 2511.760 1018.970 2511.900 1200.470 ;
        RECT 2513.110 1200.000 2513.390 1200.470 ;
        RECT 2525.990 1200.000 2526.270 1204.000 ;
        RECT 2538.870 1200.610 2539.150 1204.000 ;
        RECT 2551.290 1200.610 2551.570 1204.000 ;
        RECT 2532.460 1200.470 2539.150 1200.610 ;
        RECT 2526.020 1193.050 2526.160 1200.000 ;
        RECT 2525.960 1192.730 2526.220 1193.050 ;
        RECT 2532.460 1019.310 2532.600 1200.470 ;
        RECT 2538.870 1200.000 2539.150 1200.470 ;
        RECT 2546.260 1200.470 2551.570 1200.610 ;
        RECT 2546.260 1019.650 2546.400 1200.470 ;
        RECT 2551.290 1200.000 2551.570 1200.470 ;
        RECT 2564.170 1200.000 2564.450 1204.000 ;
        RECT 2577.050 1200.610 2577.330 1204.000 ;
        RECT 2573.860 1200.470 2577.330 1200.610 ;
        RECT 2564.200 1192.710 2564.340 1200.000 ;
        RECT 2564.140 1192.390 2564.400 1192.710 ;
        RECT 2573.860 1019.990 2574.000 1200.470 ;
        RECT 2577.050 1200.000 2577.330 1200.470 ;
        RECT 2589.930 1200.000 2590.210 1204.000 ;
        RECT 2602.810 1200.610 2603.090 1204.000 ;
        RECT 2601.460 1200.470 2603.090 1200.610 ;
        RECT 2589.960 1192.370 2590.100 1200.000 ;
        RECT 2589.900 1192.050 2590.160 1192.370 ;
        RECT 2573.800 1019.670 2574.060 1019.990 ;
        RECT 2546.200 1019.330 2546.460 1019.650 ;
        RECT 2532.400 1018.990 2532.660 1019.310 ;
        RECT 2511.700 1018.650 2511.960 1018.970 ;
        RECT 2601.460 1014.550 2601.600 1200.470 ;
        RECT 2602.810 1200.000 2603.090 1200.470 ;
        RECT 2615.690 1200.000 2615.970 1204.000 ;
        RECT 2628.570 1200.610 2628.850 1204.000 ;
        RECT 2622.160 1200.470 2628.850 1200.610 ;
        RECT 2615.720 1192.030 2615.860 1200.000 ;
        RECT 2615.660 1191.710 2615.920 1192.030 ;
        RECT 2622.160 1015.230 2622.300 1200.470 ;
        RECT 2628.570 1200.000 2628.850 1200.470 ;
        RECT 2641.450 1200.000 2641.730 1204.000 ;
        RECT 2654.330 1200.610 2654.610 1204.000 ;
        RECT 2649.760 1200.470 2654.610 1200.610 ;
        RECT 2641.480 1191.690 2641.620 1200.000 ;
        RECT 2641.420 1191.370 2641.680 1191.690 ;
        RECT 2622.100 1014.910 2622.360 1015.230 ;
        RECT 2649.760 1014.890 2649.900 1200.470 ;
        RECT 2654.330 1200.000 2654.610 1200.470 ;
        RECT 2667.210 1200.000 2667.490 1204.000 ;
        RECT 2680.090 1200.610 2680.370 1204.000 ;
        RECT 2692.970 1200.610 2693.250 1204.000 ;
        RECT 2677.360 1200.470 2680.370 1200.610 ;
        RECT 2667.240 1191.350 2667.380 1200.000 ;
        RECT 2667.180 1191.030 2667.440 1191.350 ;
        RECT 2677.360 1020.670 2677.500 1200.470 ;
        RECT 2680.090 1200.000 2680.370 1200.470 ;
        RECT 2691.160 1200.470 2693.250 1200.610 ;
        RECT 2677.300 1020.350 2677.560 1020.670 ;
        RECT 2691.160 1019.165 2691.300 1200.470 ;
        RECT 2692.970 1200.000 2693.250 1200.470 ;
        RECT 2691.090 1018.795 2691.370 1019.165 ;
        RECT 2649.700 1014.570 2649.960 1014.890 ;
        RECT 2601.400 1014.230 2601.660 1014.550 ;
        RECT 2501.120 1010.830 2501.380 1011.150 ;
        RECT 2498.820 1010.490 2499.080 1010.810 ;
        RECT 2498.360 1005.730 2498.620 1006.050 ;
        RECT 2482.250 906.850 2482.530 906.965 ;
        RECT 2481.860 906.710 2482.530 906.850 ;
        RECT 2482.250 906.595 2482.530 906.710 ;
        RECT 2498.420 579.205 2498.560 1005.730 ;
        RECT 2498.880 590.765 2499.020 1010.490 ;
        RECT 2499.280 1005.390 2499.540 1005.710 ;
        RECT 2499.340 593.485 2499.480 1005.390 ;
        RECT 2499.740 1005.050 2500.000 1005.370 ;
        RECT 2499.800 604.365 2499.940 1005.050 ;
        RECT 2500.200 1004.710 2500.460 1005.030 ;
        RECT 2500.260 610.485 2500.400 1004.710 ;
        RECT 2500.660 1004.370 2500.920 1004.690 ;
        RECT 2500.720 618.645 2500.860 1004.370 ;
        RECT 2500.650 618.275 2500.930 618.645 ;
        RECT 2500.190 610.115 2500.470 610.485 ;
        RECT 2499.730 603.995 2500.010 604.365 ;
        RECT 2499.270 593.115 2499.550 593.485 ;
        RECT 2498.810 590.395 2499.090 590.765 ;
        RECT 2498.350 578.835 2498.630 579.205 ;
        RECT 2501.180 576.485 2501.320 1010.830 ;
        RECT 2501.580 1007.770 2501.840 1008.090 ;
        RECT 2501.640 915.805 2501.780 1007.770 ;
        RECT 2501.570 915.435 2501.850 915.805 ;
        RECT 2501.110 576.115 2501.390 576.485 ;
        RECT 1503.840 554.550 1504.100 554.870 ;
        RECT 2083.900 554.550 2084.160 554.870 ;
      LAYER via2 ;
        RECT 1868.150 3063.600 1868.430 3063.880 ;
        RECT 1490.030 3033.000 1490.310 3033.280 ;
        RECT 1489.570 3026.880 1489.850 3027.160 ;
        RECT 1489.110 3018.720 1489.390 3019.000 ;
        RECT 1488.650 3012.600 1488.930 3012.880 ;
        RECT 1488.190 3004.440 1488.470 3004.720 ;
        RECT 1487.730 2999.000 1488.010 2999.280 ;
        RECT 1487.270 2990.160 1487.550 2990.440 ;
        RECT 1486.810 2701.160 1487.090 2701.440 ;
        RECT 1486.350 2692.320 1486.630 2692.600 ;
        RECT 1318.450 2410.800 1318.730 2411.080 ;
        RECT 1572.830 2593.720 1573.110 2594.000 ;
        RECT 1600.430 2593.720 1600.710 2594.000 ;
        RECT 1614.690 2593.720 1614.970 2594.000 ;
        RECT 1621.590 2593.720 1621.870 2594.000 ;
        RECT 1627.110 2593.720 1627.390 2594.000 ;
        RECT 1632.170 2593.720 1632.450 2594.000 ;
        RECT 1636.770 2593.720 1637.050 2594.000 ;
        RECT 1644.590 2593.720 1644.870 2594.000 ;
        RECT 1537.870 2587.600 1538.150 2587.880 ;
        RECT 1565.930 2593.040 1566.210 2593.320 ;
        RECT 1586.170 2593.040 1586.450 2593.320 ;
        RECT 1593.530 2593.040 1593.810 2593.320 ;
        RECT 1605.490 2593.040 1605.770 2593.320 ;
        RECT 1615.610 2593.040 1615.890 2593.320 ;
        RECT 1573.290 2592.360 1573.570 2592.640 ;
        RECT 1580.190 2592.360 1580.470 2592.640 ;
        RECT 1566.390 2591.680 1566.670 2591.960 ;
        RECT 1586.630 2592.360 1586.910 2592.640 ;
        RECT 1587.550 2592.360 1587.830 2592.640 ;
        RECT 1579.730 2590.320 1580.010 2590.600 ;
        RECT 1587.090 2589.640 1587.370 2589.920 ;
        RECT 1593.990 2591.680 1594.270 2591.960 ;
        RECT 1600.890 2591.680 1601.170 2591.960 ;
        RECT 1608.710 2591.000 1608.990 2591.280 ;
        RECT 1593.990 2590.320 1594.270 2590.600 ;
        RECT 1627.570 2592.360 1627.850 2592.640 ;
        RECT 1650.570 2593.720 1650.850 2594.000 ;
        RECT 1656.550 2593.720 1656.830 2594.000 ;
        RECT 1662.070 2593.720 1662.350 2594.000 ;
        RECT 1668.970 2593.720 1669.250 2594.000 ;
        RECT 1673.570 2593.720 1673.850 2594.000 ;
        RECT 1679.090 2593.720 1679.370 2594.000 ;
        RECT 1684.610 2593.720 1684.890 2594.000 ;
        RECT 1690.590 2593.720 1690.870 2594.000 ;
        RECT 1697.490 2593.720 1697.770 2594.000 ;
        RECT 1703.010 2593.720 1703.290 2594.000 ;
        RECT 1707.610 2593.720 1707.890 2594.000 ;
        RECT 1726.470 2593.720 1726.750 2594.000 ;
        RECT 1732.910 2593.720 1733.190 2594.000 ;
        RECT 1744.870 2593.720 1745.150 2594.000 ;
        RECT 1657.010 2593.040 1657.290 2593.320 ;
        RECT 1649.190 2592.360 1649.470 2592.640 ;
        RECT 1560.870 2588.960 1561.150 2589.240 ;
        RECT 1551.210 2588.280 1551.490 2588.560 ;
        RECT 1545.230 2587.600 1545.510 2587.880 ;
        RECT 1551.670 2587.600 1551.950 2587.880 ;
        RECT 1559.030 2587.600 1559.310 2587.880 ;
        RECT 1600.890 2410.120 1601.170 2410.400 ;
        RECT 1607.790 2410.120 1608.070 2410.400 ;
        RECT 1622.510 2588.280 1622.790 2588.560 ;
        RECT 1622.050 2587.600 1622.330 2587.880 ;
        RECT 1628.490 2588.280 1628.770 2588.560 ;
        RECT 1635.850 2588.280 1636.130 2588.560 ;
        RECT 1642.290 2588.280 1642.570 2588.560 ;
        RECT 1663.450 2591.000 1663.730 2591.280 ;
        RECT 1662.990 2588.280 1663.270 2588.560 ;
        RECT 1683.690 2591.680 1683.970 2591.960 ;
        RECT 1697.950 2593.040 1698.230 2593.320 ;
        RECT 1690.590 2591.680 1690.870 2591.960 ;
        RECT 1697.490 2591.680 1697.770 2591.960 ;
        RECT 1704.390 2591.000 1704.670 2591.280 ;
        RECT 1714.970 2592.360 1715.250 2592.640 ;
        RECT 1718.650 2591.680 1718.930 2591.960 ;
        RECT 1738.430 2593.040 1738.710 2593.320 ;
        RECT 1738.890 2592.360 1739.170 2592.640 ;
        RECT 1669.890 2588.960 1670.170 2589.240 ;
        RECT 1711.290 2588.960 1711.570 2589.240 ;
        RECT 1676.790 2588.280 1677.070 2588.560 ;
        RECT 1718.190 2588.280 1718.470 2588.560 ;
        RECT 1726.010 2588.280 1726.290 2588.560 ;
        RECT 1731.990 2588.280 1732.270 2588.560 ;
        RECT 1739.350 2588.960 1739.630 2589.240 ;
        RECT 2442.690 3063.600 2442.970 3063.880 ;
        RECT 2469.830 3063.600 2470.110 3063.880 ;
        RECT 1898.510 3047.960 1898.790 3048.240 ;
        RECT 1899.890 3047.960 1900.170 3048.240 ;
        RECT 1898.050 2746.720 1898.330 2747.000 ;
        RECT 2083.890 3030.280 2084.170 3030.560 ;
        RECT 1898.970 2704.560 1899.250 2704.840 ;
        RECT 1898.510 2410.800 1898.790 2411.080 ;
        RECT 2083.890 3024.160 2084.170 3024.440 ;
        RECT 2083.890 3016.000 2084.170 3016.280 ;
        RECT 2083.890 3009.880 2084.170 3010.160 ;
        RECT 2083.890 3002.400 2084.170 3002.680 ;
        RECT 2087.110 2996.280 2087.390 2996.560 ;
        RECT 2084.810 2698.440 2085.090 2698.720 ;
        RECT 2083.890 2691.640 2084.170 2691.920 ;
        RECT 2087.570 2988.120 2087.850 2988.400 ;
        RECT 2482.250 3049.320 2482.530 3049.600 ;
        RECT 2497.890 2747.400 2498.170 2747.680 ;
        RECT 2497.890 2710.000 2498.170 2710.280 ;
        RECT 2497.890 2704.560 2498.170 2704.840 ;
        RECT 2126.670 2598.480 2126.950 2598.760 ;
        RECT 2170.830 2598.480 2171.110 2598.760 ;
        RECT 2146.450 2593.040 2146.730 2593.320 ;
        RECT 2132.190 2592.360 2132.470 2592.640 ;
        RECT 2152.890 2591.680 2153.170 2591.960 ;
        RECT 2145.990 2591.000 2146.270 2591.280 ;
        RECT 2163.010 2588.960 2163.290 2589.240 ;
        RECT 2166.230 2588.280 2166.510 2588.560 ;
        RECT 2215.910 2593.720 2216.190 2594.000 ;
        RECT 2212.690 2593.040 2212.970 2593.320 ;
        RECT 2176.810 2591.680 2177.090 2591.960 ;
        RECT 2179.570 2591.680 2179.850 2591.960 ;
        RECT 2173.130 2588.280 2173.410 2588.560 ;
        RECT 2170.370 2477.440 2170.650 2477.720 ;
        RECT 2169.450 2463.160 2169.730 2463.440 ;
        RECT 2168.070 2414.880 2168.350 2415.160 ;
        RECT 2168.990 2414.880 2169.270 2415.160 ;
        RECT 2184.630 2591.000 2184.910 2591.280 ;
        RECT 2204.410 2591.000 2204.690 2591.280 ;
        RECT 2180.030 2588.280 2180.310 2588.560 ;
        RECT 2186.470 2588.960 2186.750 2589.240 ;
        RECT 2186.930 2588.280 2187.210 2588.560 ;
        RECT 2193.370 2588.280 2193.650 2588.560 ;
        RECT 2190.610 2587.600 2190.890 2587.880 ;
        RECT 2193.830 2587.600 2194.110 2587.880 ;
        RECT 2197.510 2587.600 2197.790 2587.880 ;
        RECT 2200.730 2587.600 2201.010 2587.880 ;
        RECT 2207.630 2587.600 2207.910 2587.880 ;
        RECT 2214.530 2587.600 2214.810 2587.880 ;
        RECT 2221.430 2593.040 2221.710 2593.320 ;
        RECT 2226.950 2593.040 2227.230 2593.320 ;
        RECT 2232.010 2593.040 2232.290 2593.320 ;
        RECT 2220.510 2592.360 2220.790 2592.640 ;
        RECT 2227.410 2592.360 2227.690 2592.640 ;
        RECT 2227.870 2591.680 2228.150 2591.960 ;
        RECT 2235.690 2592.360 2235.970 2592.640 ;
        RECT 2239.830 2592.360 2240.110 2592.640 ;
        RECT 2235.230 2591.680 2235.510 2591.960 ;
        RECT 2241.670 2591.000 2241.950 2591.280 ;
        RECT 2256.390 2593.720 2256.670 2594.000 ;
        RECT 2262.830 2593.720 2263.110 2594.000 ;
        RECT 2243.510 2592.360 2243.790 2592.640 ;
        RECT 2249.030 2587.600 2249.310 2587.880 ;
        RECT 2250.870 2591.680 2251.150 2591.960 ;
        RECT 2255.930 2587.600 2256.210 2587.880 ;
        RECT 2262.830 2587.600 2263.110 2587.880 ;
        RECT 2268.810 2592.360 2269.090 2592.640 ;
        RECT 2276.630 2592.360 2276.910 2592.640 ;
        RECT 2269.270 2588.280 2269.550 2588.560 ;
        RECT 2269.730 2587.600 2270.010 2587.880 ;
        RECT 2276.630 2587.600 2276.910 2587.880 ;
        RECT 2291.810 2593.720 2292.090 2594.000 ;
        RECT 2297.790 2593.720 2298.070 2594.000 ;
        RECT 2332.290 2593.720 2332.570 2594.000 ;
        RECT 2285.370 2593.040 2285.650 2593.320 ;
        RECT 2280.310 2592.360 2280.590 2592.640 ;
        RECT 2305.150 2593.040 2305.430 2593.320 ;
        RECT 2311.590 2592.360 2311.870 2592.640 ;
        RECT 2318.490 2592.360 2318.770 2592.640 ;
        RECT 2332.290 2592.360 2332.570 2592.640 ;
        RECT 2297.790 2591.680 2298.070 2591.960 ;
        RECT 2325.390 2591.680 2325.670 2591.960 ;
        RECT 2339.190 2591.000 2339.470 2591.280 ;
        RECT 2304.230 2588.280 2304.510 2588.560 ;
        RECT 2345.170 2588.280 2345.450 2588.560 ;
        RECT 2283.530 2587.600 2283.810 2587.880 ;
        RECT 2290.430 2587.600 2290.710 2587.880 ;
        RECT 2297.330 2587.600 2297.610 2587.880 ;
        RECT 2303.770 2587.600 2304.050 2587.880 ;
        RECT 2311.130 2587.600 2311.410 2587.880 ;
        RECT 2318.030 2587.600 2318.310 2587.880 ;
        RECT 2324.930 2587.600 2325.210 2587.880 ;
        RECT 2331.830 2587.600 2332.110 2587.880 ;
        RECT 2338.730 2587.600 2339.010 2587.880 ;
        RECT 2331.830 2412.160 2332.110 2412.440 ;
        RECT 2345.630 2587.600 2345.910 2587.880 ;
        RECT 2345.170 2411.480 2345.450 2411.760 ;
        RECT 2345.630 2410.800 2345.910 2411.080 ;
        RECT 2356.210 2408.760 2356.490 2409.040 ;
        RECT 2386.110 2408.760 2386.390 2409.040 ;
        RECT 2654.290 2412.160 2654.570 2412.440 ;
        RECT 2680.050 2411.480 2680.330 2411.760 ;
        RECT 2692.930 2410.800 2693.210 2411.080 ;
        RECT 1386.530 1020.880 1386.810 1021.160 ;
        RECT 1372.730 1020.200 1373.010 1020.480 ;
        RECT 1358.930 1019.520 1359.210 1019.800 ;
        RECT 1345.130 1018.840 1345.410 1019.120 ;
        RECT 1641.830 1018.160 1642.110 1018.440 ;
        RECT 1648.730 1018.160 1649.010 1018.440 ;
        RECT 1655.630 1018.160 1655.910 1018.440 ;
        RECT 1641.830 1016.800 1642.110 1017.080 ;
        RECT 1655.630 1016.120 1655.910 1016.400 ;
        RECT 1648.730 1015.440 1649.010 1015.720 ;
        RECT 1662.070 1016.800 1662.350 1017.080 ;
        RECT 1669.430 1016.800 1669.710 1017.080 ;
        RECT 1662.530 1016.120 1662.810 1016.400 ;
        RECT 1670.350 1018.160 1670.630 1018.440 ;
        RECT 1675.870 1017.480 1676.150 1017.760 ;
        RECT 1669.890 1016.120 1670.170 1016.400 ;
        RECT 1676.790 1016.120 1677.070 1016.400 ;
        RECT 1669.430 1015.440 1669.710 1015.720 ;
        RECT 1676.330 1015.440 1676.610 1015.720 ;
        RECT 1683.230 1016.800 1683.510 1017.080 ;
        RECT 1683.690 1016.120 1683.970 1016.400 ;
        RECT 1690.590 1016.800 1690.870 1017.080 ;
        RECT 1697.950 1017.480 1698.230 1017.760 ;
        RECT 1704.390 1017.480 1704.670 1017.760 ;
        RECT 1697.490 1016.120 1697.770 1016.400 ;
        RECT 1711.290 1018.160 1711.570 1018.440 ;
        RECT 1718.190 1018.160 1718.470 1018.440 ;
        RECT 1710.830 1015.440 1711.110 1015.720 ;
        RECT 1683.230 1014.760 1683.510 1015.040 ;
        RECT 1689.670 1014.760 1689.950 1015.040 ;
        RECT 1696.110 1014.760 1696.390 1015.040 ;
        RECT 1725.090 1016.120 1725.370 1016.400 ;
        RECT 1731.990 1015.440 1732.270 1015.720 ;
        RECT 1745.790 1018.160 1746.070 1018.440 ;
        RECT 1755.450 1018.160 1755.730 1018.440 ;
        RECT 1738.890 1015.440 1739.170 1015.720 ;
        RECT 1745.330 1017.480 1745.610 1017.760 ;
        RECT 1745.790 1016.120 1746.070 1016.400 ;
        RECT 1711.290 1014.760 1711.570 1015.040 ;
        RECT 1712.210 1014.760 1712.490 1015.040 ;
        RECT 1718.190 1014.760 1718.470 1015.040 ;
        RECT 1724.630 1014.760 1724.910 1015.040 ;
        RECT 1729.690 1014.760 1729.970 1015.040 ;
        RECT 1735.670 1014.760 1735.950 1015.040 ;
        RECT 1741.650 1014.760 1741.930 1015.040 ;
        RECT 1746.250 1014.760 1746.530 1015.040 ;
        RECT 1759.130 1018.160 1759.410 1018.440 ;
        RECT 1759.590 1015.440 1759.870 1015.720 ;
        RECT 1766.030 1015.440 1766.310 1015.720 ;
        RECT 1773.390 1015.440 1773.670 1015.720 ;
        RECT 1780.290 1015.440 1780.570 1015.720 ;
        RECT 1787.190 1016.800 1787.470 1017.080 ;
        RECT 1789.030 1015.440 1789.310 1015.720 ;
        RECT 1831.810 1020.880 1832.090 1021.160 ;
        RECT 1855.730 1020.880 1856.010 1021.160 ;
        RECT 1835.490 1020.200 1835.770 1020.480 ;
        RECT 1828.590 1019.520 1828.870 1019.800 ;
        RECT 1821.690 1018.840 1821.970 1019.120 ;
        RECT 1842.390 1016.120 1842.670 1016.400 ;
        RECT 1754.990 1014.760 1755.270 1015.040 ;
        RECT 1758.670 1014.760 1758.950 1015.040 ;
        RECT 1766.490 1014.760 1766.770 1015.040 ;
        RECT 1771.550 1014.760 1771.830 1015.040 ;
        RECT 1777.990 1014.760 1778.270 1015.040 ;
        RECT 1782.130 1014.760 1782.410 1015.040 ;
        RECT 1787.190 1014.760 1787.470 1015.040 ;
        RECT 1793.170 1014.760 1793.450 1015.040 ;
        RECT 1800.070 1014.760 1800.350 1015.040 ;
        RECT 1806.510 1014.760 1806.790 1015.040 ;
        RECT 1812.490 1014.760 1812.770 1015.040 ;
        RECT 1817.550 1014.760 1817.830 1015.040 ;
        RECT 1823.530 1014.760 1823.810 1015.040 ;
        RECT 1489.110 558.480 1489.390 558.760 ;
        RECT 1503.830 556.440 1504.110 556.720 ;
        RECT 1898.970 913.440 1899.250 913.720 ;
        RECT 1898.970 627.840 1899.250 628.120 ;
        RECT 1899.890 627.840 1900.170 628.120 ;
        RECT 1902.190 904.600 1902.470 904.880 ;
        RECT 1904.030 615.600 1904.310 615.880 ;
        RECT 1901.730 610.160 1902.010 610.440 ;
        RECT 1901.270 601.320 1901.550 601.600 ;
        RECT 1899.890 595.880 1900.170 596.160 ;
        RECT 1904.030 590.440 1904.310 590.720 ;
        RECT 2249.030 1020.200 2249.310 1020.480 ;
        RECT 2245.810 1016.800 2246.090 1017.080 ;
        RECT 2252.710 1016.800 2252.990 1017.080 ;
        RECT 2259.610 1016.800 2259.890 1017.080 ;
        RECT 2266.510 1016.800 2266.790 1017.080 ;
        RECT 2255.930 1016.120 2256.210 1016.400 ;
        RECT 2283.070 1020.880 2283.350 1021.160 ;
        RECT 2280.770 1016.800 2281.050 1017.080 ;
        RECT 2269.730 1016.120 2270.010 1016.400 ;
        RECT 2273.410 1016.120 2273.690 1016.400 ;
        RECT 2275.250 1016.120 2275.530 1016.400 ;
        RECT 2276.170 1016.120 2276.450 1016.400 ;
        RECT 2290.430 1016.120 2290.710 1016.400 ;
        RECT 2297.330 1016.800 2297.610 1017.080 ;
        RECT 2304.230 1016.120 2304.510 1016.400 ;
        RECT 2310.670 1016.800 2310.950 1017.080 ;
        RECT 2317.570 1016.800 2317.850 1017.080 ;
        RECT 2318.030 1016.120 2318.310 1016.400 ;
        RECT 2323.090 1016.120 2323.370 1016.400 ;
        RECT 2345.630 1020.880 2345.910 1021.160 ;
        RECT 2352.530 1020.880 2352.810 1021.160 ;
        RECT 2338.730 1020.200 2339.010 1020.480 ;
        RECT 2352.070 1020.200 2352.350 1020.480 ;
        RECT 2325.390 1016.120 2325.670 1016.400 ;
        RECT 2332.750 1016.120 2333.030 1016.400 ;
        RECT 2359.430 1016.120 2359.710 1016.400 ;
        RECT 2366.330 1016.120 2366.610 1016.400 ;
        RECT 2262.830 1014.760 2263.110 1015.040 ;
        RECT 2276.630 1014.760 2276.910 1015.040 ;
        RECT 2283.070 1014.760 2283.350 1015.040 ;
        RECT 2289.970 1014.760 2290.250 1015.040 ;
        RECT 2295.030 1014.760 2295.310 1015.040 ;
        RECT 2302.850 1014.760 2303.130 1015.040 ;
        RECT 2306.990 1014.760 2307.270 1015.040 ;
        RECT 2312.050 1014.760 2312.330 1015.040 ;
        RECT 2318.030 1014.760 2318.310 1015.040 ;
        RECT 2324.930 1014.760 2325.210 1015.040 ;
        RECT 2331.830 1014.760 2332.110 1015.040 ;
        RECT 2336.430 1014.760 2336.710 1015.040 ;
        RECT 2342.410 1014.760 2342.690 1015.040 ;
        RECT 2347.010 1014.760 2347.290 1015.040 ;
        RECT 2353.450 1014.760 2353.730 1015.040 ;
        RECT 2358.050 1014.760 2358.330 1015.040 ;
        RECT 2358.970 1014.760 2359.250 1015.040 ;
        RECT 2384.730 1038.560 2385.010 1038.840 ;
        RECT 2384.270 1020.200 2384.550 1020.480 ;
        RECT 2383.350 1019.520 2383.630 1019.800 ;
        RECT 2387.490 1020.880 2387.770 1021.160 ;
        RECT 2390.710 1020.880 2390.990 1021.160 ;
        RECT 2387.950 1020.200 2388.230 1020.480 ;
        RECT 2388.410 1019.520 2388.690 1019.800 ;
        RECT 2387.950 1016.800 2388.230 1017.080 ;
        RECT 2408.190 1020.880 2408.470 1021.160 ;
        RECT 2450.970 1020.880 2451.250 1021.160 ;
        RECT 2428.890 1020.200 2429.170 1020.480 ;
        RECT 2402.210 1019.520 2402.490 1019.800 ;
        RECT 2415.090 1018.160 2415.370 1018.440 ;
        RECT 2421.990 1017.480 2422.270 1017.760 ;
        RECT 2380.130 1016.120 2380.410 1016.400 ;
        RECT 2387.490 1016.120 2387.770 1016.400 ;
        RECT 2428.890 1016.120 2429.170 1016.400 ;
        RECT 2364.490 1014.760 2364.770 1015.040 ;
        RECT 2370.930 1014.760 2371.210 1015.040 ;
        RECT 2377.830 1014.760 2378.110 1015.040 ;
        RECT 2380.590 1014.760 2380.870 1015.040 ;
        RECT 2394.390 1014.760 2394.670 1015.040 ;
        RECT 2403.130 1014.760 2403.410 1015.040 ;
        RECT 2408.190 1014.760 2408.470 1015.040 ;
        RECT 2415.090 1014.760 2415.370 1015.040 ;
        RECT 2421.990 1014.760 2422.270 1015.040 ;
        RECT 2242.130 1007.280 2242.410 1007.560 ;
        RECT 1904.030 578.880 1904.310 579.160 ;
        RECT 1903.570 573.440 1903.850 573.720 ;
        RECT 2083.890 556.440 2084.170 556.720 ;
        RECT 2691.090 1018.840 2691.370 1019.120 ;
        RECT 2482.250 906.640 2482.530 906.920 ;
        RECT 2500.650 618.320 2500.930 618.600 ;
        RECT 2500.190 610.160 2500.470 610.440 ;
        RECT 2499.730 604.040 2500.010 604.320 ;
        RECT 2499.270 593.160 2499.550 593.440 ;
        RECT 2498.810 590.440 2499.090 590.720 ;
        RECT 2498.350 578.880 2498.630 579.160 ;
        RECT 2501.570 915.480 2501.850 915.760 ;
        RECT 2501.110 576.160 2501.390 576.440 ;
      LAYER met3 ;
        RECT 1868.125 3063.900 1868.455 3063.905 ;
        RECT 1867.870 3063.890 1868.455 3063.900 ;
        RECT 2442.665 3063.900 2442.995 3063.905 ;
        RECT 2469.805 3063.900 2470.135 3063.905 ;
        RECT 2442.665 3063.890 2443.250 3063.900 ;
        RECT 2469.550 3063.890 2470.135 3063.900 ;
        RECT 1867.870 3063.590 1868.680 3063.890 ;
        RECT 2442.665 3063.590 2443.450 3063.890 ;
        RECT 2469.350 3063.590 2470.135 3063.890 ;
        RECT 1867.870 3063.580 1868.455 3063.590 ;
        RECT 1868.125 3063.575 1868.455 3063.580 ;
        RECT 2442.665 3063.580 2443.250 3063.590 ;
        RECT 2469.550 3063.580 2470.135 3063.590 ;
        RECT 2442.665 3063.575 2442.995 3063.580 ;
        RECT 2469.805 3063.575 2470.135 3063.580 ;
        RECT 1845.790 3055.050 1846.170 3055.060 ;
        RECT 1865.110 3055.050 1865.490 3055.060 ;
        RECT 1845.790 3054.750 1865.490 3055.050 ;
        RECT 1845.790 3054.740 1846.170 3054.750 ;
        RECT 1865.110 3054.740 1865.490 3054.750 ;
        RECT 1859.280 3051.235 1861.020 3052.140 ;
        RECT 2459.280 3051.235 2461.020 3052.140 ;
        RECT 1490.005 3033.290 1490.335 3033.305 ;
        RECT 1490.005 3033.085 1497.450 3033.290 ;
        RECT 1490.005 3032.990 1504.600 3033.085 ;
        RECT 1490.005 3032.975 1490.335 3032.990 ;
        RECT 1497.150 3032.785 1504.600 3032.990 ;
        RECT 1489.545 3027.170 1489.875 3027.185 ;
        RECT 1497.150 3027.170 1504.600 3027.445 ;
        RECT 1489.545 3027.145 1504.600 3027.170 ;
        RECT 1489.545 3026.870 1497.450 3027.145 ;
        RECT 1489.545 3026.855 1489.875 3026.870 ;
        RECT 1489.085 3019.010 1489.415 3019.025 ;
        RECT 1489.085 3018.945 1497.450 3019.010 ;
        RECT 1489.085 3018.710 1504.600 3018.945 ;
        RECT 1489.085 3018.695 1489.415 3018.710 ;
        RECT 1497.150 3018.645 1504.600 3018.710 ;
        RECT 1497.150 3013.005 1504.600 3013.305 ;
        RECT 1488.625 3012.890 1488.955 3012.905 ;
        RECT 1497.150 3012.890 1497.450 3013.005 ;
        RECT 1488.625 3012.590 1497.450 3012.890 ;
        RECT 1488.625 3012.575 1488.955 3012.590 ;
        RECT 1488.165 3004.730 1488.495 3004.745 ;
        RECT 1497.150 3004.730 1504.600 3004.805 ;
        RECT 1488.165 3004.505 1504.600 3004.730 ;
        RECT 1488.165 3004.430 1497.450 3004.505 ;
        RECT 1488.165 3004.415 1488.495 3004.430 ;
        RECT 1487.705 2999.290 1488.035 2999.305 ;
        RECT 1487.705 2999.165 1497.450 2999.290 ;
        RECT 1487.705 2998.990 1504.600 2999.165 ;
        RECT 1487.705 2998.975 1488.035 2998.990 ;
        RECT 1497.150 2998.865 1504.600 2998.990 ;
        RECT 1487.245 2990.450 1487.575 2990.465 ;
        RECT 1497.150 2990.450 1504.600 2990.665 ;
        RECT 1487.245 2990.365 1504.600 2990.450 ;
        RECT 1487.245 2990.150 1497.450 2990.365 ;
        RECT 1487.245 2990.135 1487.575 2990.150 ;
        RECT 1486.785 2701.450 1487.115 2701.465 ;
        RECT 1486.785 2701.425 1497.450 2701.450 ;
        RECT 1486.785 2701.150 1504.600 2701.425 ;
        RECT 1486.785 2701.135 1487.115 2701.150 ;
        RECT 1497.150 2701.125 1504.600 2701.150 ;
        RECT 1497.150 2692.625 1504.600 2692.925 ;
        RECT 1486.325 2692.610 1486.655 2692.625 ;
        RECT 1497.150 2692.610 1497.450 2692.625 ;
        RECT 1486.325 2692.310 1497.450 2692.610 ;
        RECT 1486.325 2692.295 1486.655 2692.310 ;
      LAYER met3 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
      LAYER met3 ;
        RECT 1881.880 3048.265 1889.370 3048.565 ;
        RECT 1889.070 3048.250 1889.370 3048.265 ;
        RECT 1898.485 3048.250 1898.815 3048.265 ;
        RECT 1899.865 3048.250 1900.195 3048.265 ;
        RECT 1889.070 3047.950 1900.195 3048.250 ;
        RECT 1898.485 3047.935 1898.815 3047.950 ;
        RECT 1899.865 3047.935 1900.195 3047.950 ;
        RECT 2100.000 3032.785 2104.600 3033.085 ;
        RECT 2083.865 3030.570 2084.195 3030.585 ;
        RECT 2100.670 3030.570 2100.970 3032.785 ;
        RECT 2083.865 3030.270 2100.970 3030.570 ;
        RECT 2083.865 3030.255 2084.195 3030.270 ;
        RECT 2100.000 3027.145 2104.600 3027.445 ;
        RECT 2083.865 3024.450 2084.195 3024.465 ;
        RECT 2100.670 3024.450 2100.970 3027.145 ;
        RECT 2083.865 3024.150 2100.970 3024.450 ;
        RECT 2083.865 3024.135 2084.195 3024.150 ;
        RECT 2100.000 3018.645 2104.600 3018.945 ;
        RECT 2083.865 3016.290 2084.195 3016.305 ;
        RECT 2100.670 3016.290 2100.970 3018.645 ;
        RECT 2083.865 3015.990 2100.970 3016.290 ;
        RECT 2083.865 3015.975 2084.195 3015.990 ;
        RECT 2100.000 3013.005 2104.600 3013.305 ;
        RECT 2083.865 3010.170 2084.195 3010.185 ;
        RECT 2100.670 3010.170 2100.970 3013.005 ;
        RECT 2083.865 3009.870 2100.970 3010.170 ;
        RECT 2083.865 3009.855 2084.195 3009.870 ;
        RECT 2100.000 3004.505 2104.600 3004.805 ;
        RECT 2083.865 3002.690 2084.195 3002.705 ;
        RECT 2100.670 3002.690 2100.970 3004.505 ;
        RECT 2083.865 3002.390 2100.970 3002.690 ;
        RECT 2083.865 3002.375 2084.195 3002.390 ;
        RECT 2100.000 2998.865 2104.600 2999.165 ;
        RECT 2087.085 2996.570 2087.415 2996.585 ;
        RECT 2100.670 2996.570 2100.970 2998.865 ;
        RECT 2087.085 2996.270 2100.970 2996.570 ;
        RECT 2087.085 2996.255 2087.415 2996.270 ;
        RECT 2100.000 2990.365 2104.600 2990.665 ;
        RECT 2087.545 2988.410 2087.875 2988.425 ;
        RECT 2100.670 2988.410 2100.970 2990.365 ;
        RECT 2087.545 2988.110 2100.970 2988.410 ;
        RECT 2087.545 2988.095 2087.875 2988.110 ;
        RECT 1881.880 2747.010 1889.370 2747.210 ;
        RECT 1898.025 2747.010 1898.355 2747.025 ;
        RECT 1881.880 2746.910 1898.355 2747.010 ;
        RECT 1885.390 2738.710 1885.690 2746.910 ;
        RECT 1889.070 2746.710 1898.355 2746.910 ;
        RECT 1898.025 2746.695 1898.355 2746.710 ;
        RECT 1881.880 2738.410 1886.480 2738.710 ;
        RECT 1885.390 2733.070 1885.690 2738.410 ;
        RECT 1881.880 2732.770 1886.480 2733.070 ;
        RECT 1885.390 2724.570 1885.690 2732.770 ;
        RECT 1881.880 2724.270 1886.480 2724.570 ;
        RECT 1885.390 2718.930 1885.690 2724.270 ;
        RECT 1881.880 2718.630 1886.480 2718.930 ;
        RECT 1885.390 2710.430 1885.690 2718.630 ;
        RECT 1881.880 2710.130 1886.480 2710.430 ;
        RECT 1885.390 2704.790 1885.690 2710.130 ;
        RECT 1898.945 2704.850 1899.275 2704.865 ;
        RECT 1887.230 2704.790 1899.275 2704.850 ;
        RECT 1881.880 2704.550 1899.275 2704.790 ;
        RECT 1881.880 2704.490 1887.530 2704.550 ;
        RECT 1898.945 2704.535 1899.275 2704.550 ;
        RECT 2100.000 2701.125 2104.600 2701.425 ;
        RECT 2084.785 2698.730 2085.115 2698.745 ;
        RECT 2100.670 2698.730 2100.970 2701.125 ;
        RECT 2084.785 2698.430 2100.970 2698.730 ;
        RECT 2084.785 2698.415 2085.115 2698.430 ;
        RECT 2100.000 2692.625 2104.600 2692.925 ;
        RECT 2083.865 2691.930 2084.195 2691.945 ;
        RECT 2100.670 2691.930 2100.970 2692.625 ;
        RECT 2083.865 2691.630 2100.970 2691.930 ;
        RECT 2083.865 2691.615 2084.195 2691.630 ;
      LAYER met3 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met3 ;
        RECT 2482.225 3049.610 2482.555 3049.625 ;
        RECT 2482.225 3049.295 2482.770 3049.610 ;
        RECT 2482.470 3048.565 2482.770 3049.295 ;
        RECT 2481.880 3048.265 2486.480 3048.565 ;
        RECT 2497.865 2747.690 2498.195 2747.705 ;
        RECT 2488.910 2747.390 2498.195 2747.690 ;
        RECT 2488.910 2747.210 2489.210 2747.390 ;
        RECT 2497.865 2747.375 2498.195 2747.390 ;
        RECT 2481.880 2746.910 2489.210 2747.210 ;
        RECT 2485.230 2739.530 2485.530 2746.910 ;
        RECT 2485.230 2739.230 2486.450 2739.530 ;
        RECT 2486.150 2738.710 2486.450 2739.230 ;
        RECT 2481.880 2738.410 2486.480 2738.710 ;
        RECT 2486.150 2733.070 2486.450 2738.410 ;
        RECT 2481.880 2732.770 2486.480 2733.070 ;
        RECT 2486.150 2724.570 2486.450 2732.770 ;
        RECT 2481.880 2724.270 2486.480 2724.570 ;
        RECT 2486.150 2718.930 2486.450 2724.270 ;
        RECT 2481.880 2718.630 2486.480 2718.930 ;
        RECT 2486.150 2710.430 2486.450 2718.630 ;
        RECT 2481.880 2710.290 2486.480 2710.430 ;
        RECT 2497.865 2710.290 2498.195 2710.305 ;
        RECT 2481.880 2710.130 2498.195 2710.290 ;
        RECT 2486.150 2709.990 2498.195 2710.130 ;
        RECT 2497.865 2709.975 2498.195 2709.990 ;
        RECT 2497.865 2704.850 2498.195 2704.865 ;
        RECT 2486.150 2704.790 2498.195 2704.850 ;
        RECT 2481.880 2704.550 2498.195 2704.790 ;
        RECT 2481.880 2704.490 2486.480 2704.550 ;
        RECT 2497.865 2704.535 2498.195 2704.550 ;
        RECT 2126.645 2598.770 2126.975 2598.785 ;
        RECT 2139.810 2598.770 2140.190 2598.780 ;
        RECT 2126.645 2598.470 2140.190 2598.770 ;
        RECT 2126.645 2598.455 2126.975 2598.470 ;
        RECT 2139.810 2598.460 2140.190 2598.470 ;
        RECT 2169.010 2598.770 2169.390 2598.780 ;
        RECT 2170.805 2598.770 2171.135 2598.785 ;
        RECT 2169.010 2598.470 2171.135 2598.770 ;
        RECT 2169.010 2598.460 2169.390 2598.470 ;
        RECT 2170.805 2598.455 2171.135 2598.470 ;
        RECT 1568.870 2594.010 1569.250 2594.020 ;
        RECT 1572.805 2594.010 1573.135 2594.025 ;
        RECT 1568.870 2593.710 1573.135 2594.010 ;
        RECT 1568.870 2593.700 1569.250 2593.710 ;
        RECT 1572.805 2593.695 1573.135 2593.710 ;
        RECT 1598.310 2594.010 1598.690 2594.020 ;
        RECT 1600.405 2594.010 1600.735 2594.025 ;
        RECT 1598.310 2593.710 1600.735 2594.010 ;
        RECT 1598.310 2593.700 1598.690 2593.710 ;
        RECT 1600.405 2593.695 1600.735 2593.710 ;
        RECT 1614.665 2594.010 1614.995 2594.025 ;
        RECT 1621.565 2594.020 1621.895 2594.025 ;
        RECT 1617.630 2594.010 1618.010 2594.020 ;
        RECT 1621.310 2594.010 1621.895 2594.020 ;
        RECT 1614.665 2593.710 1618.010 2594.010 ;
        RECT 1621.110 2593.710 1621.895 2594.010 ;
        RECT 1614.665 2593.695 1614.995 2593.710 ;
        RECT 1617.630 2593.700 1618.010 2593.710 ;
        RECT 1621.310 2593.700 1621.895 2593.710 ;
        RECT 1625.910 2594.010 1626.290 2594.020 ;
        RECT 1627.085 2594.010 1627.415 2594.025 ;
        RECT 1625.910 2593.710 1627.415 2594.010 ;
        RECT 1625.910 2593.700 1626.290 2593.710 ;
        RECT 1621.565 2593.695 1621.895 2593.700 ;
        RECT 1627.085 2593.695 1627.415 2593.710 ;
        RECT 1632.145 2594.020 1632.475 2594.025 ;
        RECT 1636.745 2594.020 1637.075 2594.025 ;
        RECT 1644.565 2594.020 1644.895 2594.025 ;
        RECT 1632.145 2594.010 1632.730 2594.020 ;
        RECT 1636.745 2594.010 1637.330 2594.020 ;
        RECT 1644.310 2594.010 1644.895 2594.020 ;
        RECT 1632.145 2593.710 1632.930 2594.010 ;
        RECT 1636.745 2593.710 1637.530 2594.010 ;
        RECT 1644.110 2593.710 1644.895 2594.010 ;
        RECT 1632.145 2593.700 1632.730 2593.710 ;
        RECT 1636.745 2593.700 1637.330 2593.710 ;
        RECT 1644.310 2593.700 1644.895 2593.710 ;
        RECT 1632.145 2593.695 1632.475 2593.700 ;
        RECT 1636.745 2593.695 1637.075 2593.700 ;
        RECT 1644.565 2593.695 1644.895 2593.700 ;
        RECT 1650.545 2594.020 1650.875 2594.025 ;
        RECT 1650.545 2594.010 1651.130 2594.020 ;
        RECT 1656.525 2594.010 1656.855 2594.025 ;
        RECT 1662.045 2594.020 1662.375 2594.025 ;
        RECT 1658.110 2594.010 1658.490 2594.020 ;
        RECT 1661.790 2594.010 1662.375 2594.020 ;
        RECT 1650.545 2593.710 1651.330 2594.010 ;
        RECT 1656.525 2593.710 1658.490 2594.010 ;
        RECT 1661.590 2593.710 1662.375 2594.010 ;
        RECT 1650.545 2593.700 1651.130 2593.710 ;
        RECT 1650.545 2593.695 1650.875 2593.700 ;
        RECT 1656.525 2593.695 1656.855 2593.710 ;
        RECT 1658.110 2593.700 1658.490 2593.710 ;
        RECT 1661.790 2593.700 1662.375 2593.710 ;
        RECT 1668.230 2594.010 1668.610 2594.020 ;
        RECT 1668.945 2594.010 1669.275 2594.025 ;
        RECT 1668.230 2593.710 1669.275 2594.010 ;
        RECT 1668.230 2593.700 1668.610 2593.710 ;
        RECT 1662.045 2593.695 1662.375 2593.700 ;
        RECT 1668.945 2593.695 1669.275 2593.710 ;
        RECT 1672.830 2594.010 1673.210 2594.020 ;
        RECT 1673.545 2594.010 1673.875 2594.025 ;
        RECT 1672.830 2593.710 1673.875 2594.010 ;
        RECT 1672.830 2593.700 1673.210 2593.710 ;
        RECT 1673.545 2593.695 1673.875 2593.710 ;
        RECT 1679.065 2594.020 1679.395 2594.025 ;
        RECT 1684.585 2594.020 1684.915 2594.025 ;
        RECT 1690.565 2594.020 1690.895 2594.025 ;
        RECT 1679.065 2594.010 1679.650 2594.020 ;
        RECT 1684.585 2594.010 1685.170 2594.020 ;
        RECT 1690.310 2594.010 1690.895 2594.020 ;
        RECT 1679.065 2593.710 1679.850 2594.010 ;
        RECT 1684.585 2593.710 1685.370 2594.010 ;
        RECT 1690.110 2593.710 1690.895 2594.010 ;
        RECT 1679.065 2593.700 1679.650 2593.710 ;
        RECT 1684.585 2593.700 1685.170 2593.710 ;
        RECT 1690.310 2593.700 1690.895 2593.710 ;
        RECT 1679.065 2593.695 1679.395 2593.700 ;
        RECT 1684.585 2593.695 1684.915 2593.700 ;
        RECT 1690.565 2593.695 1690.895 2593.700 ;
        RECT 1697.465 2594.020 1697.795 2594.025 ;
        RECT 1697.465 2594.010 1698.050 2594.020 ;
        RECT 1702.270 2594.010 1702.650 2594.020 ;
        RECT 1702.985 2594.010 1703.315 2594.025 ;
        RECT 1697.465 2593.710 1698.250 2594.010 ;
        RECT 1702.270 2593.710 1703.315 2594.010 ;
        RECT 1697.465 2593.700 1698.050 2593.710 ;
        RECT 1702.270 2593.700 1702.650 2593.710 ;
        RECT 1697.465 2593.695 1697.795 2593.700 ;
        RECT 1702.985 2593.695 1703.315 2593.710 ;
        RECT 1707.585 2594.020 1707.915 2594.025 ;
        RECT 1707.585 2594.010 1708.170 2594.020 ;
        RECT 1725.270 2594.010 1725.650 2594.020 ;
        RECT 1726.445 2594.010 1726.775 2594.025 ;
        RECT 1732.885 2594.020 1733.215 2594.025 ;
        RECT 1744.845 2594.020 1745.175 2594.025 ;
        RECT 2215.885 2594.020 2216.215 2594.025 ;
        RECT 2256.365 2594.020 2256.695 2594.025 ;
        RECT 2262.805 2594.020 2263.135 2594.025 ;
        RECT 1732.630 2594.010 1733.215 2594.020 ;
        RECT 1744.590 2594.010 1745.175 2594.020 ;
        RECT 2215.630 2594.010 2216.215 2594.020 ;
        RECT 1707.585 2593.710 1708.370 2594.010 ;
        RECT 1725.270 2593.710 1726.775 2594.010 ;
        RECT 1732.430 2593.710 1733.215 2594.010 ;
        RECT 1744.390 2593.710 1745.175 2594.010 ;
        RECT 2215.430 2593.710 2216.215 2594.010 ;
        RECT 1707.585 2593.700 1708.170 2593.710 ;
        RECT 1725.270 2593.700 1725.650 2593.710 ;
        RECT 1707.585 2593.695 1707.915 2593.700 ;
        RECT 1726.445 2593.695 1726.775 2593.710 ;
        RECT 1732.630 2593.700 1733.215 2593.710 ;
        RECT 1744.590 2593.700 1745.175 2593.710 ;
        RECT 2215.630 2593.700 2216.215 2593.710 ;
        RECT 2256.110 2594.010 2256.695 2594.020 ;
        RECT 2262.550 2594.010 2263.135 2594.020 ;
        RECT 2256.110 2593.710 2256.920 2594.010 ;
        RECT 2262.350 2593.710 2263.135 2594.010 ;
        RECT 2256.110 2593.700 2256.695 2593.710 ;
        RECT 2262.550 2593.700 2263.135 2593.710 ;
        RECT 1732.885 2593.695 1733.215 2593.700 ;
        RECT 1744.845 2593.695 1745.175 2593.700 ;
        RECT 2215.885 2593.695 2216.215 2593.700 ;
        RECT 2256.365 2593.695 2256.695 2593.700 ;
        RECT 2262.805 2593.695 2263.135 2593.700 ;
        RECT 2291.785 2594.020 2292.115 2594.025 ;
        RECT 2291.785 2594.010 2292.370 2594.020 ;
        RECT 2297.765 2594.010 2298.095 2594.025 ;
        RECT 2332.265 2594.020 2332.595 2594.025 ;
        RECT 2302.110 2594.010 2302.490 2594.020 ;
        RECT 2332.265 2594.010 2332.850 2594.020 ;
        RECT 2291.785 2593.710 2292.570 2594.010 ;
        RECT 2297.765 2593.710 2302.490 2594.010 ;
        RECT 2332.040 2593.710 2332.850 2594.010 ;
        RECT 2291.785 2593.700 2292.370 2593.710 ;
        RECT 2291.785 2593.695 2292.115 2593.700 ;
        RECT 2297.765 2593.695 2298.095 2593.710 ;
        RECT 2302.110 2593.700 2302.490 2593.710 ;
        RECT 2332.265 2593.700 2332.850 2593.710 ;
        RECT 2332.265 2593.695 2332.595 2593.700 ;
        RECT 1562.430 2593.330 1562.810 2593.340 ;
        RECT 1565.905 2593.330 1566.235 2593.345 ;
        RECT 1562.430 2593.030 1566.235 2593.330 ;
        RECT 1562.430 2593.020 1562.810 2593.030 ;
        RECT 1565.905 2593.015 1566.235 2593.030 ;
        RECT 1580.830 2593.330 1581.210 2593.340 ;
        RECT 1586.145 2593.330 1586.475 2593.345 ;
        RECT 1580.830 2593.030 1586.475 2593.330 ;
        RECT 1580.830 2593.020 1581.210 2593.030 ;
        RECT 1586.145 2593.015 1586.475 2593.030 ;
        RECT 1592.790 2593.330 1593.170 2593.340 ;
        RECT 1593.505 2593.330 1593.835 2593.345 ;
        RECT 1592.790 2593.030 1593.835 2593.330 ;
        RECT 1592.790 2593.020 1593.170 2593.030 ;
        RECT 1593.505 2593.015 1593.835 2593.030 ;
        RECT 1603.830 2593.330 1604.210 2593.340 ;
        RECT 1605.465 2593.330 1605.795 2593.345 ;
        RECT 1603.830 2593.030 1605.795 2593.330 ;
        RECT 1603.830 2593.020 1604.210 2593.030 ;
        RECT 1605.465 2593.015 1605.795 2593.030 ;
        RECT 1615.585 2593.340 1615.915 2593.345 ;
        RECT 1615.585 2593.330 1616.170 2593.340 ;
        RECT 1656.270 2593.330 1656.650 2593.340 ;
        RECT 1656.985 2593.330 1657.315 2593.345 ;
        RECT 1615.585 2593.030 1616.370 2593.330 ;
        RECT 1656.270 2593.030 1657.315 2593.330 ;
        RECT 1615.585 2593.020 1616.170 2593.030 ;
        RECT 1656.270 2593.020 1656.650 2593.030 ;
        RECT 1615.585 2593.015 1615.915 2593.020 ;
        RECT 1656.985 2593.015 1657.315 2593.030 ;
        RECT 1697.925 2593.330 1698.255 2593.345 ;
        RECT 1738.405 2593.340 1738.735 2593.345 ;
        RECT 1703.190 2593.330 1703.570 2593.340 ;
        RECT 1738.150 2593.330 1738.735 2593.340 ;
        RECT 1697.925 2593.030 1703.570 2593.330 ;
        RECT 1737.950 2593.030 1738.735 2593.330 ;
        RECT 1697.925 2593.015 1698.255 2593.030 ;
        RECT 1703.190 2593.020 1703.570 2593.030 ;
        RECT 1738.150 2593.020 1738.735 2593.030 ;
        RECT 1738.405 2593.015 1738.735 2593.020 ;
        RECT 2146.425 2593.330 2146.755 2593.345 ;
        RECT 2148.470 2593.330 2148.850 2593.340 ;
        RECT 2146.425 2593.030 2148.850 2593.330 ;
        RECT 2146.425 2593.015 2146.755 2593.030 ;
        RECT 2148.470 2593.020 2148.850 2593.030 ;
        RECT 2208.270 2593.330 2208.650 2593.340 ;
        RECT 2212.665 2593.330 2212.995 2593.345 ;
        RECT 2208.270 2593.030 2212.995 2593.330 ;
        RECT 2208.270 2593.020 2208.650 2593.030 ;
        RECT 2212.665 2593.015 2212.995 2593.030 ;
        RECT 2220.230 2593.330 2220.610 2593.340 ;
        RECT 2221.405 2593.330 2221.735 2593.345 ;
        RECT 2226.925 2593.340 2227.255 2593.345 ;
        RECT 2226.670 2593.330 2227.255 2593.340 ;
        RECT 2220.230 2593.030 2221.735 2593.330 ;
        RECT 2226.470 2593.030 2227.255 2593.330 ;
        RECT 2220.230 2593.020 2220.610 2593.030 ;
        RECT 2221.405 2593.015 2221.735 2593.030 ;
        RECT 2226.670 2593.020 2227.255 2593.030 ;
        RECT 2226.925 2593.015 2227.255 2593.020 ;
        RECT 2231.985 2593.330 2232.315 2593.345 ;
        RECT 2285.345 2593.340 2285.675 2593.345 ;
        RECT 2233.110 2593.330 2233.490 2593.340 ;
        RECT 2231.985 2593.030 2233.490 2593.330 ;
        RECT 2231.985 2593.015 2232.315 2593.030 ;
        RECT 2233.110 2593.020 2233.490 2593.030 ;
        RECT 2285.345 2593.330 2285.930 2593.340 ;
        RECT 2305.125 2593.330 2305.455 2593.345 ;
        RECT 2305.790 2593.330 2306.170 2593.340 ;
        RECT 2285.345 2593.030 2286.130 2593.330 ;
        RECT 2305.125 2593.030 2306.170 2593.330 ;
        RECT 2285.345 2593.020 2285.930 2593.030 ;
        RECT 2285.345 2593.015 2285.675 2593.020 ;
        RECT 2305.125 2593.015 2305.455 2593.030 ;
        RECT 2305.790 2593.020 2306.170 2593.030 ;
        RECT 1573.265 2592.650 1573.595 2592.665 ;
        RECT 1575.310 2592.650 1575.690 2592.660 ;
        RECT 1573.265 2592.350 1575.690 2592.650 ;
        RECT 1573.265 2592.335 1573.595 2592.350 ;
        RECT 1575.310 2592.340 1575.690 2592.350 ;
        RECT 1580.165 2592.650 1580.495 2592.665 ;
        RECT 1586.605 2592.660 1586.935 2592.665 ;
        RECT 1582.670 2592.650 1583.050 2592.660 ;
        RECT 1580.165 2592.350 1583.050 2592.650 ;
        RECT 1580.165 2592.335 1580.495 2592.350 ;
        RECT 1582.670 2592.340 1583.050 2592.350 ;
        RECT 1586.350 2592.650 1586.935 2592.660 ;
        RECT 1587.525 2592.650 1587.855 2592.665 ;
        RECT 1592.790 2592.650 1593.170 2592.660 ;
        RECT 1608.430 2592.650 1608.810 2592.660 ;
        RECT 1627.545 2592.650 1627.875 2592.665 ;
        RECT 1586.350 2592.350 1587.160 2592.650 ;
        RECT 1587.525 2592.350 1593.170 2592.650 ;
        RECT 1586.350 2592.340 1586.935 2592.350 ;
        RECT 1586.605 2592.335 1586.935 2592.340 ;
        RECT 1587.525 2592.335 1587.855 2592.350 ;
        RECT 1592.790 2592.340 1593.170 2592.350 ;
        RECT 1593.980 2592.350 1627.875 2592.650 ;
        RECT 1593.980 2591.985 1594.280 2592.350 ;
        RECT 1608.430 2592.340 1608.810 2592.350 ;
        RECT 1627.545 2592.335 1627.875 2592.350 ;
        RECT 1649.165 2592.650 1649.495 2592.665 ;
        RECT 1714.945 2592.660 1715.275 2592.665 ;
        RECT 1651.670 2592.650 1652.050 2592.660 ;
        RECT 1649.165 2592.350 1652.050 2592.650 ;
        RECT 1649.165 2592.335 1649.495 2592.350 ;
        RECT 1651.670 2592.340 1652.050 2592.350 ;
        RECT 1714.945 2592.650 1715.530 2592.660 ;
        RECT 1738.865 2592.650 1739.195 2592.665 ;
        RECT 1744.590 2592.650 1744.970 2592.660 ;
        RECT 1714.945 2592.350 1715.730 2592.650 ;
        RECT 1738.865 2592.350 1744.970 2592.650 ;
        RECT 1714.945 2592.340 1715.530 2592.350 ;
        RECT 1714.945 2592.335 1715.275 2592.340 ;
        RECT 1738.865 2592.335 1739.195 2592.350 ;
        RECT 1744.590 2592.340 1744.970 2592.350 ;
        RECT 2132.165 2592.650 2132.495 2592.665 ;
        RECT 2132.830 2592.650 2133.210 2592.660 ;
        RECT 2132.165 2592.350 2133.210 2592.650 ;
        RECT 2132.165 2592.335 2132.495 2592.350 ;
        RECT 2132.830 2592.340 2133.210 2592.350 ;
        RECT 2219.310 2592.650 2219.690 2592.660 ;
        RECT 2220.485 2592.650 2220.815 2592.665 ;
        RECT 2219.310 2592.350 2220.815 2592.650 ;
        RECT 2219.310 2592.340 2219.690 2592.350 ;
        RECT 2220.485 2592.335 2220.815 2592.350 ;
        RECT 2224.830 2592.650 2225.210 2592.660 ;
        RECT 2227.385 2592.650 2227.715 2592.665 ;
        RECT 2224.830 2592.350 2227.715 2592.650 ;
        RECT 2224.830 2592.340 2225.210 2592.350 ;
        RECT 2227.385 2592.335 2227.715 2592.350 ;
        RECT 2235.665 2592.650 2235.995 2592.665 ;
        RECT 2238.630 2592.650 2239.010 2592.660 ;
        RECT 2239.805 2592.650 2240.135 2592.665 ;
        RECT 2235.665 2592.350 2240.135 2592.650 ;
        RECT 2235.665 2592.335 2235.995 2592.350 ;
        RECT 2238.630 2592.340 2239.010 2592.350 ;
        RECT 2239.805 2592.335 2240.135 2592.350 ;
        RECT 2243.485 2592.650 2243.815 2592.665 ;
        RECT 2244.150 2592.650 2244.530 2592.660 ;
        RECT 2243.485 2592.350 2244.530 2592.650 ;
        RECT 2243.485 2592.335 2243.815 2592.350 ;
        RECT 2244.150 2592.340 2244.530 2592.350 ;
        RECT 2268.070 2592.650 2268.450 2592.660 ;
        RECT 2268.785 2592.650 2269.115 2592.665 ;
        RECT 2268.070 2592.350 2269.115 2592.650 ;
        RECT 2268.070 2592.340 2268.450 2592.350 ;
        RECT 2268.785 2592.335 2269.115 2592.350 ;
        RECT 2273.590 2592.650 2273.970 2592.660 ;
        RECT 2276.605 2592.650 2276.935 2592.665 ;
        RECT 2280.285 2592.660 2280.615 2592.665 ;
        RECT 2280.030 2592.650 2280.615 2592.660 ;
        RECT 2273.590 2592.350 2276.935 2592.650 ;
        RECT 2279.830 2592.350 2280.615 2592.650 ;
        RECT 2273.590 2592.340 2273.970 2592.350 ;
        RECT 2276.605 2592.335 2276.935 2592.350 ;
        RECT 2280.030 2592.340 2280.615 2592.350 ;
        RECT 2280.285 2592.335 2280.615 2592.340 ;
        RECT 2311.565 2592.650 2311.895 2592.665 ;
        RECT 2312.230 2592.650 2312.610 2592.660 ;
        RECT 2311.565 2592.350 2312.610 2592.650 ;
        RECT 2311.565 2592.335 2311.895 2592.350 ;
        RECT 2312.230 2592.340 2312.610 2592.350 ;
        RECT 2318.465 2592.650 2318.795 2592.665 ;
        RECT 2319.590 2592.650 2319.970 2592.660 ;
        RECT 2318.465 2592.350 2319.970 2592.650 ;
        RECT 2318.465 2592.335 2318.795 2592.350 ;
        RECT 2319.590 2592.340 2319.970 2592.350 ;
        RECT 2332.265 2592.650 2332.595 2592.665 ;
        RECT 2337.070 2592.650 2337.450 2592.660 ;
        RECT 2332.265 2592.350 2337.450 2592.650 ;
        RECT 2332.265 2592.335 2332.595 2592.350 ;
        RECT 2337.070 2592.340 2337.450 2592.350 ;
        RECT 1566.365 2591.970 1566.695 2591.985 ;
        RECT 1569.790 2591.970 1570.170 2591.980 ;
        RECT 1566.365 2591.670 1570.170 2591.970 ;
        RECT 1566.365 2591.655 1566.695 2591.670 ;
        RECT 1569.790 2591.660 1570.170 2591.670 ;
        RECT 1593.965 2591.655 1594.295 2591.985 ;
        RECT 1600.865 2591.970 1601.195 2591.985 ;
        RECT 1604.750 2591.970 1605.130 2591.980 ;
        RECT 1600.865 2591.670 1605.130 2591.970 ;
        RECT 1600.865 2591.655 1601.195 2591.670 ;
        RECT 1604.750 2591.660 1605.130 2591.670 ;
        RECT 1683.665 2591.970 1683.995 2591.985 ;
        RECT 1686.630 2591.970 1687.010 2591.980 ;
        RECT 1683.665 2591.670 1687.010 2591.970 ;
        RECT 1683.665 2591.655 1683.995 2591.670 ;
        RECT 1686.630 2591.660 1687.010 2591.670 ;
        RECT 1690.565 2591.970 1690.895 2591.985 ;
        RECT 1692.150 2591.970 1692.530 2591.980 ;
        RECT 1690.565 2591.670 1692.530 2591.970 ;
        RECT 1690.565 2591.655 1690.895 2591.670 ;
        RECT 1692.150 2591.660 1692.530 2591.670 ;
        RECT 1697.465 2591.970 1697.795 2591.985 ;
        RECT 1718.625 2591.980 1718.955 2591.985 ;
        RECT 1699.510 2591.970 1699.890 2591.980 ;
        RECT 1697.465 2591.670 1699.890 2591.970 ;
        RECT 1697.465 2591.655 1697.795 2591.670 ;
        RECT 1699.510 2591.660 1699.890 2591.670 ;
        RECT 1718.625 2591.970 1719.210 2591.980 ;
        RECT 2152.865 2591.970 2153.195 2591.985 ;
        RECT 2153.990 2591.970 2154.370 2591.980 ;
        RECT 1718.625 2591.670 1719.410 2591.970 ;
        RECT 2152.865 2591.670 2154.370 2591.970 ;
        RECT 1718.625 2591.660 1719.210 2591.670 ;
        RECT 1718.625 2591.655 1718.955 2591.660 ;
        RECT 2152.865 2591.655 2153.195 2591.670 ;
        RECT 2153.990 2591.660 2154.370 2591.670 ;
        RECT 2175.150 2591.970 2175.530 2591.980 ;
        RECT 2176.785 2591.970 2177.115 2591.985 ;
        RECT 2179.545 2591.970 2179.875 2591.985 ;
        RECT 2227.845 2591.980 2228.175 2591.985 ;
        RECT 2235.205 2591.980 2235.535 2591.985 ;
        RECT 2250.845 2591.980 2251.175 2591.985 ;
        RECT 2297.765 2591.980 2298.095 2591.985 ;
        RECT 2227.590 2591.970 2228.175 2591.980 ;
        RECT 2234.950 2591.970 2235.535 2591.980 ;
        RECT 2250.590 2591.970 2251.175 2591.980 ;
        RECT 2297.510 2591.970 2298.095 2591.980 ;
        RECT 2175.150 2591.670 2179.875 2591.970 ;
        RECT 2227.390 2591.670 2228.175 2591.970 ;
        RECT 2234.750 2591.670 2235.535 2591.970 ;
        RECT 2250.390 2591.670 2251.175 2591.970 ;
        RECT 2297.310 2591.670 2298.095 2591.970 ;
        RECT 2175.150 2591.660 2175.530 2591.670 ;
        RECT 2176.785 2591.655 2177.115 2591.670 ;
        RECT 2179.545 2591.655 2179.875 2591.670 ;
        RECT 2227.590 2591.660 2228.175 2591.670 ;
        RECT 2234.950 2591.660 2235.535 2591.670 ;
        RECT 2250.590 2591.660 2251.175 2591.670 ;
        RECT 2297.510 2591.660 2298.095 2591.670 ;
        RECT 2227.845 2591.655 2228.175 2591.660 ;
        RECT 2235.205 2591.655 2235.535 2591.660 ;
        RECT 2250.845 2591.655 2251.175 2591.660 ;
        RECT 2297.765 2591.655 2298.095 2591.660 ;
        RECT 2325.365 2591.970 2325.695 2591.985 ;
        RECT 2326.030 2591.970 2326.410 2591.980 ;
        RECT 2325.365 2591.670 2326.410 2591.970 ;
        RECT 2325.365 2591.655 2325.695 2591.670 ;
        RECT 2326.030 2591.660 2326.410 2591.670 ;
        RECT 1608.685 2591.290 1609.015 2591.305 ;
        RECT 1610.270 2591.290 1610.650 2591.300 ;
        RECT 1608.685 2590.990 1610.650 2591.290 ;
        RECT 1608.685 2590.975 1609.015 2590.990 ;
        RECT 1610.270 2590.980 1610.650 2590.990 ;
        RECT 1663.425 2591.290 1663.755 2591.305 ;
        RECT 1669.150 2591.290 1669.530 2591.300 ;
        RECT 1663.425 2590.990 1669.530 2591.290 ;
        RECT 1663.425 2590.975 1663.755 2590.990 ;
        RECT 1669.150 2590.980 1669.530 2590.990 ;
        RECT 1704.365 2591.290 1704.695 2591.305 ;
        RECT 2145.965 2591.300 2146.295 2591.305 ;
        RECT 1709.630 2591.290 1710.010 2591.300 ;
        RECT 1704.365 2590.990 1710.010 2591.290 ;
        RECT 1704.365 2590.975 1704.695 2590.990 ;
        RECT 1709.630 2590.980 1710.010 2590.990 ;
        RECT 2145.710 2591.290 2146.295 2591.300 ;
        RECT 2180.670 2591.290 2181.050 2591.300 ;
        RECT 2184.605 2591.290 2184.935 2591.305 ;
        RECT 2145.710 2590.990 2146.520 2591.290 ;
        RECT 2180.670 2590.990 2184.935 2591.290 ;
        RECT 2145.710 2590.980 2146.295 2590.990 ;
        RECT 2180.670 2590.980 2181.050 2590.990 ;
        RECT 2145.965 2590.975 2146.295 2590.980 ;
        RECT 2184.605 2590.975 2184.935 2590.990 ;
        RECT 2203.670 2591.290 2204.050 2591.300 ;
        RECT 2204.385 2591.290 2204.715 2591.305 ;
        RECT 2241.645 2591.300 2241.975 2591.305 ;
        RECT 2241.390 2591.290 2241.975 2591.300 ;
        RECT 2203.670 2590.990 2204.715 2591.290 ;
        RECT 2241.190 2590.990 2241.975 2591.290 ;
        RECT 2203.670 2590.980 2204.050 2590.990 ;
        RECT 2204.385 2590.975 2204.715 2590.990 ;
        RECT 2241.390 2590.980 2241.975 2590.990 ;
        RECT 2241.645 2590.975 2241.975 2590.980 ;
        RECT 2339.165 2591.290 2339.495 2591.305 ;
        RECT 2342.590 2591.290 2342.970 2591.300 ;
        RECT 2339.165 2590.990 2342.970 2591.290 ;
        RECT 2339.165 2590.975 2339.495 2590.990 ;
        RECT 2342.590 2590.980 2342.970 2590.990 ;
        RECT 1573.470 2590.610 1573.850 2590.620 ;
        RECT 1579.705 2590.610 1580.035 2590.625 ;
        RECT 1573.470 2590.310 1580.035 2590.610 ;
        RECT 1573.470 2590.300 1573.850 2590.310 ;
        RECT 1579.705 2590.295 1580.035 2590.310 ;
        RECT 1593.965 2590.610 1594.295 2590.625 ;
        RECT 1600.150 2590.610 1600.530 2590.620 ;
        RECT 1593.965 2590.310 1600.530 2590.610 ;
        RECT 1593.965 2590.295 1594.295 2590.310 ;
        RECT 1600.150 2590.300 1600.530 2590.310 ;
        RECT 1587.065 2589.940 1587.395 2589.945 ;
        RECT 1587.065 2589.930 1587.650 2589.940 ;
        RECT 1586.840 2589.630 1587.650 2589.930 ;
        RECT 1587.065 2589.620 1587.650 2589.630 ;
        RECT 1587.065 2589.615 1587.395 2589.620 ;
        RECT 1560.845 2589.250 1561.175 2589.265 ;
        RECT 1563.350 2589.250 1563.730 2589.260 ;
        RECT 1560.845 2588.950 1563.730 2589.250 ;
        RECT 1560.845 2588.935 1561.175 2588.950 ;
        RECT 1563.350 2588.940 1563.730 2588.950 ;
        RECT 1669.865 2589.250 1670.195 2589.265 ;
        RECT 1674.670 2589.250 1675.050 2589.260 ;
        RECT 1669.865 2588.950 1675.050 2589.250 ;
        RECT 1669.865 2588.935 1670.195 2588.950 ;
        RECT 1674.670 2588.940 1675.050 2588.950 ;
        RECT 1711.265 2589.250 1711.595 2589.265 ;
        RECT 1739.325 2589.260 1739.655 2589.265 ;
        RECT 1716.990 2589.250 1717.370 2589.260 ;
        RECT 1711.265 2588.950 1717.370 2589.250 ;
        RECT 1711.265 2588.935 1711.595 2588.950 ;
        RECT 1716.990 2588.940 1717.370 2588.950 ;
        RECT 1739.070 2589.250 1739.655 2589.260 ;
        RECT 2162.985 2589.260 2163.315 2589.265 ;
        RECT 2186.445 2589.260 2186.775 2589.265 ;
        RECT 2162.985 2589.250 2163.570 2589.260 ;
        RECT 1739.070 2588.950 1739.880 2589.250 ;
        RECT 2162.760 2588.950 2163.570 2589.250 ;
        RECT 1739.070 2588.940 1739.655 2588.950 ;
        RECT 1739.325 2588.935 1739.655 2588.940 ;
        RECT 2162.985 2588.940 2163.570 2588.950 ;
        RECT 2186.190 2589.250 2186.775 2589.260 ;
        RECT 2186.190 2588.950 2187.000 2589.250 ;
        RECT 2186.190 2588.940 2186.775 2588.950 ;
        RECT 2162.985 2588.935 2163.315 2588.940 ;
        RECT 2186.445 2588.935 2186.775 2588.940 ;
        RECT 1548.630 2588.570 1549.010 2588.580 ;
        RECT 1551.185 2588.570 1551.515 2588.585 ;
        RECT 1622.485 2588.580 1622.815 2588.585 ;
        RECT 1548.630 2588.270 1551.515 2588.570 ;
        RECT 1548.630 2588.260 1549.010 2588.270 ;
        RECT 1551.185 2588.255 1551.515 2588.270 ;
        RECT 1622.230 2588.570 1622.815 2588.580 ;
        RECT 1628.465 2588.570 1628.795 2588.585 ;
        RECT 1633.270 2588.570 1633.650 2588.580 ;
        RECT 1622.230 2588.270 1623.040 2588.570 ;
        RECT 1628.465 2588.270 1633.650 2588.570 ;
        RECT 1622.230 2588.260 1622.815 2588.270 ;
        RECT 1622.485 2588.255 1622.815 2588.260 ;
        RECT 1628.465 2588.255 1628.795 2588.270 ;
        RECT 1633.270 2588.260 1633.650 2588.270 ;
        RECT 1635.825 2588.570 1636.155 2588.585 ;
        RECT 1639.710 2588.570 1640.090 2588.580 ;
        RECT 1635.825 2588.270 1640.090 2588.570 ;
        RECT 1635.825 2588.255 1636.155 2588.270 ;
        RECT 1639.710 2588.260 1640.090 2588.270 ;
        RECT 1642.265 2588.570 1642.595 2588.585 ;
        RECT 1662.965 2588.580 1663.295 2588.585 ;
        RECT 1645.230 2588.570 1645.610 2588.580 ;
        RECT 1642.265 2588.270 1645.610 2588.570 ;
        RECT 1642.265 2588.255 1642.595 2588.270 ;
        RECT 1645.230 2588.260 1645.610 2588.270 ;
        RECT 1662.710 2588.570 1663.295 2588.580 ;
        RECT 1676.765 2588.570 1677.095 2588.585 ;
        RECT 1680.190 2588.570 1680.570 2588.580 ;
        RECT 1662.710 2588.270 1663.520 2588.570 ;
        RECT 1676.765 2588.270 1680.570 2588.570 ;
        RECT 1662.710 2588.260 1663.295 2588.270 ;
        RECT 1662.965 2588.255 1663.295 2588.260 ;
        RECT 1676.765 2588.255 1677.095 2588.270 ;
        RECT 1680.190 2588.260 1680.570 2588.270 ;
        RECT 1718.165 2588.570 1718.495 2588.585 ;
        RECT 1721.590 2588.570 1721.970 2588.580 ;
        RECT 1718.165 2588.270 1721.970 2588.570 ;
        RECT 1718.165 2588.255 1718.495 2588.270 ;
        RECT 1721.590 2588.260 1721.970 2588.270 ;
        RECT 1725.985 2588.570 1726.315 2588.585 ;
        RECT 1727.110 2588.570 1727.490 2588.580 ;
        RECT 1725.985 2588.270 1727.490 2588.570 ;
        RECT 1725.985 2588.255 1726.315 2588.270 ;
        RECT 1727.110 2588.260 1727.490 2588.270 ;
        RECT 1731.965 2588.570 1732.295 2588.585 ;
        RECT 1733.550 2588.570 1733.930 2588.580 ;
        RECT 1731.965 2588.270 1733.930 2588.570 ;
        RECT 1731.965 2588.255 1732.295 2588.270 ;
        RECT 1733.550 2588.260 1733.930 2588.270 ;
        RECT 2165.030 2588.570 2165.410 2588.580 ;
        RECT 2166.205 2588.570 2166.535 2588.585 ;
        RECT 2165.030 2588.270 2166.535 2588.570 ;
        RECT 2165.030 2588.260 2165.410 2588.270 ;
        RECT 2166.205 2588.255 2166.535 2588.270 ;
        RECT 2169.630 2588.570 2170.010 2588.580 ;
        RECT 2173.105 2588.570 2173.435 2588.585 ;
        RECT 2169.630 2588.270 2173.435 2588.570 ;
        RECT 2169.630 2588.260 2170.010 2588.270 ;
        RECT 2173.105 2588.255 2173.435 2588.270 ;
        RECT 2178.830 2588.570 2179.210 2588.580 ;
        RECT 2180.005 2588.570 2180.335 2588.585 ;
        RECT 2178.830 2588.270 2180.335 2588.570 ;
        RECT 2178.830 2588.260 2179.210 2588.270 ;
        RECT 2180.005 2588.255 2180.335 2588.270 ;
        RECT 2184.350 2588.570 2184.730 2588.580 ;
        RECT 2186.905 2588.570 2187.235 2588.585 ;
        RECT 2184.350 2588.270 2187.235 2588.570 ;
        RECT 2184.350 2588.260 2184.730 2588.270 ;
        RECT 2186.905 2588.255 2187.235 2588.270 ;
        RECT 2189.870 2588.570 2190.250 2588.580 ;
        RECT 2193.345 2588.570 2193.675 2588.585 ;
        RECT 2189.870 2588.270 2193.675 2588.570 ;
        RECT 2189.870 2588.260 2190.250 2588.270 ;
        RECT 2193.345 2588.255 2193.675 2588.270 ;
        RECT 2266.230 2588.570 2266.610 2588.580 ;
        RECT 2269.245 2588.570 2269.575 2588.585 ;
        RECT 2266.230 2588.270 2269.575 2588.570 ;
        RECT 2266.230 2588.260 2266.610 2588.270 ;
        RECT 2269.245 2588.255 2269.575 2588.270 ;
        RECT 2301.190 2588.570 2301.570 2588.580 ;
        RECT 2304.205 2588.570 2304.535 2588.585 ;
        RECT 2301.190 2588.270 2304.535 2588.570 ;
        RECT 2301.190 2588.260 2301.570 2588.270 ;
        RECT 2304.205 2588.255 2304.535 2588.270 ;
        RECT 2341.670 2588.570 2342.050 2588.580 ;
        RECT 2345.145 2588.570 2345.475 2588.585 ;
        RECT 2341.670 2588.270 2345.475 2588.570 ;
        RECT 2341.670 2588.260 2342.050 2588.270 ;
        RECT 2345.145 2588.255 2345.475 2588.270 ;
        RECT 1536.670 2587.890 1537.050 2587.900 ;
        RECT 1537.845 2587.890 1538.175 2587.905 ;
        RECT 1536.670 2587.590 1538.175 2587.890 ;
        RECT 1536.670 2587.580 1537.050 2587.590 ;
        RECT 1537.845 2587.575 1538.175 2587.590 ;
        RECT 1543.110 2587.890 1543.490 2587.900 ;
        RECT 1545.205 2587.890 1545.535 2587.905 ;
        RECT 1551.645 2587.900 1551.975 2587.905 ;
        RECT 1559.005 2587.900 1559.335 2587.905 ;
        RECT 1551.390 2587.890 1551.975 2587.900 ;
        RECT 1558.750 2587.890 1559.335 2587.900 ;
        RECT 1543.110 2587.590 1545.535 2587.890 ;
        RECT 1551.190 2587.590 1551.975 2587.890 ;
        RECT 1558.550 2587.590 1559.335 2587.890 ;
        RECT 1543.110 2587.580 1543.490 2587.590 ;
        RECT 1545.205 2587.575 1545.535 2587.590 ;
        RECT 1551.390 2587.580 1551.975 2587.590 ;
        RECT 1558.750 2587.580 1559.335 2587.590 ;
        RECT 1551.645 2587.575 1551.975 2587.580 ;
        RECT 1559.005 2587.575 1559.335 2587.580 ;
        RECT 1622.025 2587.890 1622.355 2587.905 ;
        RECT 1627.750 2587.890 1628.130 2587.900 ;
        RECT 1622.025 2587.590 1628.130 2587.890 ;
        RECT 1622.025 2587.575 1622.355 2587.590 ;
        RECT 1627.750 2587.580 1628.130 2587.590 ;
        RECT 2190.585 2587.890 2190.915 2587.905 ;
        RECT 2193.805 2587.900 2194.135 2587.905 ;
        RECT 2191.710 2587.890 2192.090 2587.900 ;
        RECT 2193.550 2587.890 2194.135 2587.900 ;
        RECT 2190.585 2587.590 2192.090 2587.890 ;
        RECT 2193.350 2587.590 2194.135 2587.890 ;
        RECT 2190.585 2587.575 2190.915 2587.590 ;
        RECT 2191.710 2587.580 2192.090 2587.590 ;
        RECT 2193.550 2587.580 2194.135 2587.590 ;
        RECT 2193.805 2587.575 2194.135 2587.580 ;
        RECT 2197.485 2587.890 2197.815 2587.905 ;
        RECT 2198.150 2587.890 2198.530 2587.900 ;
        RECT 2197.485 2587.590 2198.530 2587.890 ;
        RECT 2197.485 2587.575 2197.815 2587.590 ;
        RECT 2198.150 2587.580 2198.530 2587.590 ;
        RECT 2199.990 2587.890 2200.370 2587.900 ;
        RECT 2200.705 2587.890 2201.035 2587.905 ;
        RECT 2207.605 2587.900 2207.935 2587.905 ;
        RECT 2207.350 2587.890 2207.935 2587.900 ;
        RECT 2199.990 2587.590 2201.035 2587.890 ;
        RECT 2207.150 2587.590 2207.935 2587.890 ;
        RECT 2199.990 2587.580 2200.370 2587.590 ;
        RECT 2200.705 2587.575 2201.035 2587.590 ;
        RECT 2207.350 2587.580 2207.935 2587.590 ;
        RECT 2213.790 2587.890 2214.170 2587.900 ;
        RECT 2214.505 2587.890 2214.835 2587.905 ;
        RECT 2249.005 2587.900 2249.335 2587.905 ;
        RECT 2248.750 2587.890 2249.335 2587.900 ;
        RECT 2213.790 2587.590 2214.835 2587.890 ;
        RECT 2248.550 2587.590 2249.335 2587.890 ;
        RECT 2213.790 2587.580 2214.170 2587.590 ;
        RECT 2207.605 2587.575 2207.935 2587.580 ;
        RECT 2214.505 2587.575 2214.835 2587.590 ;
        RECT 2248.750 2587.580 2249.335 2587.590 ;
        RECT 2254.270 2587.890 2254.650 2587.900 ;
        RECT 2255.905 2587.890 2256.235 2587.905 ;
        RECT 2254.270 2587.590 2256.235 2587.890 ;
        RECT 2254.270 2587.580 2254.650 2587.590 ;
        RECT 2249.005 2587.575 2249.335 2587.580 ;
        RECT 2255.905 2587.575 2256.235 2587.590 ;
        RECT 2259.790 2587.890 2260.170 2587.900 ;
        RECT 2262.805 2587.890 2263.135 2587.905 ;
        RECT 2259.790 2587.590 2263.135 2587.890 ;
        RECT 2259.790 2587.580 2260.170 2587.590 ;
        RECT 2262.805 2587.575 2263.135 2587.590 ;
        RECT 2268.990 2587.890 2269.370 2587.900 ;
        RECT 2269.705 2587.890 2270.035 2587.905 ;
        RECT 2276.605 2587.900 2276.935 2587.905 ;
        RECT 2276.350 2587.890 2276.935 2587.900 ;
        RECT 2268.990 2587.590 2270.035 2587.890 ;
        RECT 2276.150 2587.590 2276.935 2587.890 ;
        RECT 2268.990 2587.580 2269.370 2587.590 ;
        RECT 2269.705 2587.575 2270.035 2587.590 ;
        RECT 2276.350 2587.580 2276.935 2587.590 ;
        RECT 2281.870 2587.890 2282.250 2587.900 ;
        RECT 2283.505 2587.890 2283.835 2587.905 ;
        RECT 2281.870 2587.590 2283.835 2587.890 ;
        RECT 2281.870 2587.580 2282.250 2587.590 ;
        RECT 2276.605 2587.575 2276.935 2587.580 ;
        RECT 2283.505 2587.575 2283.835 2587.590 ;
        RECT 2289.230 2587.890 2289.610 2587.900 ;
        RECT 2290.405 2587.890 2290.735 2587.905 ;
        RECT 2289.230 2587.590 2290.735 2587.890 ;
        RECT 2289.230 2587.580 2289.610 2587.590 ;
        RECT 2290.405 2587.575 2290.735 2587.590 ;
        RECT 2295.670 2587.890 2296.050 2587.900 ;
        RECT 2297.305 2587.890 2297.635 2587.905 ;
        RECT 2303.745 2587.900 2304.075 2587.905 ;
        RECT 2303.745 2587.890 2304.330 2587.900 ;
        RECT 2295.670 2587.590 2297.635 2587.890 ;
        RECT 2303.520 2587.590 2304.330 2587.890 ;
        RECT 2295.670 2587.580 2296.050 2587.590 ;
        RECT 2297.305 2587.575 2297.635 2587.590 ;
        RECT 2303.745 2587.580 2304.330 2587.590 ;
        RECT 2310.390 2587.890 2310.770 2587.900 ;
        RECT 2311.105 2587.890 2311.435 2587.905 ;
        RECT 2318.005 2587.900 2318.335 2587.905 ;
        RECT 2317.750 2587.890 2318.335 2587.900 ;
        RECT 2310.390 2587.590 2311.435 2587.890 ;
        RECT 2317.550 2587.590 2318.335 2587.890 ;
        RECT 2310.390 2587.580 2310.770 2587.590 ;
        RECT 2303.745 2587.575 2304.075 2587.580 ;
        RECT 2311.105 2587.575 2311.435 2587.590 ;
        RECT 2317.750 2587.580 2318.335 2587.590 ;
        RECT 2324.190 2587.890 2324.570 2587.900 ;
        RECT 2324.905 2587.890 2325.235 2587.905 ;
        RECT 2324.190 2587.590 2325.235 2587.890 ;
        RECT 2324.190 2587.580 2324.570 2587.590 ;
        RECT 2318.005 2587.575 2318.335 2587.580 ;
        RECT 2324.905 2587.575 2325.235 2587.590 ;
        RECT 2330.630 2587.890 2331.010 2587.900 ;
        RECT 2331.805 2587.890 2332.135 2587.905 ;
        RECT 2330.630 2587.590 2332.135 2587.890 ;
        RECT 2330.630 2587.580 2331.010 2587.590 ;
        RECT 2331.805 2587.575 2332.135 2587.590 ;
        RECT 2336.150 2587.890 2336.530 2587.900 ;
        RECT 2338.705 2587.890 2339.035 2587.905 ;
        RECT 2345.605 2587.900 2345.935 2587.905 ;
        RECT 2345.350 2587.890 2345.935 2587.900 ;
        RECT 2336.150 2587.590 2339.035 2587.890 ;
        RECT 2345.150 2587.590 2345.935 2587.890 ;
        RECT 2336.150 2587.580 2336.530 2587.590 ;
        RECT 2338.705 2587.575 2339.035 2587.590 ;
        RECT 2345.350 2587.580 2345.935 2587.590 ;
        RECT 2345.605 2587.575 2345.935 2587.580 ;
        RECT 2169.630 2477.730 2170.010 2477.740 ;
        RECT 2170.345 2477.730 2170.675 2477.745 ;
        RECT 2169.630 2477.430 2170.675 2477.730 ;
        RECT 2169.630 2477.420 2170.010 2477.430 ;
        RECT 2170.345 2477.415 2170.675 2477.430 ;
        RECT 2169.425 2463.460 2169.755 2463.465 ;
        RECT 2169.425 2463.450 2170.010 2463.460 ;
        RECT 2169.425 2463.150 2170.210 2463.450 ;
        RECT 2169.425 2463.140 2170.010 2463.150 ;
        RECT 2169.425 2463.135 2169.755 2463.140 ;
        RECT 2168.045 2415.170 2168.375 2415.185 ;
        RECT 2168.965 2415.170 2169.295 2415.185 ;
        RECT 2168.045 2414.870 2169.295 2415.170 ;
        RECT 2168.045 2414.855 2168.375 2414.870 ;
        RECT 2168.965 2414.855 2169.295 2414.870 ;
        RECT 2331.805 2412.450 2332.135 2412.465 ;
        RECT 2654.265 2412.450 2654.595 2412.465 ;
        RECT 2331.805 2412.150 2654.595 2412.450 ;
        RECT 2331.805 2412.135 2332.135 2412.150 ;
        RECT 2654.265 2412.135 2654.595 2412.150 ;
        RECT 2345.145 2411.770 2345.475 2411.785 ;
        RECT 2680.025 2411.770 2680.355 2411.785 ;
        RECT 2345.145 2411.470 2680.355 2411.770 ;
        RECT 2345.145 2411.455 2345.475 2411.470 ;
        RECT 2680.025 2411.455 2680.355 2411.470 ;
        RECT 1318.425 2411.090 1318.755 2411.105 ;
        RECT 1898.485 2411.090 1898.815 2411.105 ;
        RECT 1318.425 2410.790 1898.815 2411.090 ;
        RECT 1318.425 2410.775 1318.755 2410.790 ;
        RECT 1898.485 2410.775 1898.815 2410.790 ;
        RECT 2345.605 2411.090 2345.935 2411.105 ;
        RECT 2692.905 2411.090 2693.235 2411.105 ;
        RECT 2345.605 2410.790 2693.235 2411.090 ;
        RECT 2345.605 2410.775 2345.935 2410.790 ;
        RECT 2692.905 2410.775 2693.235 2410.790 ;
        RECT 1600.865 2410.410 1601.195 2410.425 ;
        RECT 1607.765 2410.410 1608.095 2410.425 ;
        RECT 1600.865 2410.110 1608.095 2410.410 ;
        RECT 1600.865 2410.095 1601.195 2410.110 ;
        RECT 1607.765 2410.095 1608.095 2410.110 ;
        RECT 2356.185 2409.050 2356.515 2409.065 ;
        RECT 2386.085 2409.050 2386.415 2409.065 ;
        RECT 2356.185 2408.750 2386.415 2409.050 ;
        RECT 2356.185 2408.735 2356.515 2408.750 ;
        RECT 2386.085 2408.735 2386.415 2408.750 ;
      LAYER met3 ;
        RECT 1304.400 2393.720 2695.600 2394.585 ;
        RECT 1303.990 2384.920 2696.000 2393.720 ;
        RECT 1303.990 2384.240 2695.600 2384.920 ;
        RECT 1304.400 2383.520 2695.600 2384.240 ;
        RECT 1304.400 2382.840 2696.000 2383.520 ;
        RECT 1303.990 2374.040 2696.000 2382.840 ;
        RECT 1304.400 2372.640 2695.600 2374.040 ;
        RECT 1303.990 2363.840 2696.000 2372.640 ;
        RECT 1303.990 2363.160 2695.600 2363.840 ;
        RECT 1304.400 2362.440 2695.600 2363.160 ;
        RECT 1304.400 2361.760 2696.000 2362.440 ;
        RECT 1303.990 2352.960 2696.000 2361.760 ;
        RECT 1303.990 2352.280 2695.600 2352.960 ;
        RECT 1304.400 2351.560 2695.600 2352.280 ;
        RECT 1304.400 2350.880 2696.000 2351.560 ;
        RECT 1303.990 2342.760 2696.000 2350.880 ;
        RECT 1303.990 2342.080 2695.600 2342.760 ;
        RECT 1304.400 2341.360 2695.600 2342.080 ;
        RECT 1304.400 2340.680 2696.000 2341.360 ;
        RECT 1303.990 2331.880 2696.000 2340.680 ;
        RECT 1303.990 2331.200 2695.600 2331.880 ;
        RECT 1304.400 2330.480 2695.600 2331.200 ;
        RECT 1304.400 2329.800 2696.000 2330.480 ;
        RECT 1303.990 2321.680 2696.000 2329.800 ;
        RECT 1303.990 2321.000 2695.600 2321.680 ;
        RECT 1304.400 2320.280 2695.600 2321.000 ;
        RECT 1304.400 2319.600 2696.000 2320.280 ;
        RECT 1303.990 2310.800 2696.000 2319.600 ;
        RECT 1303.990 2310.120 2695.600 2310.800 ;
        RECT 1304.400 2309.400 2695.600 2310.120 ;
        RECT 1304.400 2308.720 2696.000 2309.400 ;
        RECT 1303.990 2300.600 2696.000 2308.720 ;
        RECT 1303.990 2299.240 2695.600 2300.600 ;
        RECT 1304.400 2299.200 2695.600 2299.240 ;
        RECT 1304.400 2297.840 2696.000 2299.200 ;
        RECT 1303.990 2289.720 2696.000 2297.840 ;
        RECT 1303.990 2289.040 2695.600 2289.720 ;
        RECT 1304.400 2288.320 2695.600 2289.040 ;
        RECT 1304.400 2287.640 2696.000 2288.320 ;
        RECT 1303.990 2279.520 2696.000 2287.640 ;
        RECT 1303.990 2278.160 2695.600 2279.520 ;
        RECT 1304.400 2278.120 2695.600 2278.160 ;
        RECT 1304.400 2276.760 2696.000 2278.120 ;
        RECT 1303.990 2268.640 2696.000 2276.760 ;
        RECT 1303.990 2267.280 2695.600 2268.640 ;
        RECT 1304.400 2267.240 2695.600 2267.280 ;
        RECT 1304.400 2265.880 2696.000 2267.240 ;
        RECT 1303.990 2258.440 2696.000 2265.880 ;
        RECT 1303.990 2257.080 2695.600 2258.440 ;
        RECT 1304.400 2257.040 2695.600 2257.080 ;
        RECT 1304.400 2255.680 2696.000 2257.040 ;
        RECT 1303.990 2247.560 2696.000 2255.680 ;
        RECT 1303.990 2246.200 2695.600 2247.560 ;
        RECT 1304.400 2246.160 2695.600 2246.200 ;
        RECT 1304.400 2244.800 2696.000 2246.160 ;
        RECT 1303.990 2237.360 2696.000 2244.800 ;
        RECT 1303.990 2236.000 2695.600 2237.360 ;
        RECT 1304.400 2235.960 2695.600 2236.000 ;
        RECT 1304.400 2234.600 2696.000 2235.960 ;
        RECT 1303.990 2226.480 2696.000 2234.600 ;
        RECT 1303.990 2225.120 2695.600 2226.480 ;
        RECT 1304.400 2225.080 2695.600 2225.120 ;
        RECT 1304.400 2223.720 2696.000 2225.080 ;
        RECT 1303.990 2216.280 2696.000 2223.720 ;
        RECT 1303.990 2214.880 2695.600 2216.280 ;
        RECT 1303.990 2214.240 2696.000 2214.880 ;
        RECT 1304.400 2212.840 2696.000 2214.240 ;
        RECT 1303.990 2205.400 2696.000 2212.840 ;
        RECT 1303.990 2204.040 2695.600 2205.400 ;
        RECT 1304.400 2204.000 2695.600 2204.040 ;
        RECT 1304.400 2202.640 2696.000 2204.000 ;
        RECT 1303.990 2195.200 2696.000 2202.640 ;
        RECT 1303.990 2193.800 2695.600 2195.200 ;
        RECT 1303.990 2193.160 2696.000 2193.800 ;
        RECT 1304.400 2191.760 2696.000 2193.160 ;
        RECT 1303.990 2184.320 2696.000 2191.760 ;
        RECT 1303.990 2182.920 2695.600 2184.320 ;
        RECT 1303.990 2182.280 2696.000 2182.920 ;
        RECT 1304.400 2180.880 2696.000 2182.280 ;
        RECT 1303.990 2174.120 2696.000 2180.880 ;
        RECT 1303.990 2172.720 2695.600 2174.120 ;
        RECT 1303.990 2172.080 2696.000 2172.720 ;
        RECT 1304.400 2170.680 2696.000 2172.080 ;
        RECT 1303.990 2163.240 2696.000 2170.680 ;
        RECT 1303.990 2161.840 2695.600 2163.240 ;
        RECT 1303.990 2161.200 2696.000 2161.840 ;
        RECT 1304.400 2159.800 2696.000 2161.200 ;
        RECT 1303.990 2153.040 2696.000 2159.800 ;
        RECT 1303.990 2151.640 2695.600 2153.040 ;
        RECT 1303.990 2151.000 2696.000 2151.640 ;
        RECT 1304.400 2149.600 2696.000 2151.000 ;
        RECT 1303.990 2142.160 2696.000 2149.600 ;
        RECT 1303.990 2140.760 2695.600 2142.160 ;
        RECT 1303.990 2140.120 2696.000 2140.760 ;
        RECT 1304.400 2138.720 2696.000 2140.120 ;
        RECT 1303.990 2131.960 2696.000 2138.720 ;
        RECT 1303.990 2130.560 2695.600 2131.960 ;
        RECT 1303.990 2129.240 2696.000 2130.560 ;
        RECT 1304.400 2127.840 2696.000 2129.240 ;
        RECT 1303.990 2121.080 2696.000 2127.840 ;
        RECT 1303.990 2119.680 2695.600 2121.080 ;
        RECT 1303.990 2119.040 2696.000 2119.680 ;
        RECT 1304.400 2117.640 2696.000 2119.040 ;
        RECT 1303.990 2110.880 2696.000 2117.640 ;
        RECT 1303.990 2109.480 2695.600 2110.880 ;
        RECT 1303.990 2108.160 2696.000 2109.480 ;
        RECT 1304.400 2106.760 2696.000 2108.160 ;
        RECT 1303.990 2100.680 2696.000 2106.760 ;
        RECT 1303.990 2099.280 2695.600 2100.680 ;
        RECT 1303.990 2097.960 2696.000 2099.280 ;
        RECT 1304.400 2096.560 2696.000 2097.960 ;
        RECT 1303.990 2089.800 2696.000 2096.560 ;
        RECT 1303.990 2088.400 2695.600 2089.800 ;
        RECT 1303.990 2087.080 2696.000 2088.400 ;
        RECT 1304.400 2085.680 2696.000 2087.080 ;
        RECT 1303.990 2079.600 2696.000 2085.680 ;
        RECT 1303.990 2078.200 2695.600 2079.600 ;
        RECT 1303.990 2076.200 2696.000 2078.200 ;
        RECT 1304.400 2074.800 2696.000 2076.200 ;
        RECT 1303.990 2068.720 2696.000 2074.800 ;
        RECT 1303.990 2067.320 2695.600 2068.720 ;
        RECT 1303.990 2066.000 2696.000 2067.320 ;
        RECT 1304.400 2064.600 2696.000 2066.000 ;
        RECT 1303.990 2058.520 2696.000 2064.600 ;
        RECT 1303.990 2057.120 2695.600 2058.520 ;
        RECT 1303.990 2055.120 2696.000 2057.120 ;
        RECT 1304.400 2053.720 2696.000 2055.120 ;
        RECT 1303.990 2047.640 2696.000 2053.720 ;
        RECT 1303.990 2046.240 2695.600 2047.640 ;
        RECT 1303.990 2044.240 2696.000 2046.240 ;
        RECT 1304.400 2042.840 2696.000 2044.240 ;
        RECT 1303.990 2037.440 2696.000 2042.840 ;
        RECT 1303.990 2036.040 2695.600 2037.440 ;
        RECT 1303.990 2034.040 2696.000 2036.040 ;
        RECT 1304.400 2032.640 2696.000 2034.040 ;
        RECT 1303.990 2026.560 2696.000 2032.640 ;
        RECT 1303.990 2025.160 2695.600 2026.560 ;
        RECT 1303.990 2023.160 2696.000 2025.160 ;
        RECT 1304.400 2021.760 2696.000 2023.160 ;
        RECT 1303.990 2016.360 2696.000 2021.760 ;
        RECT 1303.990 2014.960 2695.600 2016.360 ;
        RECT 1303.990 2012.960 2696.000 2014.960 ;
        RECT 1304.400 2011.560 2696.000 2012.960 ;
        RECT 1303.990 2005.480 2696.000 2011.560 ;
        RECT 1303.990 2004.080 2695.600 2005.480 ;
        RECT 1303.990 2002.080 2696.000 2004.080 ;
        RECT 1304.400 2000.680 2696.000 2002.080 ;
        RECT 1303.990 1995.280 2696.000 2000.680 ;
        RECT 1303.990 1993.880 2695.600 1995.280 ;
        RECT 1303.990 1991.200 2696.000 1993.880 ;
        RECT 1304.400 1989.800 2696.000 1991.200 ;
        RECT 1303.990 1984.400 2696.000 1989.800 ;
        RECT 1303.990 1983.000 2695.600 1984.400 ;
        RECT 1303.990 1981.000 2696.000 1983.000 ;
        RECT 1304.400 1979.600 2696.000 1981.000 ;
        RECT 1303.990 1974.200 2696.000 1979.600 ;
        RECT 1303.990 1972.800 2695.600 1974.200 ;
        RECT 1303.990 1970.120 2696.000 1972.800 ;
        RECT 1304.400 1968.720 2696.000 1970.120 ;
        RECT 1303.990 1963.320 2696.000 1968.720 ;
        RECT 1303.990 1961.920 2695.600 1963.320 ;
        RECT 1303.990 1959.240 2696.000 1961.920 ;
        RECT 1304.400 1957.840 2696.000 1959.240 ;
        RECT 1303.990 1953.120 2696.000 1957.840 ;
        RECT 1303.990 1951.720 2695.600 1953.120 ;
        RECT 1303.990 1949.040 2696.000 1951.720 ;
        RECT 1304.400 1947.640 2696.000 1949.040 ;
        RECT 1303.990 1942.240 2696.000 1947.640 ;
        RECT 1303.990 1940.840 2695.600 1942.240 ;
        RECT 1303.990 1938.160 2696.000 1940.840 ;
        RECT 1304.400 1936.760 2696.000 1938.160 ;
        RECT 1303.990 1932.040 2696.000 1936.760 ;
        RECT 1303.990 1930.640 2695.600 1932.040 ;
        RECT 1303.990 1927.960 2696.000 1930.640 ;
        RECT 1304.400 1926.560 2696.000 1927.960 ;
        RECT 1303.990 1921.160 2696.000 1926.560 ;
        RECT 1303.990 1919.760 2695.600 1921.160 ;
        RECT 1303.990 1917.080 2696.000 1919.760 ;
        RECT 1304.400 1915.680 2696.000 1917.080 ;
        RECT 1303.990 1910.960 2696.000 1915.680 ;
        RECT 1303.990 1909.560 2695.600 1910.960 ;
        RECT 1303.990 1906.200 2696.000 1909.560 ;
        RECT 1304.400 1904.800 2696.000 1906.200 ;
        RECT 1303.990 1900.080 2696.000 1904.800 ;
        RECT 1303.990 1898.680 2695.600 1900.080 ;
        RECT 1303.990 1896.000 2696.000 1898.680 ;
        RECT 1304.400 1894.600 2696.000 1896.000 ;
        RECT 1303.990 1889.880 2696.000 1894.600 ;
        RECT 1303.990 1888.480 2695.600 1889.880 ;
        RECT 1303.990 1885.120 2696.000 1888.480 ;
        RECT 1304.400 1883.720 2696.000 1885.120 ;
        RECT 1303.990 1879.000 2696.000 1883.720 ;
        RECT 1303.990 1877.600 2695.600 1879.000 ;
        RECT 1303.990 1874.920 2696.000 1877.600 ;
        RECT 1304.400 1873.520 2696.000 1874.920 ;
        RECT 1303.990 1868.800 2696.000 1873.520 ;
        RECT 1303.990 1867.400 2695.600 1868.800 ;
        RECT 1303.990 1864.040 2696.000 1867.400 ;
        RECT 1304.400 1862.640 2696.000 1864.040 ;
        RECT 1303.990 1857.920 2696.000 1862.640 ;
        RECT 1303.990 1856.520 2695.600 1857.920 ;
        RECT 1303.990 1853.160 2696.000 1856.520 ;
        RECT 1304.400 1851.760 2696.000 1853.160 ;
        RECT 1303.990 1847.720 2696.000 1851.760 ;
        RECT 1303.990 1846.320 2695.600 1847.720 ;
        RECT 1303.990 1842.960 2696.000 1846.320 ;
        RECT 1304.400 1841.560 2696.000 1842.960 ;
        RECT 1303.990 1836.840 2696.000 1841.560 ;
        RECT 1303.990 1835.440 2695.600 1836.840 ;
        RECT 1303.990 1832.080 2696.000 1835.440 ;
        RECT 1304.400 1830.680 2696.000 1832.080 ;
        RECT 1303.990 1826.640 2696.000 1830.680 ;
        RECT 1303.990 1825.240 2695.600 1826.640 ;
        RECT 1303.990 1821.200 2696.000 1825.240 ;
        RECT 1304.400 1819.800 2696.000 1821.200 ;
        RECT 1303.990 1815.760 2696.000 1819.800 ;
        RECT 1303.990 1814.360 2695.600 1815.760 ;
        RECT 1303.990 1811.000 2696.000 1814.360 ;
        RECT 1304.400 1809.600 2696.000 1811.000 ;
        RECT 1303.990 1805.560 2696.000 1809.600 ;
        RECT 1303.990 1804.160 2695.600 1805.560 ;
        RECT 1303.990 1800.120 2696.000 1804.160 ;
        RECT 1304.400 1798.720 2696.000 1800.120 ;
        RECT 1303.990 1795.360 2696.000 1798.720 ;
        RECT 1303.990 1793.960 2695.600 1795.360 ;
        RECT 1303.990 1789.920 2696.000 1793.960 ;
        RECT 1304.400 1788.520 2696.000 1789.920 ;
        RECT 1303.990 1784.480 2696.000 1788.520 ;
        RECT 1303.990 1783.080 2695.600 1784.480 ;
        RECT 1303.990 1779.040 2696.000 1783.080 ;
        RECT 1304.400 1777.640 2696.000 1779.040 ;
        RECT 1303.990 1774.280 2696.000 1777.640 ;
        RECT 1303.990 1772.880 2695.600 1774.280 ;
        RECT 1303.990 1768.160 2696.000 1772.880 ;
        RECT 1304.400 1766.760 2696.000 1768.160 ;
        RECT 1303.990 1763.400 2696.000 1766.760 ;
        RECT 1303.990 1762.000 2695.600 1763.400 ;
        RECT 1303.990 1757.960 2696.000 1762.000 ;
        RECT 1304.400 1756.560 2696.000 1757.960 ;
        RECT 1303.990 1753.200 2696.000 1756.560 ;
        RECT 1303.990 1751.800 2695.600 1753.200 ;
        RECT 1303.990 1747.080 2696.000 1751.800 ;
        RECT 1304.400 1745.680 2696.000 1747.080 ;
        RECT 1303.990 1742.320 2696.000 1745.680 ;
        RECT 1303.990 1740.920 2695.600 1742.320 ;
        RECT 1303.990 1736.200 2696.000 1740.920 ;
        RECT 1304.400 1734.800 2696.000 1736.200 ;
        RECT 1303.990 1732.120 2696.000 1734.800 ;
        RECT 1303.990 1730.720 2695.600 1732.120 ;
        RECT 1303.990 1726.000 2696.000 1730.720 ;
        RECT 1304.400 1724.600 2696.000 1726.000 ;
        RECT 1303.990 1721.240 2696.000 1724.600 ;
        RECT 1303.990 1719.840 2695.600 1721.240 ;
        RECT 1303.990 1715.120 2696.000 1719.840 ;
        RECT 1304.400 1713.720 2696.000 1715.120 ;
        RECT 1303.990 1711.040 2696.000 1713.720 ;
        RECT 1303.990 1709.640 2695.600 1711.040 ;
        RECT 1303.990 1704.920 2696.000 1709.640 ;
        RECT 1304.400 1703.520 2696.000 1704.920 ;
        RECT 1303.990 1700.160 2696.000 1703.520 ;
        RECT 1303.990 1698.760 2695.600 1700.160 ;
        RECT 1303.990 1694.040 2696.000 1698.760 ;
        RECT 1304.400 1692.640 2696.000 1694.040 ;
        RECT 1303.990 1689.960 2696.000 1692.640 ;
        RECT 1303.990 1688.560 2695.600 1689.960 ;
        RECT 1303.990 1683.160 2696.000 1688.560 ;
        RECT 1304.400 1681.760 2696.000 1683.160 ;
        RECT 1303.990 1679.080 2696.000 1681.760 ;
        RECT 1303.990 1677.680 2695.600 1679.080 ;
        RECT 1303.990 1672.960 2696.000 1677.680 ;
        RECT 1304.400 1671.560 2696.000 1672.960 ;
        RECT 1303.990 1668.880 2696.000 1671.560 ;
        RECT 1303.990 1667.480 2695.600 1668.880 ;
        RECT 1303.990 1662.080 2696.000 1667.480 ;
        RECT 1304.400 1660.680 2696.000 1662.080 ;
        RECT 1303.990 1658.000 2696.000 1660.680 ;
        RECT 1303.990 1656.600 2695.600 1658.000 ;
        RECT 1303.990 1651.880 2696.000 1656.600 ;
        RECT 1304.400 1650.480 2696.000 1651.880 ;
        RECT 1303.990 1647.800 2696.000 1650.480 ;
        RECT 1303.990 1646.400 2695.600 1647.800 ;
        RECT 1303.990 1641.000 2696.000 1646.400 ;
        RECT 1304.400 1639.600 2696.000 1641.000 ;
        RECT 1303.990 1636.920 2696.000 1639.600 ;
        RECT 1303.990 1635.520 2695.600 1636.920 ;
        RECT 1303.990 1630.120 2696.000 1635.520 ;
        RECT 1304.400 1628.720 2696.000 1630.120 ;
        RECT 1303.990 1626.720 2696.000 1628.720 ;
        RECT 1303.990 1625.320 2695.600 1626.720 ;
        RECT 1303.990 1619.920 2696.000 1625.320 ;
        RECT 1304.400 1618.520 2696.000 1619.920 ;
        RECT 1303.990 1615.840 2696.000 1618.520 ;
        RECT 1303.990 1614.440 2695.600 1615.840 ;
        RECT 1303.990 1609.040 2696.000 1614.440 ;
        RECT 1304.400 1607.640 2696.000 1609.040 ;
        RECT 1303.990 1605.640 2696.000 1607.640 ;
        RECT 1303.990 1604.240 2695.600 1605.640 ;
        RECT 1303.990 1598.160 2696.000 1604.240 ;
        RECT 1304.400 1596.760 2696.000 1598.160 ;
        RECT 1303.990 1594.760 2696.000 1596.760 ;
        RECT 1303.990 1593.360 2695.600 1594.760 ;
        RECT 1303.990 1587.960 2696.000 1593.360 ;
        RECT 1304.400 1586.560 2696.000 1587.960 ;
        RECT 1303.990 1584.560 2696.000 1586.560 ;
        RECT 1303.990 1583.160 2695.600 1584.560 ;
        RECT 1303.990 1577.080 2696.000 1583.160 ;
        RECT 1304.400 1575.680 2696.000 1577.080 ;
        RECT 1303.990 1573.680 2696.000 1575.680 ;
        RECT 1303.990 1572.280 2695.600 1573.680 ;
        RECT 1303.990 1566.880 2696.000 1572.280 ;
        RECT 1304.400 1565.480 2696.000 1566.880 ;
        RECT 1303.990 1563.480 2696.000 1565.480 ;
        RECT 1303.990 1562.080 2695.600 1563.480 ;
        RECT 1303.990 1556.000 2696.000 1562.080 ;
        RECT 1304.400 1554.600 2696.000 1556.000 ;
        RECT 1303.990 1552.600 2696.000 1554.600 ;
        RECT 1303.990 1551.200 2695.600 1552.600 ;
        RECT 1303.990 1545.120 2696.000 1551.200 ;
        RECT 1304.400 1543.720 2696.000 1545.120 ;
        RECT 1303.990 1542.400 2696.000 1543.720 ;
        RECT 1303.990 1541.000 2695.600 1542.400 ;
        RECT 1303.990 1534.920 2696.000 1541.000 ;
        RECT 1304.400 1533.520 2696.000 1534.920 ;
        RECT 1303.990 1531.520 2696.000 1533.520 ;
        RECT 1303.990 1530.120 2695.600 1531.520 ;
        RECT 1303.990 1524.040 2696.000 1530.120 ;
        RECT 1304.400 1522.640 2696.000 1524.040 ;
        RECT 1303.990 1521.320 2696.000 1522.640 ;
        RECT 1303.990 1519.920 2695.600 1521.320 ;
        RECT 1303.990 1513.160 2696.000 1519.920 ;
        RECT 1304.400 1511.760 2696.000 1513.160 ;
        RECT 1303.990 1510.440 2696.000 1511.760 ;
        RECT 1303.990 1509.040 2695.600 1510.440 ;
        RECT 1303.990 1502.960 2696.000 1509.040 ;
        RECT 1304.400 1501.560 2696.000 1502.960 ;
        RECT 1303.990 1500.240 2696.000 1501.560 ;
        RECT 1303.990 1498.840 2695.600 1500.240 ;
        RECT 1303.990 1492.080 2696.000 1498.840 ;
        RECT 1304.400 1490.680 2696.000 1492.080 ;
        RECT 1303.990 1490.040 2696.000 1490.680 ;
        RECT 1303.990 1488.640 2695.600 1490.040 ;
        RECT 1303.990 1481.880 2696.000 1488.640 ;
        RECT 1304.400 1480.480 2696.000 1481.880 ;
        RECT 1303.990 1479.160 2696.000 1480.480 ;
        RECT 1303.990 1477.760 2695.600 1479.160 ;
        RECT 1303.990 1471.000 2696.000 1477.760 ;
        RECT 1304.400 1469.600 2696.000 1471.000 ;
        RECT 1303.990 1468.960 2696.000 1469.600 ;
        RECT 1303.990 1467.560 2695.600 1468.960 ;
        RECT 1303.990 1460.120 2696.000 1467.560 ;
        RECT 1304.400 1458.720 2696.000 1460.120 ;
        RECT 1303.990 1458.080 2696.000 1458.720 ;
        RECT 1303.990 1456.680 2695.600 1458.080 ;
        RECT 1303.990 1449.920 2696.000 1456.680 ;
        RECT 1304.400 1448.520 2696.000 1449.920 ;
        RECT 1303.990 1447.880 2696.000 1448.520 ;
        RECT 1303.990 1446.480 2695.600 1447.880 ;
        RECT 1303.990 1439.040 2696.000 1446.480 ;
        RECT 1304.400 1437.640 2696.000 1439.040 ;
        RECT 1303.990 1437.000 2696.000 1437.640 ;
        RECT 1303.990 1435.600 2695.600 1437.000 ;
        RECT 1303.990 1428.840 2696.000 1435.600 ;
        RECT 1304.400 1427.440 2696.000 1428.840 ;
        RECT 1303.990 1426.800 2696.000 1427.440 ;
        RECT 1303.990 1425.400 2695.600 1426.800 ;
        RECT 1303.990 1417.960 2696.000 1425.400 ;
        RECT 1304.400 1416.560 2696.000 1417.960 ;
        RECT 1303.990 1415.920 2696.000 1416.560 ;
        RECT 1303.990 1414.520 2695.600 1415.920 ;
        RECT 1303.990 1407.080 2696.000 1414.520 ;
        RECT 1304.400 1405.720 2696.000 1407.080 ;
        RECT 1304.400 1405.680 2695.600 1405.720 ;
        RECT 1303.990 1404.320 2695.600 1405.680 ;
        RECT 1303.990 1396.880 2696.000 1404.320 ;
        RECT 1304.400 1395.480 2696.000 1396.880 ;
        RECT 1303.990 1394.840 2696.000 1395.480 ;
        RECT 1303.990 1393.440 2695.600 1394.840 ;
        RECT 1303.990 1386.000 2696.000 1393.440 ;
        RECT 1304.400 1384.640 2696.000 1386.000 ;
        RECT 1304.400 1384.600 2695.600 1384.640 ;
        RECT 1303.990 1383.240 2695.600 1384.600 ;
        RECT 1303.990 1375.120 2696.000 1383.240 ;
        RECT 1304.400 1373.760 2696.000 1375.120 ;
        RECT 1304.400 1373.720 2695.600 1373.760 ;
        RECT 1303.990 1372.360 2695.600 1373.720 ;
        RECT 1303.990 1364.920 2696.000 1372.360 ;
        RECT 1304.400 1363.560 2696.000 1364.920 ;
        RECT 1304.400 1363.520 2695.600 1363.560 ;
        RECT 1303.990 1362.160 2695.600 1363.520 ;
        RECT 1303.990 1354.040 2696.000 1362.160 ;
        RECT 1304.400 1352.680 2696.000 1354.040 ;
        RECT 1304.400 1352.640 2695.600 1352.680 ;
        RECT 1303.990 1351.280 2695.600 1352.640 ;
        RECT 1303.990 1343.840 2696.000 1351.280 ;
        RECT 1304.400 1342.480 2696.000 1343.840 ;
        RECT 1304.400 1342.440 2695.600 1342.480 ;
        RECT 1303.990 1341.080 2695.600 1342.440 ;
        RECT 1303.990 1332.960 2696.000 1341.080 ;
        RECT 1304.400 1331.600 2696.000 1332.960 ;
        RECT 1304.400 1331.560 2695.600 1331.600 ;
        RECT 1303.990 1330.200 2695.600 1331.560 ;
        RECT 1303.990 1322.080 2696.000 1330.200 ;
        RECT 1304.400 1321.400 2696.000 1322.080 ;
        RECT 1304.400 1320.680 2695.600 1321.400 ;
        RECT 1303.990 1320.000 2695.600 1320.680 ;
        RECT 1303.990 1311.880 2696.000 1320.000 ;
        RECT 1304.400 1310.520 2696.000 1311.880 ;
        RECT 1304.400 1310.480 2695.600 1310.520 ;
        RECT 1303.990 1309.120 2695.600 1310.480 ;
        RECT 1303.990 1301.000 2696.000 1309.120 ;
        RECT 1304.400 1300.320 2696.000 1301.000 ;
        RECT 1304.400 1299.600 2695.600 1300.320 ;
        RECT 1303.990 1298.920 2695.600 1299.600 ;
        RECT 1303.990 1290.120 2696.000 1298.920 ;
        RECT 1304.400 1289.440 2696.000 1290.120 ;
        RECT 1304.400 1288.720 2695.600 1289.440 ;
        RECT 1303.990 1288.040 2695.600 1288.720 ;
        RECT 1303.990 1279.920 2696.000 1288.040 ;
        RECT 1304.400 1279.240 2696.000 1279.920 ;
        RECT 1304.400 1278.520 2695.600 1279.240 ;
        RECT 1303.990 1277.840 2695.600 1278.520 ;
        RECT 1303.990 1269.040 2696.000 1277.840 ;
        RECT 1304.400 1268.360 2696.000 1269.040 ;
        RECT 1304.400 1267.640 2695.600 1268.360 ;
        RECT 1303.990 1266.960 2695.600 1267.640 ;
        RECT 1303.990 1258.840 2696.000 1266.960 ;
        RECT 1304.400 1258.160 2696.000 1258.840 ;
        RECT 1304.400 1257.440 2695.600 1258.160 ;
        RECT 1303.990 1256.760 2695.600 1257.440 ;
        RECT 1303.990 1247.960 2696.000 1256.760 ;
        RECT 1304.400 1247.280 2696.000 1247.960 ;
        RECT 1304.400 1246.560 2695.600 1247.280 ;
        RECT 1303.990 1245.880 2695.600 1246.560 ;
        RECT 1303.990 1237.080 2696.000 1245.880 ;
        RECT 1304.400 1235.680 2695.600 1237.080 ;
        RECT 1303.990 1226.880 2696.000 1235.680 ;
        RECT 1304.400 1226.200 2696.000 1226.880 ;
        RECT 1304.400 1225.480 2695.600 1226.200 ;
        RECT 1303.990 1224.800 2695.600 1225.480 ;
        RECT 1303.990 1216.000 2696.000 1224.800 ;
        RECT 1304.400 1214.600 2695.600 1216.000 ;
        RECT 1303.990 1205.800 2696.000 1214.600 ;
        RECT 1304.400 1204.950 2695.600 1205.800 ;
      LAYER met3 ;
        RECT 2370.190 1038.850 2370.570 1038.860 ;
        RECT 2384.705 1038.850 2385.035 1038.865 ;
        RECT 2370.190 1038.550 2385.035 1038.850 ;
        RECT 2370.190 1038.540 2370.570 1038.550 ;
        RECT 2384.705 1038.535 2385.035 1038.550 ;
        RECT 1386.505 1021.170 1386.835 1021.185 ;
        RECT 1796.110 1021.170 1796.490 1021.180 ;
        RECT 1386.505 1020.870 1796.490 1021.170 ;
        RECT 1386.505 1020.855 1386.835 1020.870 ;
        RECT 1796.110 1020.860 1796.490 1020.870 ;
        RECT 1830.150 1021.170 1830.530 1021.180 ;
        RECT 1831.785 1021.170 1832.115 1021.185 ;
        RECT 1830.150 1020.870 1832.115 1021.170 ;
        RECT 1830.150 1020.860 1830.530 1020.870 ;
        RECT 1831.785 1020.855 1832.115 1020.870 ;
        RECT 1854.990 1021.170 1855.370 1021.180 ;
        RECT 1855.705 1021.170 1856.035 1021.185 ;
        RECT 2283.045 1021.180 2283.375 1021.185 ;
        RECT 1854.990 1020.870 1856.035 1021.170 ;
        RECT 1854.990 1020.860 1855.370 1020.870 ;
        RECT 1855.705 1020.855 1856.035 1020.870 ;
        RECT 2282.790 1021.170 2283.375 1021.180 ;
        RECT 2340.750 1021.170 2341.130 1021.180 ;
        RECT 2345.605 1021.170 2345.935 1021.185 ;
        RECT 2282.790 1020.870 2283.600 1021.170 ;
        RECT 2340.750 1020.870 2345.935 1021.170 ;
        RECT 2282.790 1020.860 2283.375 1020.870 ;
        RECT 2340.750 1020.860 2341.130 1020.870 ;
        RECT 2283.045 1020.855 2283.375 1020.860 ;
        RECT 2345.605 1020.855 2345.935 1020.870 ;
        RECT 2351.790 1021.170 2352.170 1021.180 ;
        RECT 2352.505 1021.170 2352.835 1021.185 ;
        RECT 2387.465 1021.180 2387.795 1021.185 ;
        RECT 2387.465 1021.170 2388.050 1021.180 ;
        RECT 2351.790 1020.870 2352.835 1021.170 ;
        RECT 2387.240 1020.870 2388.050 1021.170 ;
        RECT 2351.790 1020.860 2352.170 1020.870 ;
        RECT 2352.505 1020.855 2352.835 1020.870 ;
        RECT 2387.465 1020.860 2388.050 1020.870 ;
        RECT 2390.685 1021.170 2391.015 1021.185 ;
        RECT 2395.950 1021.170 2396.330 1021.180 ;
        RECT 2390.685 1020.870 2396.330 1021.170 ;
        RECT 2387.465 1020.855 2387.795 1020.860 ;
        RECT 2390.685 1020.855 2391.015 1020.870 ;
        RECT 2395.950 1020.860 2396.330 1020.870 ;
        RECT 2408.165 1021.170 2408.495 1021.185 ;
        RECT 2450.945 1021.180 2451.275 1021.185 ;
        RECT 2408.830 1021.170 2409.210 1021.180 ;
        RECT 2450.945 1021.170 2451.530 1021.180 ;
        RECT 2408.165 1020.870 2409.210 1021.170 ;
        RECT 2450.720 1020.870 2451.530 1021.170 ;
        RECT 2408.165 1020.855 2408.495 1020.870 ;
        RECT 2408.830 1020.860 2409.210 1020.870 ;
        RECT 2450.945 1020.860 2451.530 1020.870 ;
        RECT 2450.945 1020.855 2451.275 1020.860 ;
        RECT 1372.705 1020.490 1373.035 1020.505 ;
        RECT 1801.630 1020.490 1802.010 1020.500 ;
        RECT 1372.705 1020.190 1802.010 1020.490 ;
        RECT 1372.705 1020.175 1373.035 1020.190 ;
        RECT 1801.630 1020.180 1802.010 1020.190 ;
        RECT 1835.465 1020.490 1835.795 1020.505 ;
        RECT 1837.510 1020.490 1837.890 1020.500 ;
        RECT 1835.465 1020.190 1837.890 1020.490 ;
        RECT 1835.465 1020.175 1835.795 1020.190 ;
        RECT 1837.510 1020.180 1837.890 1020.190 ;
        RECT 2246.910 1020.490 2247.290 1020.500 ;
        RECT 2249.005 1020.490 2249.335 1020.505 ;
        RECT 2246.910 1020.190 2249.335 1020.490 ;
        RECT 2246.910 1020.180 2247.290 1020.190 ;
        RECT 2249.005 1020.175 2249.335 1020.190 ;
        RECT 2335.230 1020.490 2335.610 1020.500 ;
        RECT 2338.705 1020.490 2339.035 1020.505 ;
        RECT 2335.230 1020.190 2339.035 1020.490 ;
        RECT 2335.230 1020.180 2335.610 1020.190 ;
        RECT 2338.705 1020.175 2339.035 1020.190 ;
        RECT 2346.270 1020.490 2346.650 1020.500 ;
        RECT 2352.045 1020.490 2352.375 1020.505 ;
        RECT 2346.270 1020.190 2352.375 1020.490 ;
        RECT 2346.270 1020.180 2346.650 1020.190 ;
        RECT 2352.045 1020.175 2352.375 1020.190 ;
        RECT 2381.230 1020.490 2381.610 1020.500 ;
        RECT 2384.245 1020.490 2384.575 1020.505 ;
        RECT 2381.230 1020.190 2384.575 1020.490 ;
        RECT 2381.230 1020.180 2381.610 1020.190 ;
        RECT 2384.245 1020.175 2384.575 1020.190 ;
        RECT 2387.925 1020.490 2388.255 1020.505 ;
        RECT 2428.865 1020.500 2429.195 1020.505 ;
        RECT 2390.430 1020.490 2390.810 1020.500 ;
        RECT 2428.865 1020.490 2429.450 1020.500 ;
        RECT 2387.925 1020.190 2390.810 1020.490 ;
        RECT 2428.640 1020.190 2429.450 1020.490 ;
        RECT 2387.925 1020.175 2388.255 1020.190 ;
        RECT 2390.430 1020.180 2390.810 1020.190 ;
        RECT 2428.865 1020.180 2429.450 1020.190 ;
        RECT 2428.865 1020.175 2429.195 1020.180 ;
        RECT 1358.905 1019.810 1359.235 1019.825 ;
        RECT 1808.070 1019.810 1808.450 1019.820 ;
        RECT 1358.905 1019.510 1808.450 1019.810 ;
        RECT 1358.905 1019.495 1359.235 1019.510 ;
        RECT 1808.070 1019.500 1808.450 1019.510 ;
        RECT 1828.565 1019.810 1828.895 1019.825 ;
        RECT 1831.990 1019.810 1832.370 1019.820 ;
        RECT 1828.565 1019.510 1832.370 1019.810 ;
        RECT 1828.565 1019.495 1828.895 1019.510 ;
        RECT 1831.990 1019.500 1832.370 1019.510 ;
        RECT 2383.325 1019.810 2383.655 1019.825 ;
        RECT 2388.385 1019.810 2388.715 1019.825 ;
        RECT 2402.185 1019.820 2402.515 1019.825 ;
        RECT 2402.185 1019.810 2402.770 1019.820 ;
        RECT 2383.325 1019.510 2388.715 1019.810 ;
        RECT 2401.960 1019.510 2402.770 1019.810 ;
        RECT 2383.325 1019.495 2383.655 1019.510 ;
        RECT 2388.385 1019.495 2388.715 1019.510 ;
        RECT 2402.185 1019.500 2402.770 1019.510 ;
        RECT 2402.185 1019.495 2402.515 1019.500 ;
        RECT 1345.105 1019.130 1345.435 1019.145 ;
        RECT 1821.665 1019.140 1821.995 1019.145 ;
        RECT 1814.510 1019.130 1814.890 1019.140 ;
        RECT 1345.105 1018.830 1814.890 1019.130 ;
        RECT 1345.105 1018.815 1345.435 1018.830 ;
        RECT 1814.510 1018.820 1814.890 1018.830 ;
        RECT 1821.665 1019.130 1822.250 1019.140 ;
        RECT 2241.390 1019.130 2241.770 1019.140 ;
        RECT 2691.065 1019.130 2691.395 1019.145 ;
        RECT 1821.665 1018.830 1822.450 1019.130 ;
        RECT 2241.390 1018.830 2691.395 1019.130 ;
        RECT 1821.665 1018.820 1822.250 1018.830 ;
        RECT 2241.390 1018.820 2241.770 1018.830 ;
        RECT 1821.665 1018.815 1821.995 1018.820 ;
        RECT 2691.065 1018.815 2691.395 1018.830 ;
        RECT 1640.630 1018.450 1641.010 1018.460 ;
        RECT 1641.805 1018.450 1642.135 1018.465 ;
        RECT 1640.630 1018.150 1642.135 1018.450 ;
        RECT 1640.630 1018.140 1641.010 1018.150 ;
        RECT 1641.805 1018.135 1642.135 1018.150 ;
        RECT 1647.070 1018.450 1647.450 1018.460 ;
        RECT 1648.705 1018.450 1649.035 1018.465 ;
        RECT 1647.070 1018.150 1649.035 1018.450 ;
        RECT 1647.070 1018.140 1647.450 1018.150 ;
        RECT 1648.705 1018.135 1649.035 1018.150 ;
        RECT 1653.510 1018.450 1653.890 1018.460 ;
        RECT 1655.605 1018.450 1655.935 1018.465 ;
        RECT 1653.510 1018.150 1655.935 1018.450 ;
        RECT 1653.510 1018.140 1653.890 1018.150 ;
        RECT 1655.605 1018.135 1655.935 1018.150 ;
        RECT 1670.325 1018.450 1670.655 1018.465 ;
        RECT 1674.670 1018.450 1675.050 1018.460 ;
        RECT 1670.325 1018.150 1675.050 1018.450 ;
        RECT 1670.325 1018.135 1670.655 1018.150 ;
        RECT 1674.670 1018.140 1675.050 1018.150 ;
        RECT 1711.265 1018.450 1711.595 1018.465 ;
        RECT 1714.230 1018.450 1714.610 1018.460 ;
        RECT 1711.265 1018.150 1714.610 1018.450 ;
        RECT 1711.265 1018.135 1711.595 1018.150 ;
        RECT 1714.230 1018.140 1714.610 1018.150 ;
        RECT 1718.165 1018.450 1718.495 1018.465 ;
        RECT 1745.765 1018.460 1746.095 1018.465 ;
        RECT 1719.750 1018.450 1720.130 1018.460 ;
        RECT 1718.165 1018.150 1720.130 1018.450 ;
        RECT 1718.165 1018.135 1718.495 1018.150 ;
        RECT 1719.750 1018.140 1720.130 1018.150 ;
        RECT 1745.510 1018.450 1746.095 1018.460 ;
        RECT 1755.425 1018.460 1755.755 1018.465 ;
        RECT 1755.425 1018.450 1756.010 1018.460 ;
        RECT 1745.510 1018.150 1746.320 1018.450 ;
        RECT 1755.200 1018.150 1756.010 1018.450 ;
        RECT 1745.510 1018.140 1746.095 1018.150 ;
        RECT 1745.765 1018.135 1746.095 1018.140 ;
        RECT 1755.425 1018.140 1756.010 1018.150 ;
        RECT 1759.105 1018.450 1759.435 1018.465 ;
        RECT 2415.065 1018.460 2415.395 1018.465 ;
        RECT 2415.065 1018.450 2415.650 1018.460 ;
        RECT 2437.350 1018.450 2437.730 1018.460 ;
        RECT 1759.105 1018.150 2413.770 1018.450 ;
        RECT 2414.840 1018.150 2415.650 1018.450 ;
        RECT 1755.425 1018.135 1755.755 1018.140 ;
        RECT 1759.105 1018.135 1759.435 1018.150 ;
        RECT 1675.845 1017.770 1676.175 1017.785 ;
        RECT 1697.925 1017.770 1698.255 1017.785 ;
        RECT 1704.365 1017.780 1704.695 1017.785 ;
        RECT 1700.430 1017.770 1700.810 1017.780 ;
        RECT 1675.845 1017.470 1700.810 1017.770 ;
        RECT 1675.845 1017.455 1676.175 1017.470 ;
        RECT 1697.925 1017.455 1698.255 1017.470 ;
        RECT 1700.430 1017.460 1700.810 1017.470 ;
        RECT 1704.110 1017.770 1704.695 1017.780 ;
        RECT 1745.305 1017.770 1745.635 1017.785 ;
        RECT 2413.470 1017.770 2413.770 1018.150 ;
        RECT 2415.065 1018.140 2415.650 1018.150 ;
        RECT 2416.230 1018.150 2437.730 1018.450 ;
        RECT 2415.065 1018.135 2415.395 1018.140 ;
        RECT 2416.230 1017.770 2416.530 1018.150 ;
        RECT 2437.350 1018.140 2437.730 1018.150 ;
        RECT 2421.965 1017.780 2422.295 1017.785 ;
        RECT 1704.110 1017.470 1704.920 1017.770 ;
        RECT 1745.305 1017.470 2412.850 1017.770 ;
        RECT 2413.470 1017.470 2416.530 1017.770 ;
        RECT 2421.710 1017.770 2422.295 1017.780 ;
        RECT 2442.870 1017.770 2443.250 1017.780 ;
        RECT 2421.710 1017.470 2422.520 1017.770 ;
        RECT 2422.970 1017.470 2443.250 1017.770 ;
        RECT 1704.110 1017.460 1704.695 1017.470 ;
        RECT 1704.365 1017.455 1704.695 1017.460 ;
        RECT 1745.305 1017.455 1745.635 1017.470 ;
        RECT 1641.805 1017.100 1642.135 1017.105 ;
        RECT 1662.045 1017.100 1662.375 1017.105 ;
        RECT 1641.550 1017.090 1642.135 1017.100 ;
        RECT 1661.790 1017.090 1662.375 1017.100 ;
        RECT 1664.550 1017.090 1664.930 1017.100 ;
        RECT 1669.405 1017.090 1669.735 1017.105 ;
        RECT 1683.205 1017.100 1683.535 1017.105 ;
        RECT 1641.550 1016.790 1642.360 1017.090 ;
        RECT 1661.790 1016.790 1662.600 1017.090 ;
        RECT 1664.550 1016.790 1669.735 1017.090 ;
        RECT 1641.550 1016.780 1642.135 1016.790 ;
        RECT 1661.790 1016.780 1662.375 1016.790 ;
        RECT 1664.550 1016.780 1664.930 1016.790 ;
        RECT 1641.805 1016.775 1642.135 1016.780 ;
        RECT 1662.045 1016.775 1662.375 1016.780 ;
        RECT 1669.405 1016.775 1669.735 1016.790 ;
        RECT 1682.950 1017.090 1683.535 1017.100 ;
        RECT 1690.565 1017.090 1690.895 1017.105 ;
        RECT 1787.165 1017.100 1787.495 1017.105 ;
        RECT 1691.230 1017.090 1691.610 1017.100 ;
        RECT 1682.950 1016.790 1683.760 1017.090 ;
        RECT 1690.565 1016.790 1691.610 1017.090 ;
        RECT 1682.950 1016.780 1683.535 1016.790 ;
        RECT 1683.205 1016.775 1683.535 1016.780 ;
        RECT 1690.565 1016.775 1690.895 1016.790 ;
        RECT 1691.230 1016.780 1691.610 1016.790 ;
        RECT 1786.910 1017.090 1787.495 1017.100 ;
        RECT 2245.785 1017.090 2246.115 1017.105 ;
        RECT 2247.830 1017.090 2248.210 1017.100 ;
        RECT 1786.910 1016.790 1787.720 1017.090 ;
        RECT 2245.785 1016.790 2248.210 1017.090 ;
        RECT 1786.910 1016.780 1787.495 1016.790 ;
        RECT 1787.165 1016.775 1787.495 1016.780 ;
        RECT 2245.785 1016.775 2246.115 1016.790 ;
        RECT 2247.830 1016.780 2248.210 1016.790 ;
        RECT 2252.685 1017.090 2253.015 1017.105 ;
        RECT 2254.270 1017.090 2254.650 1017.100 ;
        RECT 2252.685 1016.790 2254.650 1017.090 ;
        RECT 2252.685 1016.775 2253.015 1016.790 ;
        RECT 2254.270 1016.780 2254.650 1016.790 ;
        RECT 2259.585 1017.090 2259.915 1017.105 ;
        RECT 2266.485 1017.100 2266.815 1017.105 ;
        RECT 2260.710 1017.090 2261.090 1017.100 ;
        RECT 2259.585 1016.790 2261.090 1017.090 ;
        RECT 2259.585 1016.775 2259.915 1016.790 ;
        RECT 2260.710 1016.780 2261.090 1016.790 ;
        RECT 2266.230 1017.090 2266.815 1017.100 ;
        RECT 2280.030 1017.090 2280.410 1017.100 ;
        RECT 2280.745 1017.090 2281.075 1017.105 ;
        RECT 2266.230 1016.790 2267.040 1017.090 ;
        RECT 2280.030 1016.790 2281.075 1017.090 ;
        RECT 2266.230 1016.780 2266.815 1016.790 ;
        RECT 2280.030 1016.780 2280.410 1016.790 ;
        RECT 2266.485 1016.775 2266.815 1016.780 ;
        RECT 2280.745 1016.775 2281.075 1016.790 ;
        RECT 2293.830 1017.090 2294.210 1017.100 ;
        RECT 2297.305 1017.090 2297.635 1017.105 ;
        RECT 2293.830 1016.790 2297.635 1017.090 ;
        RECT 2293.830 1016.780 2294.210 1016.790 ;
        RECT 2297.305 1016.775 2297.635 1016.790 ;
        RECT 2304.870 1017.090 2305.250 1017.100 ;
        RECT 2310.645 1017.090 2310.975 1017.105 ;
        RECT 2304.870 1016.790 2310.975 1017.090 ;
        RECT 2304.870 1016.780 2305.250 1016.790 ;
        RECT 2310.645 1016.775 2310.975 1016.790 ;
        RECT 2311.310 1017.090 2311.690 1017.100 ;
        RECT 2317.545 1017.090 2317.875 1017.105 ;
        RECT 2311.310 1016.790 2317.875 1017.090 ;
        RECT 2311.310 1016.780 2311.690 1016.790 ;
        RECT 2317.545 1016.775 2317.875 1016.790 ;
        RECT 2387.925 1017.090 2388.255 1017.105 ;
        RECT 2393.190 1017.090 2393.570 1017.100 ;
        RECT 2387.925 1016.790 2393.570 1017.090 ;
        RECT 2387.925 1016.775 2388.255 1016.790 ;
        RECT 2393.190 1016.780 2393.570 1016.790 ;
        RECT 1655.605 1016.420 1655.935 1016.425 ;
        RECT 1655.350 1016.410 1655.935 1016.420 ;
        RECT 1658.110 1016.410 1658.490 1016.420 ;
        RECT 1662.505 1016.410 1662.835 1016.425 ;
        RECT 1669.865 1016.420 1670.195 1016.425 ;
        RECT 1669.865 1016.410 1670.450 1016.420 ;
        RECT 1655.350 1016.110 1656.160 1016.410 ;
        RECT 1658.110 1016.110 1662.835 1016.410 ;
        RECT 1669.640 1016.110 1670.450 1016.410 ;
        RECT 1655.350 1016.100 1655.935 1016.110 ;
        RECT 1658.110 1016.100 1658.490 1016.110 ;
        RECT 1655.605 1016.095 1655.935 1016.100 ;
        RECT 1662.505 1016.095 1662.835 1016.110 ;
        RECT 1669.865 1016.100 1670.450 1016.110 ;
        RECT 1676.765 1016.410 1677.095 1016.425 ;
        RECT 1681.110 1016.410 1681.490 1016.420 ;
        RECT 1676.765 1016.110 1681.490 1016.410 ;
        RECT 1669.865 1016.095 1670.195 1016.100 ;
        RECT 1676.765 1016.095 1677.095 1016.110 ;
        RECT 1681.110 1016.100 1681.490 1016.110 ;
        RECT 1683.665 1016.410 1683.995 1016.425 ;
        RECT 1697.465 1016.420 1697.795 1016.425 ;
        RECT 1684.790 1016.410 1685.170 1016.420 ;
        RECT 1697.465 1016.410 1698.050 1016.420 ;
        RECT 1683.665 1016.110 1685.170 1016.410 ;
        RECT 1697.240 1016.110 1698.050 1016.410 ;
        RECT 1683.665 1016.095 1683.995 1016.110 ;
        RECT 1684.790 1016.100 1685.170 1016.110 ;
        RECT 1697.465 1016.100 1698.050 1016.110 ;
        RECT 1725.065 1016.410 1725.395 1016.425 ;
        RECT 1726.190 1016.410 1726.570 1016.420 ;
        RECT 1725.065 1016.110 1726.570 1016.410 ;
        RECT 1697.465 1016.095 1697.795 1016.100 ;
        RECT 1725.065 1016.095 1725.395 1016.110 ;
        RECT 1726.190 1016.100 1726.570 1016.110 ;
        RECT 1745.765 1016.410 1746.095 1016.425 ;
        RECT 1749.190 1016.410 1749.570 1016.420 ;
        RECT 1745.765 1016.110 1749.570 1016.410 ;
        RECT 1745.765 1016.095 1746.095 1016.110 ;
        RECT 1749.190 1016.100 1749.570 1016.110 ;
        RECT 1842.365 1016.410 1842.695 1016.425 ;
        RECT 1843.030 1016.410 1843.410 1016.420 ;
        RECT 1842.365 1016.110 1843.410 1016.410 ;
        RECT 1842.365 1016.095 1842.695 1016.110 ;
        RECT 1843.030 1016.100 1843.410 1016.110 ;
        RECT 2253.350 1016.410 2253.730 1016.420 ;
        RECT 2255.905 1016.410 2256.235 1016.425 ;
        RECT 2253.350 1016.110 2256.235 1016.410 ;
        RECT 2253.350 1016.100 2253.730 1016.110 ;
        RECT 2255.905 1016.095 2256.235 1016.110 ;
        RECT 2264.390 1016.410 2264.770 1016.420 ;
        RECT 2269.705 1016.410 2270.035 1016.425 ;
        RECT 2264.390 1016.110 2270.035 1016.410 ;
        RECT 2264.390 1016.100 2264.770 1016.110 ;
        RECT 2269.705 1016.095 2270.035 1016.110 ;
        RECT 2273.385 1016.410 2273.715 1016.425 ;
        RECT 2274.510 1016.410 2274.890 1016.420 ;
        RECT 2275.225 1016.410 2275.555 1016.425 ;
        RECT 2276.145 1016.420 2276.475 1016.425 ;
        RECT 2276.145 1016.410 2276.730 1016.420 ;
        RECT 2273.385 1016.110 2275.555 1016.410 ;
        RECT 2275.920 1016.110 2276.730 1016.410 ;
        RECT 2273.385 1016.095 2273.715 1016.110 ;
        RECT 2274.510 1016.100 2274.890 1016.110 ;
        RECT 2275.225 1016.095 2275.555 1016.110 ;
        RECT 2276.145 1016.100 2276.730 1016.110 ;
        RECT 2287.390 1016.410 2287.770 1016.420 ;
        RECT 2290.405 1016.410 2290.735 1016.425 ;
        RECT 2287.390 1016.110 2290.735 1016.410 ;
        RECT 2287.390 1016.100 2287.770 1016.110 ;
        RECT 2276.145 1016.095 2276.475 1016.100 ;
        RECT 2290.405 1016.095 2290.735 1016.110 ;
        RECT 2300.270 1016.410 2300.650 1016.420 ;
        RECT 2304.205 1016.410 2304.535 1016.425 ;
        RECT 2300.270 1016.110 2304.535 1016.410 ;
        RECT 2300.270 1016.100 2300.650 1016.110 ;
        RECT 2304.205 1016.095 2304.535 1016.110 ;
        RECT 2315.910 1016.410 2316.290 1016.420 ;
        RECT 2318.005 1016.410 2318.335 1016.425 ;
        RECT 2315.910 1016.110 2318.335 1016.410 ;
        RECT 2315.910 1016.100 2316.290 1016.110 ;
        RECT 2318.005 1016.095 2318.335 1016.110 ;
        RECT 2323.065 1016.420 2323.395 1016.425 ;
        RECT 2323.065 1016.410 2323.650 1016.420 ;
        RECT 2325.365 1016.410 2325.695 1016.425 ;
        RECT 2329.710 1016.410 2330.090 1016.420 ;
        RECT 2332.725 1016.410 2333.055 1016.425 ;
        RECT 2323.065 1016.110 2323.850 1016.410 ;
        RECT 2325.365 1016.110 2333.055 1016.410 ;
        RECT 2323.065 1016.100 2323.650 1016.110 ;
        RECT 2323.065 1016.095 2323.395 1016.100 ;
        RECT 2325.365 1016.095 2325.695 1016.110 ;
        RECT 2329.710 1016.100 2330.090 1016.110 ;
        RECT 2332.725 1016.095 2333.055 1016.110 ;
        RECT 2358.230 1016.410 2358.610 1016.420 ;
        RECT 2359.405 1016.410 2359.735 1016.425 ;
        RECT 2358.230 1016.110 2359.735 1016.410 ;
        RECT 2358.230 1016.100 2358.610 1016.110 ;
        RECT 2359.405 1016.095 2359.735 1016.110 ;
        RECT 2363.750 1016.410 2364.130 1016.420 ;
        RECT 2366.305 1016.410 2366.635 1016.425 ;
        RECT 2363.750 1016.110 2366.635 1016.410 ;
        RECT 2363.750 1016.100 2364.130 1016.110 ;
        RECT 2366.305 1016.095 2366.635 1016.110 ;
        RECT 2375.710 1016.410 2376.090 1016.420 ;
        RECT 2380.105 1016.410 2380.435 1016.425 ;
        RECT 2375.710 1016.110 2380.435 1016.410 ;
        RECT 2375.710 1016.100 2376.090 1016.110 ;
        RECT 2380.105 1016.095 2380.435 1016.110 ;
        RECT 2387.465 1016.410 2387.795 1016.425 ;
        RECT 2388.590 1016.410 2388.970 1016.420 ;
        RECT 2387.465 1016.110 2388.970 1016.410 ;
        RECT 2412.550 1016.410 2412.850 1017.470 ;
        RECT 2421.710 1017.460 2422.295 1017.470 ;
        RECT 2421.965 1017.455 2422.295 1017.460 ;
        RECT 2422.970 1016.410 2423.270 1017.470 ;
        RECT 2442.870 1017.460 2443.250 1017.470 ;
        RECT 2412.550 1016.110 2423.270 1016.410 ;
        RECT 2428.865 1016.410 2429.195 1016.425 ;
        RECT 2431.830 1016.410 2432.210 1016.420 ;
        RECT 2428.865 1016.110 2432.210 1016.410 ;
        RECT 2387.465 1016.095 2387.795 1016.110 ;
        RECT 2388.590 1016.100 2388.970 1016.110 ;
        RECT 2428.865 1016.095 2429.195 1016.110 ;
        RECT 2431.830 1016.100 2432.210 1016.110 ;
        RECT 1647.990 1015.730 1648.370 1015.740 ;
        RECT 1648.705 1015.730 1649.035 1015.745 ;
        RECT 1647.990 1015.430 1649.035 1015.730 ;
        RECT 1647.990 1015.420 1648.370 1015.430 ;
        RECT 1648.705 1015.415 1649.035 1015.430 ;
        RECT 1668.230 1015.730 1668.610 1015.740 ;
        RECT 1669.405 1015.730 1669.735 1015.745 ;
        RECT 1668.230 1015.430 1669.735 1015.730 ;
        RECT 1668.230 1015.420 1668.610 1015.430 ;
        RECT 1669.405 1015.415 1669.735 1015.430 ;
        RECT 1673.750 1015.730 1674.130 1015.740 ;
        RECT 1676.305 1015.730 1676.635 1015.745 ;
        RECT 1673.750 1015.430 1676.635 1015.730 ;
        RECT 1673.750 1015.420 1674.130 1015.430 ;
        RECT 1676.305 1015.415 1676.635 1015.430 ;
        RECT 1708.710 1015.730 1709.090 1015.740 ;
        RECT 1710.805 1015.730 1711.135 1015.745 ;
        RECT 1708.710 1015.430 1711.135 1015.730 ;
        RECT 1708.710 1015.420 1709.090 1015.430 ;
        RECT 1710.805 1015.415 1711.135 1015.430 ;
        RECT 1731.965 1015.730 1732.295 1015.745 ;
        RECT 1738.865 1015.740 1739.195 1015.745 ;
        RECT 1732.630 1015.730 1733.010 1015.740 ;
        RECT 1738.865 1015.730 1739.450 1015.740 ;
        RECT 1731.965 1015.430 1733.010 1015.730 ;
        RECT 1738.640 1015.430 1739.450 1015.730 ;
        RECT 1731.965 1015.415 1732.295 1015.430 ;
        RECT 1732.630 1015.420 1733.010 1015.430 ;
        RECT 1738.865 1015.420 1739.450 1015.430 ;
        RECT 1759.565 1015.730 1759.895 1015.745 ;
        RECT 1766.005 1015.740 1766.335 1015.745 ;
        RECT 1763.910 1015.730 1764.290 1015.740 ;
        RECT 1765.750 1015.730 1766.335 1015.740 ;
        RECT 1759.565 1015.430 1764.290 1015.730 ;
        RECT 1765.550 1015.430 1766.335 1015.730 ;
        RECT 1738.865 1015.415 1739.195 1015.420 ;
        RECT 1759.565 1015.415 1759.895 1015.430 ;
        RECT 1763.910 1015.420 1764.290 1015.430 ;
        RECT 1765.750 1015.420 1766.335 1015.430 ;
        RECT 1766.005 1015.415 1766.335 1015.420 ;
        RECT 1773.365 1015.730 1773.695 1015.745 ;
        RECT 1780.265 1015.740 1780.595 1015.745 ;
        RECT 1789.005 1015.740 1789.335 1015.745 ;
        RECT 1774.030 1015.730 1774.410 1015.740 ;
        RECT 1780.265 1015.730 1780.850 1015.740 ;
        RECT 1788.750 1015.730 1789.335 1015.740 ;
        RECT 1773.365 1015.430 1774.410 1015.730 ;
        RECT 1780.040 1015.430 1780.850 1015.730 ;
        RECT 1788.550 1015.430 1789.335 1015.730 ;
        RECT 1773.365 1015.415 1773.695 1015.430 ;
        RECT 1774.030 1015.420 1774.410 1015.430 ;
        RECT 1780.265 1015.420 1780.850 1015.430 ;
        RECT 1788.750 1015.420 1789.335 1015.430 ;
        RECT 1780.265 1015.415 1780.595 1015.420 ;
        RECT 1789.005 1015.415 1789.335 1015.420 ;
        RECT 1680.190 1015.050 1680.570 1015.060 ;
        RECT 1683.205 1015.050 1683.535 1015.065 ;
        RECT 1689.645 1015.060 1689.975 1015.065 ;
        RECT 1696.085 1015.060 1696.415 1015.065 ;
        RECT 1689.390 1015.050 1689.975 1015.060 ;
        RECT 1695.830 1015.050 1696.415 1015.060 ;
        RECT 1711.265 1015.060 1711.595 1015.065 ;
        RECT 1712.185 1015.060 1712.515 1015.065 ;
        RECT 1718.165 1015.060 1718.495 1015.065 ;
        RECT 1724.605 1015.060 1724.935 1015.065 ;
        RECT 1711.265 1015.050 1711.850 1015.060 ;
        RECT 1680.190 1014.750 1683.535 1015.050 ;
        RECT 1689.190 1014.750 1689.975 1015.050 ;
        RECT 1695.630 1014.750 1696.415 1015.050 ;
        RECT 1711.040 1014.750 1711.850 1015.050 ;
        RECT 1680.190 1014.740 1680.570 1014.750 ;
        RECT 1683.205 1014.735 1683.535 1014.750 ;
        RECT 1689.390 1014.740 1689.975 1014.750 ;
        RECT 1695.830 1014.740 1696.415 1014.750 ;
        RECT 1689.645 1014.735 1689.975 1014.740 ;
        RECT 1696.085 1014.735 1696.415 1014.740 ;
        RECT 1711.265 1014.740 1711.850 1014.750 ;
        RECT 1712.185 1015.050 1712.770 1015.060 ;
        RECT 1717.910 1015.050 1718.495 1015.060 ;
        RECT 1724.350 1015.050 1724.935 1015.060 ;
        RECT 1712.185 1014.750 1712.970 1015.050 ;
        RECT 1717.710 1014.750 1718.495 1015.050 ;
        RECT 1724.150 1014.750 1724.935 1015.050 ;
        RECT 1712.185 1014.740 1712.770 1014.750 ;
        RECT 1717.910 1014.740 1718.495 1014.750 ;
        RECT 1724.350 1014.740 1724.935 1014.750 ;
        RECT 1711.265 1014.735 1711.595 1014.740 ;
        RECT 1712.185 1014.735 1712.515 1014.740 ;
        RECT 1718.165 1014.735 1718.495 1014.740 ;
        RECT 1724.605 1014.735 1724.935 1014.740 ;
        RECT 1729.665 1015.060 1729.995 1015.065 ;
        RECT 1735.645 1015.060 1735.975 1015.065 ;
        RECT 1729.665 1015.050 1730.250 1015.060 ;
        RECT 1735.390 1015.050 1735.975 1015.060 ;
        RECT 1729.665 1014.750 1730.450 1015.050 ;
        RECT 1735.190 1014.750 1735.975 1015.050 ;
        RECT 1729.665 1014.740 1730.250 1014.750 ;
        RECT 1735.390 1014.740 1735.975 1014.750 ;
        RECT 1729.665 1014.735 1729.995 1014.740 ;
        RECT 1735.645 1014.735 1735.975 1014.740 ;
        RECT 1741.625 1015.060 1741.955 1015.065 ;
        RECT 1741.625 1015.050 1742.210 1015.060 ;
        RECT 1746.225 1015.050 1746.555 1015.065 ;
        RECT 1754.965 1015.060 1755.295 1015.065 ;
        RECT 1758.645 1015.060 1758.975 1015.065 ;
        RECT 1748.270 1015.050 1748.650 1015.060 ;
        RECT 1754.710 1015.050 1755.295 1015.060 ;
        RECT 1758.390 1015.050 1758.975 1015.060 ;
        RECT 1766.465 1015.060 1766.795 1015.065 ;
        RECT 1771.525 1015.060 1771.855 1015.065 ;
        RECT 1777.965 1015.060 1778.295 1015.065 ;
        RECT 1766.465 1015.050 1767.050 1015.060 ;
        RECT 1771.270 1015.050 1771.855 1015.060 ;
        RECT 1777.710 1015.050 1778.295 1015.060 ;
        RECT 1741.625 1014.750 1742.410 1015.050 ;
        RECT 1746.225 1014.750 1748.650 1015.050 ;
        RECT 1754.510 1014.750 1755.295 1015.050 ;
        RECT 1758.190 1014.750 1758.975 1015.050 ;
        RECT 1766.240 1014.750 1767.050 1015.050 ;
        RECT 1771.070 1014.750 1771.855 1015.050 ;
        RECT 1777.510 1014.750 1778.295 1015.050 ;
        RECT 1741.625 1014.740 1742.210 1014.750 ;
        RECT 1741.625 1014.735 1741.955 1014.740 ;
        RECT 1746.225 1014.735 1746.555 1014.750 ;
        RECT 1748.270 1014.740 1748.650 1014.750 ;
        RECT 1754.710 1014.740 1755.295 1014.750 ;
        RECT 1758.390 1014.740 1758.975 1014.750 ;
        RECT 1754.965 1014.735 1755.295 1014.740 ;
        RECT 1758.645 1014.735 1758.975 1014.740 ;
        RECT 1766.465 1014.740 1767.050 1014.750 ;
        RECT 1771.270 1014.740 1771.855 1014.750 ;
        RECT 1777.710 1014.740 1778.295 1014.750 ;
        RECT 1766.465 1014.735 1766.795 1014.740 ;
        RECT 1771.525 1014.735 1771.855 1014.740 ;
        RECT 1777.965 1014.735 1778.295 1014.740 ;
        RECT 1782.105 1015.060 1782.435 1015.065 ;
        RECT 1782.105 1015.050 1782.690 1015.060 ;
        RECT 1787.165 1015.050 1787.495 1015.065 ;
        RECT 1793.145 1015.060 1793.475 1015.065 ;
        RECT 1800.045 1015.060 1800.375 1015.065 ;
        RECT 1806.485 1015.060 1806.815 1015.065 ;
        RECT 1789.670 1015.050 1790.050 1015.060 ;
        RECT 1782.105 1014.750 1782.890 1015.050 ;
        RECT 1787.165 1014.750 1790.050 1015.050 ;
        RECT 1782.105 1014.740 1782.690 1014.750 ;
        RECT 1782.105 1014.735 1782.435 1014.740 ;
        RECT 1787.165 1014.735 1787.495 1014.750 ;
        RECT 1789.670 1014.740 1790.050 1014.750 ;
        RECT 1793.145 1015.050 1793.730 1015.060 ;
        RECT 1799.790 1015.050 1800.375 1015.060 ;
        RECT 1806.230 1015.050 1806.815 1015.060 ;
        RECT 1793.145 1014.750 1793.930 1015.050 ;
        RECT 1799.590 1014.750 1800.375 1015.050 ;
        RECT 1806.030 1014.750 1806.815 1015.050 ;
        RECT 1793.145 1014.740 1793.730 1014.750 ;
        RECT 1799.790 1014.740 1800.375 1014.750 ;
        RECT 1806.230 1014.740 1806.815 1014.750 ;
        RECT 1793.145 1014.735 1793.475 1014.740 ;
        RECT 1800.045 1014.735 1800.375 1014.740 ;
        RECT 1806.485 1014.735 1806.815 1014.740 ;
        RECT 1812.465 1015.060 1812.795 1015.065 ;
        RECT 1817.525 1015.060 1817.855 1015.065 ;
        RECT 1812.465 1015.050 1813.050 1015.060 ;
        RECT 1817.270 1015.050 1817.855 1015.060 ;
        RECT 1812.465 1014.750 1813.250 1015.050 ;
        RECT 1817.070 1014.750 1817.855 1015.050 ;
        RECT 1812.465 1014.740 1813.050 1014.750 ;
        RECT 1817.270 1014.740 1817.855 1014.750 ;
        RECT 1812.465 1014.735 1812.795 1014.740 ;
        RECT 1817.525 1014.735 1817.855 1014.740 ;
        RECT 1823.505 1015.060 1823.835 1015.065 ;
        RECT 1823.505 1015.050 1824.090 1015.060 ;
        RECT 2258.870 1015.050 2259.250 1015.060 ;
        RECT 2262.805 1015.050 2263.135 1015.065 ;
        RECT 1823.505 1014.750 1824.290 1015.050 ;
        RECT 2258.870 1014.750 2263.135 1015.050 ;
        RECT 1823.505 1014.740 1824.090 1014.750 ;
        RECT 2258.870 1014.740 2259.250 1014.750 ;
        RECT 1823.505 1014.735 1823.835 1014.740 ;
        RECT 2262.805 1014.735 2263.135 1014.750 ;
        RECT 2270.830 1015.050 2271.210 1015.060 ;
        RECT 2276.605 1015.050 2276.935 1015.065 ;
        RECT 2270.830 1014.750 2276.935 1015.050 ;
        RECT 2270.830 1014.740 2271.210 1014.750 ;
        RECT 2276.605 1014.735 2276.935 1014.750 ;
        RECT 2281.870 1015.050 2282.250 1015.060 ;
        RECT 2283.045 1015.050 2283.375 1015.065 ;
        RECT 2281.870 1014.750 2283.375 1015.050 ;
        RECT 2281.870 1014.740 2282.250 1014.750 ;
        RECT 2283.045 1014.735 2283.375 1014.750 ;
        RECT 2289.230 1015.050 2289.610 1015.060 ;
        RECT 2289.945 1015.050 2290.275 1015.065 ;
        RECT 2295.005 1015.060 2295.335 1015.065 ;
        RECT 2294.750 1015.050 2295.335 1015.060 ;
        RECT 2289.230 1014.750 2290.275 1015.050 ;
        RECT 2294.550 1014.750 2295.335 1015.050 ;
        RECT 2289.230 1014.740 2289.610 1014.750 ;
        RECT 2289.945 1014.735 2290.275 1014.750 ;
        RECT 2294.750 1014.740 2295.335 1014.750 ;
        RECT 2302.110 1015.050 2302.490 1015.060 ;
        RECT 2302.825 1015.050 2303.155 1015.065 ;
        RECT 2302.110 1014.750 2303.155 1015.050 ;
        RECT 2302.110 1014.740 2302.490 1014.750 ;
        RECT 2295.005 1014.735 2295.335 1014.740 ;
        RECT 2302.825 1014.735 2303.155 1014.750 ;
        RECT 2306.965 1015.050 2307.295 1015.065 ;
        RECT 2312.025 1015.060 2312.355 1015.065 ;
        RECT 2318.005 1015.060 2318.335 1015.065 ;
        RECT 2307.630 1015.050 2308.010 1015.060 ;
        RECT 2306.965 1014.750 2308.010 1015.050 ;
        RECT 2306.965 1014.735 2307.295 1014.750 ;
        RECT 2307.630 1014.740 2308.010 1014.750 ;
        RECT 2312.025 1015.050 2312.610 1015.060 ;
        RECT 2317.750 1015.050 2318.335 1015.060 ;
        RECT 2312.025 1014.750 2312.810 1015.050 ;
        RECT 2317.550 1014.750 2318.335 1015.050 ;
        RECT 2312.025 1014.740 2312.610 1014.750 ;
        RECT 2317.750 1014.740 2318.335 1014.750 ;
        RECT 2322.350 1015.050 2322.730 1015.060 ;
        RECT 2324.905 1015.050 2325.235 1015.065 ;
        RECT 2322.350 1014.750 2325.235 1015.050 ;
        RECT 2322.350 1014.740 2322.730 1014.750 ;
        RECT 2312.025 1014.735 2312.355 1014.740 ;
        RECT 2318.005 1014.735 2318.335 1014.740 ;
        RECT 2324.905 1014.735 2325.235 1014.750 ;
        RECT 2328.790 1015.050 2329.170 1015.060 ;
        RECT 2331.805 1015.050 2332.135 1015.065 ;
        RECT 2336.405 1015.060 2336.735 1015.065 ;
        RECT 2336.150 1015.050 2336.735 1015.060 ;
        RECT 2328.790 1014.750 2332.135 1015.050 ;
        RECT 2335.950 1014.750 2336.735 1015.050 ;
        RECT 2328.790 1014.740 2329.170 1014.750 ;
        RECT 2331.805 1014.735 2332.135 1014.750 ;
        RECT 2336.150 1014.740 2336.735 1014.750 ;
        RECT 2336.405 1014.735 2336.735 1014.740 ;
        RECT 2342.385 1015.060 2342.715 1015.065 ;
        RECT 2346.985 1015.060 2347.315 1015.065 ;
        RECT 2353.425 1015.060 2353.755 1015.065 ;
        RECT 2342.385 1015.050 2342.970 1015.060 ;
        RECT 2346.985 1015.050 2347.570 1015.060 ;
        RECT 2353.425 1015.050 2354.010 1015.060 ;
        RECT 2358.025 1015.050 2358.355 1015.065 ;
        RECT 2342.385 1014.750 2343.170 1015.050 ;
        RECT 2346.985 1014.750 2347.770 1015.050 ;
        RECT 2353.425 1014.750 2358.355 1015.050 ;
        RECT 2342.385 1014.740 2342.970 1014.750 ;
        RECT 2346.985 1014.740 2347.570 1014.750 ;
        RECT 2353.425 1014.740 2354.010 1014.750 ;
        RECT 2342.385 1014.735 2342.715 1014.740 ;
        RECT 2346.985 1014.735 2347.315 1014.740 ;
        RECT 2353.425 1014.735 2353.755 1014.740 ;
        RECT 2358.025 1014.735 2358.355 1014.750 ;
        RECT 2358.945 1015.060 2359.275 1015.065 ;
        RECT 2364.465 1015.060 2364.795 1015.065 ;
        RECT 2370.905 1015.060 2371.235 1015.065 ;
        RECT 2377.805 1015.060 2378.135 1015.065 ;
        RECT 2358.945 1015.050 2359.530 1015.060 ;
        RECT 2364.465 1015.050 2365.050 1015.060 ;
        RECT 2370.905 1015.050 2371.490 1015.060 ;
        RECT 2377.550 1015.050 2378.135 1015.060 ;
        RECT 2358.945 1014.750 2359.730 1015.050 ;
        RECT 2364.465 1014.750 2365.250 1015.050 ;
        RECT 2370.905 1014.750 2371.690 1015.050 ;
        RECT 2377.350 1014.750 2378.135 1015.050 ;
        RECT 2358.945 1014.740 2359.530 1014.750 ;
        RECT 2364.465 1014.740 2365.050 1014.750 ;
        RECT 2370.905 1014.740 2371.490 1014.750 ;
        RECT 2377.550 1014.740 2378.135 1014.750 ;
        RECT 2358.945 1014.735 2359.275 1014.740 ;
        RECT 2364.465 1014.735 2364.795 1014.740 ;
        RECT 2370.905 1014.735 2371.235 1014.740 ;
        RECT 2377.805 1014.735 2378.135 1014.740 ;
        RECT 2380.565 1015.050 2380.895 1015.065 ;
        RECT 2382.150 1015.050 2382.530 1015.060 ;
        RECT 2380.565 1014.750 2382.530 1015.050 ;
        RECT 2380.565 1014.735 2380.895 1014.750 ;
        RECT 2382.150 1014.740 2382.530 1014.750 ;
        RECT 2394.365 1015.050 2394.695 1015.065 ;
        RECT 2399.630 1015.050 2400.010 1015.060 ;
        RECT 2394.365 1014.750 2400.010 1015.050 ;
        RECT 2394.365 1014.735 2394.695 1014.750 ;
        RECT 2399.630 1014.740 2400.010 1014.750 ;
        RECT 2403.105 1015.050 2403.435 1015.065 ;
        RECT 2406.070 1015.050 2406.450 1015.060 ;
        RECT 2403.105 1014.750 2406.450 1015.050 ;
        RECT 2403.105 1014.735 2403.435 1014.750 ;
        RECT 2406.070 1014.740 2406.450 1014.750 ;
        RECT 2408.165 1015.050 2408.495 1015.065 ;
        RECT 2410.670 1015.050 2411.050 1015.060 ;
        RECT 2408.165 1014.750 2411.050 1015.050 ;
        RECT 2408.165 1014.735 2408.495 1014.750 ;
        RECT 2410.670 1014.740 2411.050 1014.750 ;
        RECT 2415.065 1015.050 2415.395 1015.065 ;
        RECT 2417.110 1015.050 2417.490 1015.060 ;
        RECT 2415.065 1014.750 2417.490 1015.050 ;
        RECT 2415.065 1014.735 2415.395 1014.750 ;
        RECT 2417.110 1014.740 2417.490 1014.750 ;
        RECT 2421.965 1015.050 2422.295 1015.065 ;
        RECT 2423.550 1015.050 2423.930 1015.060 ;
        RECT 2421.965 1014.750 2423.930 1015.050 ;
        RECT 2421.965 1014.735 2422.295 1014.750 ;
        RECT 2423.550 1014.740 2423.930 1014.750 ;
        RECT 1711.470 1008.620 1711.850 1008.940 ;
        RECT 1711.510 1007.580 1711.810 1008.620 ;
        RECT 2242.105 1007.580 2242.435 1007.585 ;
        RECT 1711.350 1007.270 1711.810 1007.580 ;
        RECT 2241.890 1007.570 2242.435 1007.580 ;
        RECT 2241.650 1007.270 2242.435 1007.570 ;
        RECT 1711.350 1007.260 1711.730 1007.270 ;
        RECT 2241.890 1007.260 2242.435 1007.270 ;
        RECT 2242.105 1007.255 2242.435 1007.260 ;
        RECT 1489.085 558.770 1489.415 558.785 ;
        RECT 1489.085 558.470 1503.890 558.770 ;
        RECT 1489.085 558.455 1489.415 558.470 ;
        RECT 1503.590 557.970 1503.890 558.470 ;
        RECT 1500.000 557.670 1504.600 557.970 ;
        RECT 1503.590 556.745 1503.890 557.670 ;
        RECT 1503.590 556.430 1504.135 556.745 ;
        RECT 1503.805 556.415 1504.135 556.430 ;
      LAYER met3 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
      LAYER met3 ;
        RECT 1898.945 913.730 1899.275 913.745 ;
        RECT 1889.070 913.610 1899.275 913.730 ;
        RECT 1881.880 913.430 1899.275 913.610 ;
        RECT 1881.880 913.310 1889.370 913.430 ;
        RECT 1898.945 913.415 1899.275 913.430 ;
        RECT 1881.880 904.890 1889.370 905.110 ;
        RECT 1902.165 904.890 1902.495 904.905 ;
        RECT 1881.880 904.810 1902.495 904.890 ;
        RECT 1889.070 904.590 1902.495 904.810 ;
        RECT 1902.165 904.575 1902.495 904.590 ;
        RECT 1898.945 628.130 1899.275 628.145 ;
        RECT 1899.865 628.130 1900.195 628.145 ;
        RECT 1898.945 627.830 1900.195 628.130 ;
        RECT 1898.945 627.815 1899.275 627.830 ;
        RECT 1899.865 627.815 1900.195 627.830 ;
        RECT 1904.005 615.890 1904.335 615.905 ;
        RECT 1889.070 615.870 1904.335 615.890 ;
        RECT 1881.880 615.590 1904.335 615.870 ;
        RECT 1881.880 615.570 1889.370 615.590 ;
        RECT 1904.005 615.575 1904.335 615.590 ;
        RECT 1901.705 610.450 1902.035 610.465 ;
        RECT 1885.390 610.150 1902.035 610.450 ;
        RECT 1885.390 607.370 1885.690 610.150 ;
        RECT 1901.705 610.135 1902.035 610.150 ;
        RECT 1881.880 607.070 1886.480 607.370 ;
        RECT 1881.880 601.610 1889.370 601.730 ;
        RECT 1901.245 601.610 1901.575 601.625 ;
        RECT 1881.880 601.430 1901.575 601.610 ;
        RECT 1889.070 601.310 1901.575 601.430 ;
        RECT 1901.245 601.295 1901.575 601.310 ;
        RECT 1899.865 596.170 1900.195 596.185 ;
        RECT 1885.390 595.870 1900.195 596.170 ;
        RECT 1885.390 593.230 1885.690 595.870 ;
        RECT 1899.865 595.855 1900.195 595.870 ;
        RECT 1881.880 592.930 1886.480 593.230 ;
        RECT 1904.005 590.730 1904.335 590.745 ;
        RECT 1885.390 590.430 1904.335 590.730 ;
        RECT 1885.390 587.590 1885.690 590.430 ;
        RECT 1904.005 590.415 1904.335 590.430 ;
        RECT 1881.880 587.290 1886.480 587.590 ;
        RECT 1904.005 579.170 1904.335 579.185 ;
        RECT 1889.070 579.090 1904.335 579.170 ;
        RECT 1881.880 578.870 1904.335 579.090 ;
        RECT 1881.880 578.790 1889.370 578.870 ;
        RECT 1904.005 578.855 1904.335 578.870 ;
        RECT 1903.545 573.730 1903.875 573.745 ;
        RECT 1889.070 573.450 1903.875 573.730 ;
        RECT 1881.880 573.430 1903.875 573.450 ;
        RECT 1881.880 573.150 1889.370 573.430 ;
        RECT 1903.545 573.415 1903.875 573.430 ;
        RECT 2100.000 557.670 2104.600 557.970 ;
        RECT 2083.865 556.730 2084.195 556.745 ;
        RECT 2100.670 556.730 2100.970 557.670 ;
        RECT 2083.865 556.430 2100.970 556.730 ;
        RECT 2083.865 556.415 2084.195 556.430 ;
      LAYER met3 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met3 ;
        RECT 2501.545 915.770 2501.875 915.785 ;
        RECT 2486.150 915.470 2501.875 915.770 ;
        RECT 2486.150 913.610 2486.450 915.470 ;
        RECT 2501.545 915.455 2501.875 915.470 ;
        RECT 2481.880 913.310 2486.480 913.610 ;
        RECT 2482.225 906.930 2482.555 906.945 ;
        RECT 2482.225 906.615 2482.770 906.930 ;
        RECT 2482.470 905.110 2482.770 906.615 ;
        RECT 2481.880 904.810 2486.480 905.110 ;
        RECT 2500.625 618.610 2500.955 618.625 ;
        RECT 2486.150 618.310 2500.955 618.610 ;
        RECT 2486.150 615.870 2486.450 618.310 ;
        RECT 2500.625 618.295 2500.955 618.310 ;
        RECT 2481.880 615.570 2486.480 615.870 ;
        RECT 2500.165 610.450 2500.495 610.465 ;
        RECT 2486.150 610.150 2500.495 610.450 ;
        RECT 2486.150 607.370 2486.450 610.150 ;
        RECT 2500.165 610.135 2500.495 610.150 ;
        RECT 2481.880 607.070 2486.480 607.370 ;
        RECT 2499.705 604.330 2500.035 604.345 ;
        RECT 2486.150 604.030 2500.035 604.330 ;
        RECT 2486.150 601.730 2486.450 604.030 ;
        RECT 2499.705 604.015 2500.035 604.030 ;
        RECT 2481.880 601.430 2486.480 601.730 ;
        RECT 2499.245 593.450 2499.575 593.465 ;
        RECT 2486.150 593.230 2499.575 593.450 ;
        RECT 2481.880 593.150 2499.575 593.230 ;
        RECT 2481.880 592.930 2486.480 593.150 ;
        RECT 2499.245 593.135 2499.575 593.150 ;
        RECT 2498.785 590.730 2499.115 590.745 ;
        RECT 2486.150 590.430 2499.115 590.730 ;
        RECT 2486.150 587.590 2486.450 590.430 ;
        RECT 2498.785 590.415 2499.115 590.430 ;
        RECT 2481.880 587.290 2486.480 587.590 ;
        RECT 2498.325 579.170 2498.655 579.185 ;
        RECT 2486.150 579.090 2498.655 579.170 ;
        RECT 2481.880 578.870 2498.655 579.090 ;
        RECT 2481.880 578.790 2486.480 578.870 ;
        RECT 2498.325 578.855 2498.655 578.870 ;
        RECT 2501.085 576.450 2501.415 576.465 ;
        RECT 2486.150 576.150 2501.415 576.450 ;
        RECT 2486.150 573.450 2486.450 576.150 ;
        RECT 2501.085 576.135 2501.415 576.150 ;
        RECT 2481.880 573.150 2486.480 573.450 ;
        RECT 1525.460 554.095 1527.200 555.000 ;
        RECT 2125.460 554.095 2127.200 555.000 ;
      LAYER via3 ;
        RECT 1867.900 3063.580 1868.220 3063.900 ;
        RECT 2442.900 3063.580 2443.220 3063.900 ;
        RECT 2469.580 3063.580 2469.900 3063.900 ;
        RECT 1845.820 3054.740 1846.140 3055.060 ;
        RECT 1865.140 3054.740 1865.460 3055.060 ;
        RECT 2139.840 2598.460 2140.160 2598.780 ;
        RECT 2169.040 2598.460 2169.360 2598.780 ;
        RECT 1568.900 2593.700 1569.220 2594.020 ;
        RECT 1598.340 2593.700 1598.660 2594.020 ;
        RECT 1617.660 2593.700 1617.980 2594.020 ;
        RECT 1621.340 2593.700 1621.660 2594.020 ;
        RECT 1625.940 2593.700 1626.260 2594.020 ;
        RECT 1632.380 2593.700 1632.700 2594.020 ;
        RECT 1636.980 2593.700 1637.300 2594.020 ;
        RECT 1644.340 2593.700 1644.660 2594.020 ;
        RECT 1650.780 2593.700 1651.100 2594.020 ;
        RECT 1658.140 2593.700 1658.460 2594.020 ;
        RECT 1661.820 2593.700 1662.140 2594.020 ;
        RECT 1668.260 2593.700 1668.580 2594.020 ;
        RECT 1672.860 2593.700 1673.180 2594.020 ;
        RECT 1679.300 2593.700 1679.620 2594.020 ;
        RECT 1684.820 2593.700 1685.140 2594.020 ;
        RECT 1690.340 2593.700 1690.660 2594.020 ;
        RECT 1697.700 2593.700 1698.020 2594.020 ;
        RECT 1702.300 2593.700 1702.620 2594.020 ;
        RECT 1707.820 2593.700 1708.140 2594.020 ;
        RECT 1725.300 2593.700 1725.620 2594.020 ;
        RECT 1732.660 2593.700 1732.980 2594.020 ;
        RECT 1744.620 2593.700 1744.940 2594.020 ;
        RECT 2215.660 2593.700 2215.980 2594.020 ;
        RECT 2256.140 2593.700 2256.460 2594.020 ;
        RECT 2262.580 2593.700 2262.900 2594.020 ;
        RECT 2292.020 2593.700 2292.340 2594.020 ;
        RECT 2302.140 2593.700 2302.460 2594.020 ;
        RECT 2332.500 2593.700 2332.820 2594.020 ;
        RECT 1562.460 2593.020 1562.780 2593.340 ;
        RECT 1580.860 2593.020 1581.180 2593.340 ;
        RECT 1592.820 2593.020 1593.140 2593.340 ;
        RECT 1603.860 2593.020 1604.180 2593.340 ;
        RECT 1615.820 2593.020 1616.140 2593.340 ;
        RECT 1656.300 2593.020 1656.620 2593.340 ;
        RECT 1703.220 2593.020 1703.540 2593.340 ;
        RECT 1738.180 2593.020 1738.500 2593.340 ;
        RECT 2148.500 2593.020 2148.820 2593.340 ;
        RECT 2208.300 2593.020 2208.620 2593.340 ;
        RECT 2220.260 2593.020 2220.580 2593.340 ;
        RECT 2226.700 2593.020 2227.020 2593.340 ;
        RECT 2233.140 2593.020 2233.460 2593.340 ;
        RECT 2285.580 2593.020 2285.900 2593.340 ;
        RECT 2305.820 2593.020 2306.140 2593.340 ;
        RECT 1575.340 2592.340 1575.660 2592.660 ;
        RECT 1582.700 2592.340 1583.020 2592.660 ;
        RECT 1586.380 2592.340 1586.700 2592.660 ;
        RECT 1592.820 2592.340 1593.140 2592.660 ;
        RECT 1608.460 2592.340 1608.780 2592.660 ;
        RECT 1651.700 2592.340 1652.020 2592.660 ;
        RECT 1715.180 2592.340 1715.500 2592.660 ;
        RECT 1744.620 2592.340 1744.940 2592.660 ;
        RECT 2132.860 2592.340 2133.180 2592.660 ;
        RECT 2219.340 2592.340 2219.660 2592.660 ;
        RECT 2224.860 2592.340 2225.180 2592.660 ;
        RECT 2238.660 2592.340 2238.980 2592.660 ;
        RECT 2244.180 2592.340 2244.500 2592.660 ;
        RECT 2268.100 2592.340 2268.420 2592.660 ;
        RECT 2273.620 2592.340 2273.940 2592.660 ;
        RECT 2280.060 2592.340 2280.380 2592.660 ;
        RECT 2312.260 2592.340 2312.580 2592.660 ;
        RECT 2319.620 2592.340 2319.940 2592.660 ;
        RECT 2337.100 2592.340 2337.420 2592.660 ;
        RECT 1569.820 2591.660 1570.140 2591.980 ;
        RECT 1604.780 2591.660 1605.100 2591.980 ;
        RECT 1686.660 2591.660 1686.980 2591.980 ;
        RECT 1692.180 2591.660 1692.500 2591.980 ;
        RECT 1699.540 2591.660 1699.860 2591.980 ;
        RECT 1718.860 2591.660 1719.180 2591.980 ;
        RECT 2154.020 2591.660 2154.340 2591.980 ;
        RECT 2175.180 2591.660 2175.500 2591.980 ;
        RECT 2227.620 2591.660 2227.940 2591.980 ;
        RECT 2234.980 2591.660 2235.300 2591.980 ;
        RECT 2250.620 2591.660 2250.940 2591.980 ;
        RECT 2297.540 2591.660 2297.860 2591.980 ;
        RECT 2326.060 2591.660 2326.380 2591.980 ;
        RECT 1610.300 2590.980 1610.620 2591.300 ;
        RECT 1669.180 2590.980 1669.500 2591.300 ;
        RECT 1709.660 2590.980 1709.980 2591.300 ;
        RECT 2145.740 2590.980 2146.060 2591.300 ;
        RECT 2180.700 2590.980 2181.020 2591.300 ;
        RECT 2203.700 2590.980 2204.020 2591.300 ;
        RECT 2241.420 2590.980 2241.740 2591.300 ;
        RECT 2342.620 2590.980 2342.940 2591.300 ;
        RECT 1573.500 2590.300 1573.820 2590.620 ;
        RECT 1600.180 2590.300 1600.500 2590.620 ;
        RECT 1587.300 2589.620 1587.620 2589.940 ;
        RECT 1563.380 2588.940 1563.700 2589.260 ;
        RECT 1674.700 2588.940 1675.020 2589.260 ;
        RECT 1717.020 2588.940 1717.340 2589.260 ;
        RECT 1739.100 2588.940 1739.420 2589.260 ;
        RECT 2163.220 2588.940 2163.540 2589.260 ;
        RECT 2186.220 2588.940 2186.540 2589.260 ;
        RECT 1548.660 2588.260 1548.980 2588.580 ;
        RECT 1622.260 2588.260 1622.580 2588.580 ;
        RECT 1633.300 2588.260 1633.620 2588.580 ;
        RECT 1639.740 2588.260 1640.060 2588.580 ;
        RECT 1645.260 2588.260 1645.580 2588.580 ;
        RECT 1662.740 2588.260 1663.060 2588.580 ;
        RECT 1680.220 2588.260 1680.540 2588.580 ;
        RECT 1721.620 2588.260 1721.940 2588.580 ;
        RECT 1727.140 2588.260 1727.460 2588.580 ;
        RECT 1733.580 2588.260 1733.900 2588.580 ;
        RECT 2165.060 2588.260 2165.380 2588.580 ;
        RECT 2169.660 2588.260 2169.980 2588.580 ;
        RECT 2178.860 2588.260 2179.180 2588.580 ;
        RECT 2184.380 2588.260 2184.700 2588.580 ;
        RECT 2189.900 2588.260 2190.220 2588.580 ;
        RECT 2266.260 2588.260 2266.580 2588.580 ;
        RECT 2301.220 2588.260 2301.540 2588.580 ;
        RECT 2341.700 2588.260 2342.020 2588.580 ;
        RECT 1536.700 2587.580 1537.020 2587.900 ;
        RECT 1543.140 2587.580 1543.460 2587.900 ;
        RECT 1551.420 2587.580 1551.740 2587.900 ;
        RECT 1558.780 2587.580 1559.100 2587.900 ;
        RECT 1627.780 2587.580 1628.100 2587.900 ;
        RECT 2191.740 2587.580 2192.060 2587.900 ;
        RECT 2193.580 2587.580 2193.900 2587.900 ;
        RECT 2198.180 2587.580 2198.500 2587.900 ;
        RECT 2200.020 2587.580 2200.340 2587.900 ;
        RECT 2207.380 2587.580 2207.700 2587.900 ;
        RECT 2213.820 2587.580 2214.140 2587.900 ;
        RECT 2248.780 2587.580 2249.100 2587.900 ;
        RECT 2254.300 2587.580 2254.620 2587.900 ;
        RECT 2259.820 2587.580 2260.140 2587.900 ;
        RECT 2269.020 2587.580 2269.340 2587.900 ;
        RECT 2276.380 2587.580 2276.700 2587.900 ;
        RECT 2281.900 2587.580 2282.220 2587.900 ;
        RECT 2289.260 2587.580 2289.580 2587.900 ;
        RECT 2295.700 2587.580 2296.020 2587.900 ;
        RECT 2303.980 2587.580 2304.300 2587.900 ;
        RECT 2310.420 2587.580 2310.740 2587.900 ;
        RECT 2317.780 2587.580 2318.100 2587.900 ;
        RECT 2324.220 2587.580 2324.540 2587.900 ;
        RECT 2330.660 2587.580 2330.980 2587.900 ;
        RECT 2336.180 2587.580 2336.500 2587.900 ;
        RECT 2345.380 2587.580 2345.700 2587.900 ;
        RECT 2169.660 2477.420 2169.980 2477.740 ;
        RECT 2169.660 2463.140 2169.980 2463.460 ;
        RECT 2370.220 1038.540 2370.540 1038.860 ;
        RECT 1796.140 1020.860 1796.460 1021.180 ;
        RECT 1830.180 1020.860 1830.500 1021.180 ;
        RECT 1855.020 1020.860 1855.340 1021.180 ;
        RECT 2282.820 1020.860 2283.140 1021.180 ;
        RECT 2340.780 1020.860 2341.100 1021.180 ;
        RECT 2351.820 1020.860 2352.140 1021.180 ;
        RECT 2387.700 1020.860 2388.020 1021.180 ;
        RECT 2395.980 1020.860 2396.300 1021.180 ;
        RECT 2408.860 1020.860 2409.180 1021.180 ;
        RECT 2451.180 1020.860 2451.500 1021.180 ;
        RECT 1801.660 1020.180 1801.980 1020.500 ;
        RECT 1837.540 1020.180 1837.860 1020.500 ;
        RECT 2246.940 1020.180 2247.260 1020.500 ;
        RECT 2335.260 1020.180 2335.580 1020.500 ;
        RECT 2346.300 1020.180 2346.620 1020.500 ;
        RECT 2381.260 1020.180 2381.580 1020.500 ;
        RECT 2390.460 1020.180 2390.780 1020.500 ;
        RECT 2429.100 1020.180 2429.420 1020.500 ;
        RECT 1808.100 1019.500 1808.420 1019.820 ;
        RECT 1832.020 1019.500 1832.340 1019.820 ;
        RECT 2402.420 1019.500 2402.740 1019.820 ;
        RECT 1814.540 1018.820 1814.860 1019.140 ;
        RECT 1821.900 1018.820 1822.220 1019.140 ;
        RECT 2241.420 1018.820 2241.740 1019.140 ;
        RECT 1640.660 1018.140 1640.980 1018.460 ;
        RECT 1647.100 1018.140 1647.420 1018.460 ;
        RECT 1653.540 1018.140 1653.860 1018.460 ;
        RECT 1674.700 1018.140 1675.020 1018.460 ;
        RECT 1714.260 1018.140 1714.580 1018.460 ;
        RECT 1719.780 1018.140 1720.100 1018.460 ;
        RECT 1745.540 1018.140 1745.860 1018.460 ;
        RECT 1755.660 1018.140 1755.980 1018.460 ;
        RECT 1700.460 1017.460 1700.780 1017.780 ;
        RECT 1704.140 1017.460 1704.460 1017.780 ;
        RECT 2415.300 1018.140 2415.620 1018.460 ;
        RECT 2437.380 1018.140 2437.700 1018.460 ;
        RECT 1641.580 1016.780 1641.900 1017.100 ;
        RECT 1661.820 1016.780 1662.140 1017.100 ;
        RECT 1664.580 1016.780 1664.900 1017.100 ;
        RECT 1682.980 1016.780 1683.300 1017.100 ;
        RECT 1691.260 1016.780 1691.580 1017.100 ;
        RECT 1786.940 1016.780 1787.260 1017.100 ;
        RECT 2247.860 1016.780 2248.180 1017.100 ;
        RECT 2254.300 1016.780 2254.620 1017.100 ;
        RECT 2260.740 1016.780 2261.060 1017.100 ;
        RECT 2266.260 1016.780 2266.580 1017.100 ;
        RECT 2280.060 1016.780 2280.380 1017.100 ;
        RECT 2293.860 1016.780 2294.180 1017.100 ;
        RECT 2304.900 1016.780 2305.220 1017.100 ;
        RECT 2311.340 1016.780 2311.660 1017.100 ;
        RECT 2393.220 1016.780 2393.540 1017.100 ;
        RECT 1655.380 1016.100 1655.700 1016.420 ;
        RECT 1658.140 1016.100 1658.460 1016.420 ;
        RECT 1670.100 1016.100 1670.420 1016.420 ;
        RECT 1681.140 1016.100 1681.460 1016.420 ;
        RECT 1684.820 1016.100 1685.140 1016.420 ;
        RECT 1697.700 1016.100 1698.020 1016.420 ;
        RECT 1726.220 1016.100 1726.540 1016.420 ;
        RECT 1749.220 1016.100 1749.540 1016.420 ;
        RECT 1843.060 1016.100 1843.380 1016.420 ;
        RECT 2253.380 1016.100 2253.700 1016.420 ;
        RECT 2264.420 1016.100 2264.740 1016.420 ;
        RECT 2274.540 1016.100 2274.860 1016.420 ;
        RECT 2276.380 1016.100 2276.700 1016.420 ;
        RECT 2287.420 1016.100 2287.740 1016.420 ;
        RECT 2300.300 1016.100 2300.620 1016.420 ;
        RECT 2315.940 1016.100 2316.260 1016.420 ;
        RECT 2323.300 1016.100 2323.620 1016.420 ;
        RECT 2329.740 1016.100 2330.060 1016.420 ;
        RECT 2358.260 1016.100 2358.580 1016.420 ;
        RECT 2363.780 1016.100 2364.100 1016.420 ;
        RECT 2375.740 1016.100 2376.060 1016.420 ;
        RECT 2388.620 1016.100 2388.940 1016.420 ;
        RECT 2421.740 1017.460 2422.060 1017.780 ;
        RECT 2442.900 1017.460 2443.220 1017.780 ;
        RECT 2431.860 1016.100 2432.180 1016.420 ;
        RECT 1648.020 1015.420 1648.340 1015.740 ;
        RECT 1668.260 1015.420 1668.580 1015.740 ;
        RECT 1673.780 1015.420 1674.100 1015.740 ;
        RECT 1708.740 1015.420 1709.060 1015.740 ;
        RECT 1732.660 1015.420 1732.980 1015.740 ;
        RECT 1739.100 1015.420 1739.420 1015.740 ;
        RECT 1763.940 1015.420 1764.260 1015.740 ;
        RECT 1765.780 1015.420 1766.100 1015.740 ;
        RECT 1774.060 1015.420 1774.380 1015.740 ;
        RECT 1780.500 1015.420 1780.820 1015.740 ;
        RECT 1788.780 1015.420 1789.100 1015.740 ;
        RECT 1680.220 1014.740 1680.540 1015.060 ;
        RECT 1689.420 1014.740 1689.740 1015.060 ;
        RECT 1695.860 1014.740 1696.180 1015.060 ;
        RECT 1711.500 1014.740 1711.820 1015.060 ;
        RECT 1712.420 1014.740 1712.740 1015.060 ;
        RECT 1717.940 1014.740 1718.260 1015.060 ;
        RECT 1724.380 1014.740 1724.700 1015.060 ;
        RECT 1729.900 1014.740 1730.220 1015.060 ;
        RECT 1735.420 1014.740 1735.740 1015.060 ;
        RECT 1741.860 1014.740 1742.180 1015.060 ;
        RECT 1748.300 1014.740 1748.620 1015.060 ;
        RECT 1754.740 1014.740 1755.060 1015.060 ;
        RECT 1758.420 1014.740 1758.740 1015.060 ;
        RECT 1766.700 1014.740 1767.020 1015.060 ;
        RECT 1771.300 1014.740 1771.620 1015.060 ;
        RECT 1777.740 1014.740 1778.060 1015.060 ;
        RECT 1782.340 1014.740 1782.660 1015.060 ;
        RECT 1789.700 1014.740 1790.020 1015.060 ;
        RECT 1793.380 1014.740 1793.700 1015.060 ;
        RECT 1799.820 1014.740 1800.140 1015.060 ;
        RECT 1806.260 1014.740 1806.580 1015.060 ;
        RECT 1812.700 1014.740 1813.020 1015.060 ;
        RECT 1817.300 1014.740 1817.620 1015.060 ;
        RECT 1823.740 1014.740 1824.060 1015.060 ;
        RECT 2258.900 1014.740 2259.220 1015.060 ;
        RECT 2270.860 1014.740 2271.180 1015.060 ;
        RECT 2281.900 1014.740 2282.220 1015.060 ;
        RECT 2289.260 1014.740 2289.580 1015.060 ;
        RECT 2294.780 1014.740 2295.100 1015.060 ;
        RECT 2302.140 1014.740 2302.460 1015.060 ;
        RECT 2307.660 1014.740 2307.980 1015.060 ;
        RECT 2312.260 1014.740 2312.580 1015.060 ;
        RECT 2317.780 1014.740 2318.100 1015.060 ;
        RECT 2322.380 1014.740 2322.700 1015.060 ;
        RECT 2328.820 1014.740 2329.140 1015.060 ;
        RECT 2336.180 1014.740 2336.500 1015.060 ;
        RECT 2342.620 1014.740 2342.940 1015.060 ;
        RECT 2347.220 1014.740 2347.540 1015.060 ;
        RECT 2353.660 1014.740 2353.980 1015.060 ;
        RECT 2359.180 1014.740 2359.500 1015.060 ;
        RECT 2364.700 1014.740 2365.020 1015.060 ;
        RECT 2371.140 1014.740 2371.460 1015.060 ;
        RECT 2377.580 1014.740 2377.900 1015.060 ;
        RECT 2382.180 1014.740 2382.500 1015.060 ;
        RECT 2399.660 1014.740 2399.980 1015.060 ;
        RECT 2406.100 1014.740 2406.420 1015.060 ;
        RECT 2410.700 1014.740 2411.020 1015.060 ;
        RECT 2417.140 1014.740 2417.460 1015.060 ;
        RECT 2423.580 1014.740 2423.900 1015.060 ;
        RECT 1711.500 1008.620 1711.820 1008.940 ;
        RECT 1711.380 1007.260 1711.700 1007.580 ;
        RECT 2241.920 1007.260 2242.240 1007.580 ;
      LAYER met4 ;
        RECT 1867.895 3063.575 1868.225 3063.905 ;
        RECT 2442.895 3063.575 2443.225 3063.905 ;
        RECT 2469.575 3063.575 2469.905 3063.905 ;
        RECT 1867.910 3056.235 1868.210 3063.575 ;
        RECT 2442.910 3056.235 2443.210 3063.575 ;
        RECT 1594.025 3051.635 1594.325 3056.235 ;
        RECT 1600.265 3051.635 1600.565 3056.235 ;
        RECT 1606.505 3051.635 1606.805 3056.235 ;
        RECT 1612.745 3051.635 1613.045 3056.235 ;
        RECT 1618.985 3051.635 1619.285 3056.235 ;
        RECT 1625.225 3051.635 1625.525 3056.235 ;
        RECT 1631.465 3051.635 1631.765 3056.235 ;
        RECT 1637.705 3051.635 1638.005 3056.235 ;
        RECT 1643.945 3051.635 1644.245 3056.235 ;
        RECT 1650.185 3051.635 1650.485 3056.235 ;
        RECT 1656.425 3051.635 1656.725 3056.235 ;
        RECT 1662.665 3051.635 1662.965 3056.235 ;
        RECT 1668.905 3051.635 1669.205 3056.235 ;
        RECT 1675.145 3051.635 1675.445 3056.235 ;
        RECT 1681.385 3051.635 1681.685 3056.235 ;
        RECT 1687.625 3051.635 1687.925 3056.235 ;
        RECT 1693.865 3051.635 1694.165 3056.235 ;
        RECT 1700.105 3051.635 1700.405 3056.235 ;
        RECT 1706.345 3051.635 1706.645 3056.235 ;
        RECT 1712.585 3051.635 1712.885 3056.235 ;
        RECT 1718.825 3051.635 1719.125 3056.235 ;
        RECT 1725.065 3051.635 1725.365 3056.235 ;
        RECT 1731.305 3051.635 1731.605 3056.235 ;
        RECT 1737.545 3051.635 1737.845 3056.235 ;
        RECT 1743.785 3051.635 1744.085 3056.235 ;
        RECT 1750.025 3051.635 1750.325 3056.235 ;
        RECT 1756.265 3051.635 1756.565 3056.235 ;
        RECT 1762.505 3051.635 1762.805 3056.235 ;
        RECT 1768.745 3051.635 1769.045 3056.235 ;
        RECT 1774.985 3051.635 1775.285 3056.235 ;
        RECT 1781.225 3051.635 1781.525 3056.235 ;
        RECT 1787.465 3051.635 1787.765 3056.235 ;
        RECT 1842.890 3055.050 1843.190 3056.235 ;
        RECT 1845.815 3055.050 1846.145 3055.065 ;
        RECT 1842.890 3054.750 1846.145 3055.050 ;
        RECT 1842.890 3051.635 1843.190 3054.750 ;
        RECT 1845.815 3054.735 1846.145 3054.750 ;
        RECT 1865.135 3055.050 1865.465 3055.065 ;
        RECT 1867.865 3055.050 1868.210 3056.235 ;
        RECT 1865.135 3054.750 1868.210 3055.050 ;
        RECT 1865.135 3054.735 1865.465 3054.750 ;
        RECT 1867.865 3051.635 1868.165 3054.750 ;
        RECT 2194.025 3051.635 2194.325 3056.235 ;
        RECT 2200.265 3051.635 2200.565 3056.235 ;
        RECT 2206.505 3051.635 2206.805 3056.235 ;
        RECT 2212.745 3051.635 2213.045 3056.235 ;
        RECT 2218.985 3051.635 2219.285 3056.235 ;
        RECT 2225.225 3051.635 2225.525 3056.235 ;
        RECT 2231.465 3051.635 2231.765 3056.235 ;
        RECT 2237.705 3051.635 2238.005 3056.235 ;
        RECT 2243.945 3051.635 2244.245 3056.235 ;
        RECT 2250.185 3051.635 2250.485 3056.235 ;
        RECT 2256.425 3051.635 2256.725 3056.235 ;
        RECT 2262.665 3051.635 2262.965 3056.235 ;
        RECT 2268.905 3051.635 2269.205 3056.235 ;
        RECT 2275.145 3051.635 2275.445 3056.235 ;
        RECT 2281.385 3051.635 2281.685 3056.235 ;
        RECT 2287.625 3051.635 2287.925 3056.235 ;
        RECT 2293.865 3051.635 2294.165 3056.235 ;
        RECT 2300.105 3051.635 2300.405 3056.235 ;
        RECT 2306.345 3051.635 2306.645 3056.235 ;
        RECT 2312.585 3051.635 2312.885 3056.235 ;
        RECT 2318.825 3051.635 2319.125 3056.235 ;
        RECT 2325.065 3051.635 2325.365 3056.235 ;
        RECT 2331.305 3051.635 2331.605 3056.235 ;
        RECT 2337.545 3051.635 2337.845 3056.235 ;
        RECT 2343.785 3051.635 2344.085 3056.235 ;
        RECT 2350.025 3051.635 2350.325 3056.235 ;
        RECT 2356.265 3051.635 2356.565 3056.235 ;
        RECT 2362.505 3051.635 2362.805 3056.235 ;
        RECT 2368.745 3051.635 2369.045 3056.235 ;
        RECT 2374.985 3051.635 2375.285 3056.235 ;
        RECT 2381.225 3051.635 2381.525 3056.235 ;
        RECT 2387.465 3051.635 2387.765 3056.235 ;
        RECT 2442.890 3054.750 2443.210 3056.235 ;
        RECT 2467.865 3055.050 2468.165 3056.235 ;
        RECT 2469.590 3055.050 2469.890 3063.575 ;
        RECT 2467.865 3054.750 2469.890 3055.050 ;
        RECT 2442.890 3051.635 2443.190 3054.750 ;
        RECT 2467.865 3051.635 2468.165 3054.750 ;
      LAYER met4 ;
        RECT 1505.000 2605.000 1881.480 3051.235 ;
        RECT 2105.000 2605.000 2481.480 3051.235 ;
      LAYER met4 ;
        RECT 1534.010 2601.150 1534.310 2604.600 ;
        RECT 1539.850 2601.150 1540.150 2604.600 ;
        RECT 1545.690 2601.150 1545.990 2604.600 ;
        RECT 1551.530 2601.150 1551.830 2604.600 ;
        RECT 1534.010 2600.850 1537.010 2601.150 ;
        RECT 1534.010 2600.000 1534.310 2600.850 ;
        RECT 1536.710 2587.905 1537.010 2600.850 ;
        RECT 1539.850 2600.850 1543.450 2601.150 ;
        RECT 1539.850 2600.000 1540.150 2600.850 ;
        RECT 1543.150 2587.905 1543.450 2600.850 ;
        RECT 1545.690 2600.850 1548.970 2601.150 ;
        RECT 1545.690 2600.000 1545.990 2600.850 ;
        RECT 1548.670 2588.585 1548.970 2600.850 ;
        RECT 1551.430 2600.000 1551.830 2601.150 ;
        RECT 1557.370 2601.150 1557.670 2604.600 ;
        RECT 1563.210 2601.150 1563.510 2604.600 ;
        RECT 1557.370 2600.850 1559.090 2601.150 ;
        RECT 1557.370 2600.000 1557.670 2600.850 ;
        RECT 1548.655 2588.255 1548.985 2588.585 ;
        RECT 1551.430 2587.905 1551.730 2600.000 ;
        RECT 1558.790 2587.905 1559.090 2600.850 ;
        RECT 1562.470 2600.850 1563.510 2601.150 ;
        RECT 1562.470 2593.345 1562.770 2600.850 ;
        RECT 1563.210 2600.000 1563.510 2600.850 ;
        RECT 1563.830 2599.450 1564.130 2604.600 ;
        RECT 1569.050 2601.150 1569.350 2604.600 ;
        RECT 1563.390 2599.150 1564.130 2599.450 ;
        RECT 1568.910 2600.000 1569.350 2601.150 ;
        RECT 1569.670 2601.150 1569.970 2604.600 ;
        RECT 1574.890 2602.850 1575.190 2604.600 ;
        RECT 1573.510 2602.550 1575.190 2602.850 ;
        RECT 1569.670 2600.000 1570.130 2601.150 ;
        RECT 1562.455 2593.015 1562.785 2593.345 ;
        RECT 1563.390 2589.265 1563.690 2599.150 ;
        RECT 1568.910 2594.025 1569.210 2600.000 ;
        RECT 1568.895 2593.695 1569.225 2594.025 ;
        RECT 1569.830 2591.985 1570.130 2600.000 ;
        RECT 1569.815 2591.655 1570.145 2591.985 ;
        RECT 1573.510 2590.625 1573.810 2602.550 ;
        RECT 1574.890 2600.000 1575.190 2602.550 ;
        RECT 1575.510 2599.450 1575.810 2604.600 ;
        RECT 1575.350 2599.150 1575.810 2599.450 ;
        RECT 1580.730 2599.450 1581.030 2604.600 ;
        RECT 1581.350 2602.850 1581.650 2604.600 ;
        RECT 1581.350 2602.550 1583.010 2602.850 ;
        RECT 1581.350 2600.000 1581.650 2602.550 ;
        RECT 1580.730 2599.150 1581.170 2599.450 ;
        RECT 1575.350 2592.665 1575.650 2599.150 ;
        RECT 1580.870 2593.345 1581.170 2599.150 ;
        RECT 1580.855 2593.015 1581.185 2593.345 ;
        RECT 1582.710 2592.665 1583.010 2602.550 ;
        RECT 1586.570 2601.150 1586.870 2604.600 ;
        RECT 1586.390 2600.000 1586.870 2601.150 ;
        RECT 1587.190 2601.150 1587.490 2604.600 ;
        RECT 1587.190 2600.000 1587.610 2601.150 ;
        RECT 1586.390 2592.665 1586.690 2600.000 ;
        RECT 1575.335 2592.335 1575.665 2592.665 ;
        RECT 1582.695 2592.335 1583.025 2592.665 ;
        RECT 1586.375 2592.335 1586.705 2592.665 ;
        RECT 1573.495 2590.295 1573.825 2590.625 ;
        RECT 1587.310 2589.945 1587.610 2600.000 ;
        RECT 1592.410 2599.450 1592.710 2604.600 ;
        RECT 1593.030 2601.150 1593.330 2604.600 ;
        RECT 1593.030 2600.850 1594.050 2601.150 ;
        RECT 1593.030 2600.000 1593.330 2600.850 ;
        RECT 1592.410 2599.150 1593.130 2599.450 ;
        RECT 1592.830 2593.345 1593.130 2599.150 ;
        RECT 1592.815 2593.015 1593.145 2593.345 ;
        RECT 1592.815 2592.650 1593.145 2592.665 ;
        RECT 1593.750 2592.650 1594.050 2600.850 ;
        RECT 1598.250 2599.450 1598.550 2604.600 ;
        RECT 1598.870 2602.850 1599.170 2604.600 ;
        RECT 1598.870 2602.550 1600.490 2602.850 ;
        RECT 1598.870 2600.000 1599.170 2602.550 ;
        RECT 1598.250 2599.150 1598.650 2599.450 ;
        RECT 1598.350 2594.025 1598.650 2599.150 ;
        RECT 1598.335 2593.695 1598.665 2594.025 ;
        RECT 1592.815 2592.350 1594.050 2592.650 ;
        RECT 1592.815 2592.335 1593.145 2592.350 ;
        RECT 1600.190 2590.625 1600.490 2602.550 ;
        RECT 1604.090 2601.150 1604.390 2604.600 ;
        RECT 1603.870 2600.000 1604.390 2601.150 ;
        RECT 1604.710 2601.150 1605.010 2604.600 ;
        RECT 1609.930 2602.850 1610.230 2604.600 ;
        RECT 1608.470 2602.550 1610.230 2602.850 ;
        RECT 1604.710 2600.000 1605.090 2601.150 ;
        RECT 1603.870 2593.345 1604.170 2600.000 ;
        RECT 1603.855 2593.015 1604.185 2593.345 ;
        RECT 1604.790 2591.985 1605.090 2600.000 ;
        RECT 1608.470 2592.665 1608.770 2602.550 ;
        RECT 1609.930 2600.000 1610.230 2602.550 ;
        RECT 1610.550 2599.450 1610.850 2604.600 ;
        RECT 1610.310 2599.150 1610.850 2599.450 ;
        RECT 1615.770 2599.450 1616.070 2604.600 ;
        RECT 1616.390 2602.850 1616.690 2604.600 ;
        RECT 1616.390 2602.550 1617.970 2602.850 ;
        RECT 1616.390 2600.000 1616.690 2602.550 ;
        RECT 1615.770 2599.150 1616.130 2599.450 ;
        RECT 1608.455 2592.335 1608.785 2592.665 ;
        RECT 1604.775 2591.655 1605.105 2591.985 ;
        RECT 1610.310 2591.305 1610.610 2599.150 ;
        RECT 1615.830 2593.345 1616.130 2599.150 ;
        RECT 1617.670 2594.025 1617.970 2602.550 ;
        RECT 1621.610 2601.150 1621.910 2604.600 ;
        RECT 1621.350 2600.000 1621.910 2601.150 ;
        RECT 1622.230 2601.150 1622.530 2604.600 ;
        RECT 1627.450 2602.850 1627.750 2604.600 ;
        RECT 1625.950 2602.550 1627.750 2602.850 ;
        RECT 1622.230 2600.000 1622.570 2601.150 ;
        RECT 1621.350 2594.025 1621.650 2600.000 ;
        RECT 1617.655 2593.695 1617.985 2594.025 ;
        RECT 1621.335 2593.695 1621.665 2594.025 ;
        RECT 1615.815 2593.015 1616.145 2593.345 ;
        RECT 1610.295 2590.975 1610.625 2591.305 ;
        RECT 1600.175 2590.295 1600.505 2590.625 ;
        RECT 1587.295 2589.615 1587.625 2589.945 ;
        RECT 1563.375 2588.935 1563.705 2589.265 ;
        RECT 1622.270 2588.585 1622.570 2600.000 ;
        RECT 1625.950 2594.025 1626.250 2602.550 ;
        RECT 1627.450 2600.000 1627.750 2602.550 ;
        RECT 1628.070 2599.450 1628.370 2604.600 ;
        RECT 1633.290 2601.150 1633.590 2604.600 ;
        RECT 1627.790 2599.150 1628.370 2599.450 ;
        RECT 1632.390 2600.850 1633.590 2601.150 ;
        RECT 1625.935 2593.695 1626.265 2594.025 ;
        RECT 1622.255 2588.255 1622.585 2588.585 ;
        RECT 1627.790 2587.905 1628.090 2599.150 ;
        RECT 1632.390 2594.025 1632.690 2600.850 ;
        RECT 1633.290 2600.000 1633.590 2600.850 ;
        RECT 1633.910 2599.450 1634.210 2604.600 ;
        RECT 1639.130 2601.150 1639.430 2604.600 ;
        RECT 1633.310 2599.150 1634.210 2599.450 ;
        RECT 1636.990 2600.850 1639.430 2601.150 ;
        RECT 1632.375 2593.695 1632.705 2594.025 ;
        RECT 1633.310 2588.585 1633.610 2599.150 ;
        RECT 1636.990 2594.025 1637.290 2600.850 ;
        RECT 1639.130 2600.000 1639.430 2600.850 ;
        RECT 1636.975 2593.695 1637.305 2594.025 ;
        RECT 1639.750 2588.585 1640.050 2604.600 ;
        RECT 1644.970 2601.150 1645.270 2604.600 ;
        RECT 1644.350 2600.850 1645.270 2601.150 ;
        RECT 1644.350 2594.025 1644.650 2600.850 ;
        RECT 1644.970 2600.000 1645.270 2600.850 ;
        RECT 1645.590 2599.450 1645.890 2604.600 ;
        RECT 1650.810 2601.150 1651.110 2604.600 ;
        RECT 1645.270 2599.150 1645.890 2599.450 ;
        RECT 1650.790 2600.000 1651.110 2601.150 ;
        RECT 1651.430 2601.150 1651.730 2604.600 ;
        RECT 1651.430 2600.000 1652.010 2601.150 ;
        RECT 1644.335 2593.695 1644.665 2594.025 ;
        RECT 1645.270 2588.585 1645.570 2599.150 ;
        RECT 1650.790 2594.025 1651.090 2600.000 ;
        RECT 1650.775 2593.695 1651.105 2594.025 ;
        RECT 1651.710 2592.665 1652.010 2600.000 ;
        RECT 1656.650 2599.450 1656.950 2604.600 ;
        RECT 1657.270 2601.150 1657.570 2604.600 ;
        RECT 1662.490 2601.150 1662.790 2604.600 ;
        RECT 1657.270 2600.850 1658.450 2601.150 ;
        RECT 1657.270 2600.000 1657.570 2600.850 ;
        RECT 1656.310 2599.150 1656.950 2599.450 ;
        RECT 1656.310 2593.345 1656.610 2599.150 ;
        RECT 1658.150 2594.025 1658.450 2600.850 ;
        RECT 1661.830 2600.850 1662.790 2601.150 ;
        RECT 1661.830 2594.025 1662.130 2600.850 ;
        RECT 1662.490 2600.000 1662.790 2600.850 ;
        RECT 1663.110 2599.450 1663.410 2604.600 ;
        RECT 1668.330 2601.150 1668.630 2604.600 ;
        RECT 1662.750 2599.150 1663.410 2599.450 ;
        RECT 1668.270 2600.000 1668.630 2601.150 ;
        RECT 1668.950 2601.150 1669.250 2604.600 ;
        RECT 1674.170 2602.850 1674.470 2604.600 ;
        RECT 1672.870 2602.550 1674.470 2602.850 ;
        RECT 1668.950 2600.000 1669.490 2601.150 ;
        RECT 1658.135 2593.695 1658.465 2594.025 ;
        RECT 1661.815 2593.695 1662.145 2594.025 ;
        RECT 1656.295 2593.015 1656.625 2593.345 ;
        RECT 1651.695 2592.335 1652.025 2592.665 ;
        RECT 1662.750 2588.585 1663.050 2599.150 ;
        RECT 1668.270 2594.025 1668.570 2600.000 ;
        RECT 1668.255 2593.695 1668.585 2594.025 ;
        RECT 1669.190 2591.305 1669.490 2600.000 ;
        RECT 1672.870 2594.025 1673.170 2602.550 ;
        RECT 1674.170 2600.000 1674.470 2602.550 ;
        RECT 1674.790 2599.450 1675.090 2604.600 ;
        RECT 1680.010 2601.150 1680.310 2604.600 ;
        RECT 1674.710 2599.150 1675.090 2599.450 ;
        RECT 1679.310 2600.850 1680.310 2601.150 ;
        RECT 1672.855 2593.695 1673.185 2594.025 ;
        RECT 1669.175 2590.975 1669.505 2591.305 ;
        RECT 1674.710 2589.265 1675.010 2599.150 ;
        RECT 1679.310 2594.025 1679.610 2600.850 ;
        RECT 1680.010 2600.000 1680.310 2600.850 ;
        RECT 1680.630 2599.450 1680.930 2604.600 ;
        RECT 1685.850 2601.150 1686.150 2604.600 ;
        RECT 1680.230 2599.150 1680.930 2599.450 ;
        RECT 1684.830 2600.850 1686.150 2601.150 ;
        RECT 1679.295 2593.695 1679.625 2594.025 ;
        RECT 1674.695 2588.935 1675.025 2589.265 ;
        RECT 1680.230 2588.585 1680.530 2599.150 ;
        RECT 1684.830 2594.025 1685.130 2600.850 ;
        RECT 1685.850 2600.000 1686.150 2600.850 ;
        RECT 1686.470 2601.150 1686.770 2604.600 ;
        RECT 1691.690 2602.850 1691.990 2604.600 ;
        RECT 1690.350 2602.550 1691.990 2602.850 ;
        RECT 1686.470 2600.000 1686.970 2601.150 ;
        RECT 1684.815 2593.695 1685.145 2594.025 ;
        RECT 1686.670 2591.985 1686.970 2600.000 ;
        RECT 1690.350 2594.025 1690.650 2602.550 ;
        RECT 1691.690 2600.000 1691.990 2602.550 ;
        RECT 1692.310 2599.450 1692.610 2604.600 ;
        RECT 1692.190 2599.150 1692.610 2599.450 ;
        RECT 1697.530 2599.450 1697.830 2604.600 ;
        RECT 1698.150 2602.850 1698.450 2604.600 ;
        RECT 1698.150 2602.550 1699.850 2602.850 ;
        RECT 1698.150 2600.000 1698.450 2602.550 ;
        RECT 1697.530 2599.150 1698.010 2599.450 ;
        RECT 1690.335 2593.695 1690.665 2594.025 ;
        RECT 1692.190 2591.985 1692.490 2599.150 ;
        RECT 1697.710 2594.025 1698.010 2599.150 ;
        RECT 1697.695 2593.695 1698.025 2594.025 ;
        RECT 1699.550 2591.985 1699.850 2602.550 ;
        RECT 1703.370 2601.150 1703.670 2604.600 ;
        RECT 1702.310 2600.850 1703.670 2601.150 ;
        RECT 1702.310 2594.025 1702.610 2600.850 ;
        RECT 1703.370 2600.000 1703.670 2600.850 ;
        RECT 1703.990 2599.450 1704.290 2604.600 ;
        RECT 1709.210 2602.850 1709.510 2604.600 ;
        RECT 1703.230 2599.150 1704.290 2599.450 ;
        RECT 1707.830 2602.550 1709.510 2602.850 ;
        RECT 1702.295 2593.695 1702.625 2594.025 ;
        RECT 1703.230 2593.345 1703.530 2599.150 ;
        RECT 1707.830 2594.025 1708.130 2602.550 ;
        RECT 1709.210 2600.000 1709.510 2602.550 ;
        RECT 1709.830 2599.450 1710.130 2604.600 ;
        RECT 1709.670 2599.150 1710.130 2599.450 ;
        RECT 1715.050 2599.450 1715.350 2604.600 ;
        RECT 1715.670 2602.850 1715.970 2604.600 ;
        RECT 1715.670 2602.550 1717.330 2602.850 ;
        RECT 1715.670 2600.000 1715.970 2602.550 ;
        RECT 1715.050 2599.150 1715.490 2599.450 ;
        RECT 1707.815 2593.695 1708.145 2594.025 ;
        RECT 1703.215 2593.015 1703.545 2593.345 ;
        RECT 1686.655 2591.655 1686.985 2591.985 ;
        RECT 1692.175 2591.655 1692.505 2591.985 ;
        RECT 1699.535 2591.655 1699.865 2591.985 ;
        RECT 1709.670 2591.305 1709.970 2599.150 ;
        RECT 1715.190 2592.665 1715.490 2599.150 ;
        RECT 1715.175 2592.335 1715.505 2592.665 ;
        RECT 1709.655 2590.975 1709.985 2591.305 ;
        RECT 1717.030 2589.265 1717.330 2602.550 ;
        RECT 1720.890 2601.150 1721.190 2604.600 ;
        RECT 1718.870 2600.850 1721.190 2601.150 ;
        RECT 1718.870 2591.985 1719.170 2600.850 ;
        RECT 1720.890 2600.000 1721.190 2600.850 ;
        RECT 1721.510 2601.150 1721.810 2604.600 ;
        RECT 1726.730 2601.150 1727.030 2604.600 ;
        RECT 1721.510 2600.000 1721.930 2601.150 ;
        RECT 1718.855 2591.655 1719.185 2591.985 ;
        RECT 1717.015 2588.935 1717.345 2589.265 ;
        RECT 1721.630 2588.585 1721.930 2600.000 ;
        RECT 1725.310 2600.850 1727.030 2601.150 ;
        RECT 1725.310 2594.025 1725.610 2600.850 ;
        RECT 1726.730 2600.000 1727.030 2600.850 ;
        RECT 1727.350 2599.450 1727.650 2604.600 ;
        RECT 1727.150 2599.150 1727.650 2599.450 ;
        RECT 1725.295 2593.695 1725.625 2594.025 ;
        RECT 1727.150 2588.585 1727.450 2599.150 ;
        RECT 1732.570 2596.050 1732.870 2604.600 ;
        RECT 1733.190 2599.450 1733.490 2604.600 ;
        RECT 1738.410 2601.150 1738.710 2604.600 ;
        RECT 1738.190 2600.000 1738.710 2601.150 ;
        RECT 1739.030 2601.150 1739.330 2604.600 ;
        RECT 1739.030 2600.000 1739.410 2601.150 ;
        RECT 1733.190 2599.150 1733.890 2599.450 ;
        RECT 1732.570 2595.750 1732.970 2596.050 ;
        RECT 1732.670 2594.025 1732.970 2595.750 ;
        RECT 1732.655 2593.695 1732.985 2594.025 ;
        RECT 1733.590 2588.585 1733.890 2599.150 ;
        RECT 1738.190 2593.345 1738.490 2600.000 ;
        RECT 1738.175 2593.015 1738.505 2593.345 ;
        RECT 1739.110 2589.265 1739.410 2600.000 ;
        RECT 1744.250 2599.450 1744.550 2604.600 ;
        RECT 1744.870 2601.150 1745.170 2604.600 ;
        RECT 2134.010 2601.150 2134.310 2604.600 ;
        RECT 1744.870 2600.850 1745.850 2601.150 ;
        RECT 1744.870 2600.000 1745.170 2600.850 ;
        RECT 1744.250 2599.150 1744.930 2599.450 ;
        RECT 1744.630 2594.025 1744.930 2599.150 ;
        RECT 1744.615 2593.695 1744.945 2594.025 ;
        RECT 1744.615 2592.650 1744.945 2592.665 ;
        RECT 1745.550 2592.650 1745.850 2600.850 ;
        RECT 2132.870 2600.850 2134.310 2601.150 ;
        RECT 2132.870 2592.665 2133.170 2600.850 ;
        RECT 2134.010 2600.000 2134.310 2600.850 ;
        RECT 2139.850 2598.785 2140.150 2604.600 ;
        RECT 2145.690 2601.150 2145.990 2604.600 ;
        RECT 2151.530 2601.150 2151.830 2604.600 ;
        RECT 2157.370 2601.150 2157.670 2604.600 ;
        RECT 2145.690 2600.000 2146.050 2601.150 ;
        RECT 2139.835 2598.455 2140.165 2598.785 ;
        RECT 1744.615 2592.350 1745.850 2592.650 ;
        RECT 1744.615 2592.335 1744.945 2592.350 ;
        RECT 2132.855 2592.335 2133.185 2592.665 ;
        RECT 2145.750 2591.305 2146.050 2600.000 ;
        RECT 2148.510 2600.850 2151.830 2601.150 ;
        RECT 2148.510 2593.345 2148.810 2600.850 ;
        RECT 2151.530 2600.000 2151.830 2600.850 ;
        RECT 2154.030 2600.850 2157.670 2601.150 ;
        RECT 2148.495 2593.015 2148.825 2593.345 ;
        RECT 2154.030 2591.985 2154.330 2600.850 ;
        RECT 2157.370 2600.000 2157.670 2600.850 ;
        RECT 2163.210 2599.450 2163.510 2604.600 ;
        RECT 2163.830 2601.150 2164.130 2604.600 ;
        RECT 2163.830 2600.850 2165.370 2601.150 ;
        RECT 2163.830 2600.000 2164.130 2600.850 ;
        RECT 2163.210 2599.150 2163.530 2599.450 ;
        RECT 2154.015 2591.655 2154.345 2591.985 ;
        RECT 2145.735 2590.975 2146.065 2591.305 ;
        RECT 2163.230 2589.265 2163.530 2599.150 ;
        RECT 1739.095 2588.935 1739.425 2589.265 ;
        RECT 2163.215 2588.935 2163.545 2589.265 ;
        RECT 2165.070 2588.585 2165.370 2600.850 ;
        RECT 2169.050 2598.785 2169.350 2604.600 ;
        RECT 2169.035 2598.455 2169.365 2598.785 ;
        RECT 2169.670 2588.585 2169.970 2604.600 ;
        RECT 2174.890 2599.450 2175.190 2604.600 ;
        RECT 2175.510 2601.150 2175.810 2604.600 ;
        RECT 2180.730 2601.150 2181.030 2604.600 ;
        RECT 2175.510 2600.850 2179.170 2601.150 ;
        RECT 2175.510 2600.000 2175.810 2600.850 ;
        RECT 2174.890 2599.150 2175.490 2599.450 ;
        RECT 2175.190 2591.985 2175.490 2599.150 ;
        RECT 2175.175 2591.655 2175.505 2591.985 ;
        RECT 2178.870 2588.585 2179.170 2600.850 ;
        RECT 2180.710 2600.000 2181.030 2601.150 ;
        RECT 2181.350 2601.150 2181.650 2604.600 ;
        RECT 2181.350 2600.850 2184.690 2601.150 ;
        RECT 2181.350 2600.000 2181.650 2600.850 ;
        RECT 2180.710 2591.305 2181.010 2600.000 ;
        RECT 2180.695 2590.975 2181.025 2591.305 ;
        RECT 2184.390 2588.585 2184.690 2600.850 ;
        RECT 2186.570 2599.450 2186.870 2604.600 ;
        RECT 2187.190 2601.150 2187.490 2604.600 ;
        RECT 2192.410 2601.150 2192.710 2604.600 ;
        RECT 2187.190 2600.850 2190.210 2601.150 ;
        RECT 2187.190 2600.000 2187.490 2600.850 ;
        RECT 2186.230 2599.150 2186.870 2599.450 ;
        RECT 2186.230 2589.265 2186.530 2599.150 ;
        RECT 2186.215 2588.935 2186.545 2589.265 ;
        RECT 2189.910 2588.585 2190.210 2600.850 ;
        RECT 2191.750 2600.850 2192.710 2601.150 ;
        RECT 1633.295 2588.255 1633.625 2588.585 ;
        RECT 1639.735 2588.255 1640.065 2588.585 ;
        RECT 1645.255 2588.255 1645.585 2588.585 ;
        RECT 1662.735 2588.255 1663.065 2588.585 ;
        RECT 1680.215 2588.255 1680.545 2588.585 ;
        RECT 1721.615 2588.255 1721.945 2588.585 ;
        RECT 1727.135 2588.255 1727.465 2588.585 ;
        RECT 1733.575 2588.255 1733.905 2588.585 ;
        RECT 2165.055 2588.255 2165.385 2588.585 ;
        RECT 2169.655 2588.255 2169.985 2588.585 ;
        RECT 2178.855 2588.255 2179.185 2588.585 ;
        RECT 2184.375 2588.255 2184.705 2588.585 ;
        RECT 2189.895 2588.255 2190.225 2588.585 ;
        RECT 2191.750 2587.905 2192.050 2600.850 ;
        RECT 2192.410 2600.000 2192.710 2600.850 ;
        RECT 2193.030 2599.450 2193.330 2604.600 ;
        RECT 2198.250 2601.150 2198.550 2604.600 ;
        RECT 2198.190 2600.000 2198.550 2601.150 ;
        RECT 2198.870 2601.150 2199.170 2604.600 ;
        RECT 2198.870 2600.850 2200.330 2601.150 ;
        RECT 2198.870 2600.000 2199.170 2600.850 ;
        RECT 2193.030 2599.150 2193.890 2599.450 ;
        RECT 2193.590 2587.905 2193.890 2599.150 ;
        RECT 2198.190 2587.905 2198.490 2600.000 ;
        RECT 2200.030 2587.905 2200.330 2600.850 ;
        RECT 2204.090 2599.450 2204.390 2604.600 ;
        RECT 2204.710 2601.150 2205.010 2604.600 ;
        RECT 2209.930 2601.150 2210.230 2604.600 ;
        RECT 2204.710 2600.850 2207.690 2601.150 ;
        RECT 2204.710 2600.000 2205.010 2600.850 ;
        RECT 2203.710 2599.150 2204.390 2599.450 ;
        RECT 2203.710 2591.305 2204.010 2599.150 ;
        RECT 2203.695 2590.975 2204.025 2591.305 ;
        RECT 2207.390 2587.905 2207.690 2600.850 ;
        RECT 2208.310 2600.850 2210.230 2601.150 ;
        RECT 2208.310 2593.345 2208.610 2600.850 ;
        RECT 2209.930 2600.000 2210.230 2600.850 ;
        RECT 2210.550 2601.150 2210.850 2604.600 ;
        RECT 2215.770 2601.150 2216.070 2604.600 ;
        RECT 2210.550 2600.850 2214.130 2601.150 ;
        RECT 2210.550 2600.000 2210.850 2600.850 ;
        RECT 2208.295 2593.015 2208.625 2593.345 ;
        RECT 2213.830 2587.905 2214.130 2600.850 ;
        RECT 2215.670 2600.000 2216.070 2601.150 ;
        RECT 2216.390 2601.150 2216.690 2604.600 ;
        RECT 2221.610 2601.150 2221.910 2604.600 ;
        RECT 2216.390 2600.850 2219.650 2601.150 ;
        RECT 2216.390 2600.000 2216.690 2600.850 ;
        RECT 2215.670 2594.025 2215.970 2600.000 ;
        RECT 2215.655 2593.695 2215.985 2594.025 ;
        RECT 2219.350 2592.665 2219.650 2600.850 ;
        RECT 2220.270 2600.850 2221.910 2601.150 ;
        RECT 2220.270 2593.345 2220.570 2600.850 ;
        RECT 2221.610 2600.000 2221.910 2600.850 ;
        RECT 2222.230 2601.150 2222.530 2604.600 ;
        RECT 2227.450 2601.150 2227.750 2604.600 ;
        RECT 2222.230 2600.850 2225.170 2601.150 ;
        RECT 2222.230 2600.000 2222.530 2600.850 ;
        RECT 2220.255 2593.015 2220.585 2593.345 ;
        RECT 2224.870 2592.665 2225.170 2600.850 ;
        RECT 2226.710 2600.850 2227.750 2601.150 ;
        RECT 2226.710 2593.345 2227.010 2600.850 ;
        RECT 2227.450 2600.000 2227.750 2600.850 ;
        RECT 2228.070 2599.450 2228.370 2604.600 ;
        RECT 2233.290 2601.150 2233.590 2604.600 ;
        RECT 2227.630 2599.150 2228.370 2599.450 ;
        RECT 2233.150 2600.000 2233.590 2601.150 ;
        RECT 2233.910 2601.150 2234.210 2604.600 ;
        RECT 2233.910 2600.850 2235.290 2601.150 ;
        RECT 2233.910 2600.000 2234.210 2600.850 ;
        RECT 2226.695 2593.015 2227.025 2593.345 ;
        RECT 2219.335 2592.335 2219.665 2592.665 ;
        RECT 2224.855 2592.335 2225.185 2592.665 ;
        RECT 2227.630 2591.985 2227.930 2599.150 ;
        RECT 2233.150 2593.345 2233.450 2600.000 ;
        RECT 2233.135 2593.015 2233.465 2593.345 ;
        RECT 2234.990 2591.985 2235.290 2600.850 ;
        RECT 2239.130 2599.450 2239.430 2604.600 ;
        RECT 2239.750 2601.150 2240.050 2604.600 ;
        RECT 2244.970 2601.150 2245.270 2604.600 ;
        RECT 2239.750 2600.850 2241.730 2601.150 ;
        RECT 2239.750 2600.000 2240.050 2600.850 ;
        RECT 2238.670 2599.150 2239.430 2599.450 ;
        RECT 2238.670 2592.665 2238.970 2599.150 ;
        RECT 2238.655 2592.335 2238.985 2592.665 ;
        RECT 2227.615 2591.655 2227.945 2591.985 ;
        RECT 2234.975 2591.655 2235.305 2591.985 ;
        RECT 2241.430 2591.305 2241.730 2600.850 ;
        RECT 2244.190 2600.850 2245.270 2601.150 ;
        RECT 2244.190 2592.665 2244.490 2600.850 ;
        RECT 2244.970 2600.000 2245.270 2600.850 ;
        RECT 2245.590 2601.150 2245.890 2604.600 ;
        RECT 2250.810 2601.150 2251.110 2604.600 ;
        RECT 2245.590 2600.850 2249.090 2601.150 ;
        RECT 2245.590 2600.000 2245.890 2600.850 ;
        RECT 2244.175 2592.335 2244.505 2592.665 ;
        RECT 2241.415 2590.975 2241.745 2591.305 ;
        RECT 2248.790 2587.905 2249.090 2600.850 ;
        RECT 2250.630 2600.000 2251.110 2601.150 ;
        RECT 2251.430 2601.150 2251.730 2604.600 ;
        RECT 2251.430 2600.850 2254.610 2601.150 ;
        RECT 2251.430 2600.000 2251.730 2600.850 ;
        RECT 2250.630 2591.985 2250.930 2600.000 ;
        RECT 2250.615 2591.655 2250.945 2591.985 ;
        RECT 2254.310 2587.905 2254.610 2600.850 ;
        RECT 2256.650 2599.450 2256.950 2604.600 ;
        RECT 2257.270 2601.150 2257.570 2604.600 ;
        RECT 2257.270 2600.850 2260.130 2601.150 ;
        RECT 2257.270 2600.000 2257.570 2600.850 ;
        RECT 2256.150 2599.150 2256.950 2599.450 ;
        RECT 2256.150 2594.025 2256.450 2599.150 ;
        RECT 2256.135 2593.695 2256.465 2594.025 ;
        RECT 2259.830 2587.905 2260.130 2600.850 ;
        RECT 2262.490 2599.450 2262.790 2604.600 ;
        RECT 2263.110 2601.150 2263.410 2604.600 ;
        RECT 2268.330 2601.150 2268.630 2604.600 ;
        RECT 2263.110 2600.850 2266.570 2601.150 ;
        RECT 2263.110 2600.000 2263.410 2600.850 ;
        RECT 2262.490 2599.150 2262.890 2599.450 ;
        RECT 2262.590 2594.025 2262.890 2599.150 ;
        RECT 2262.575 2593.695 2262.905 2594.025 ;
        RECT 2266.270 2588.585 2266.570 2600.850 ;
        RECT 2268.110 2600.000 2268.630 2601.150 ;
        RECT 2268.950 2601.150 2269.250 2604.600 ;
        RECT 2268.950 2600.000 2269.330 2601.150 ;
        RECT 2268.110 2592.665 2268.410 2600.000 ;
        RECT 2268.095 2592.335 2268.425 2592.665 ;
        RECT 2266.255 2588.255 2266.585 2588.585 ;
        RECT 2269.030 2587.905 2269.330 2600.000 ;
        RECT 2274.170 2599.450 2274.470 2604.600 ;
        RECT 2274.790 2601.150 2275.090 2604.600 ;
        RECT 2274.790 2600.850 2276.690 2601.150 ;
        RECT 2274.790 2600.000 2275.090 2600.850 ;
        RECT 2273.630 2599.150 2274.470 2599.450 ;
        RECT 2273.630 2592.665 2273.930 2599.150 ;
        RECT 2273.615 2592.335 2273.945 2592.665 ;
        RECT 2276.390 2587.905 2276.690 2600.850 ;
        RECT 2280.010 2599.450 2280.310 2604.600 ;
        RECT 2280.630 2601.150 2280.930 2604.600 ;
        RECT 2285.850 2601.150 2286.150 2604.600 ;
        RECT 2280.630 2600.850 2282.210 2601.150 ;
        RECT 2280.630 2600.000 2280.930 2600.850 ;
        RECT 2280.010 2599.150 2280.370 2599.450 ;
        RECT 2280.070 2592.665 2280.370 2599.150 ;
        RECT 2280.055 2592.335 2280.385 2592.665 ;
        RECT 2281.910 2587.905 2282.210 2600.850 ;
        RECT 2285.590 2600.000 2286.150 2601.150 ;
        RECT 2286.470 2601.150 2286.770 2604.600 ;
        RECT 2286.470 2600.850 2289.570 2601.150 ;
        RECT 2286.470 2600.000 2286.770 2600.850 ;
        RECT 2285.590 2593.345 2285.890 2600.000 ;
        RECT 2285.575 2593.015 2285.905 2593.345 ;
        RECT 2289.270 2587.905 2289.570 2600.850 ;
        RECT 2291.690 2599.450 2291.990 2604.600 ;
        RECT 2292.310 2601.150 2292.610 2604.600 ;
        RECT 2292.310 2600.850 2296.010 2601.150 ;
        RECT 2292.310 2600.000 2292.610 2600.850 ;
        RECT 2291.690 2599.150 2292.330 2599.450 ;
        RECT 2292.030 2594.025 2292.330 2599.150 ;
        RECT 2292.015 2593.695 2292.345 2594.025 ;
        RECT 2295.710 2587.905 2296.010 2600.850 ;
        RECT 2297.530 2599.450 2297.830 2604.600 ;
        RECT 2298.150 2601.150 2298.450 2604.600 ;
        RECT 2303.370 2601.150 2303.670 2604.600 ;
        RECT 2298.150 2600.850 2301.530 2601.150 ;
        RECT 2298.150 2600.000 2298.450 2600.850 ;
        RECT 2297.530 2599.150 2297.850 2599.450 ;
        RECT 2297.550 2591.985 2297.850 2599.150 ;
        RECT 2297.535 2591.655 2297.865 2591.985 ;
        RECT 2301.230 2588.585 2301.530 2600.850 ;
        RECT 2302.150 2600.850 2303.670 2601.150 ;
        RECT 2302.150 2594.025 2302.450 2600.850 ;
        RECT 2303.370 2600.000 2303.670 2600.850 ;
        RECT 2302.135 2593.695 2302.465 2594.025 ;
        RECT 2301.215 2588.255 2301.545 2588.585 ;
        RECT 2303.990 2587.905 2304.290 2604.600 ;
        RECT 2309.210 2601.150 2309.510 2604.600 ;
        RECT 2305.830 2600.850 2309.510 2601.150 ;
        RECT 2305.830 2593.345 2306.130 2600.850 ;
        RECT 2309.210 2600.000 2309.510 2600.850 ;
        RECT 2309.830 2601.150 2310.130 2604.600 ;
        RECT 2315.050 2601.150 2315.350 2604.600 ;
        RECT 2309.830 2600.850 2310.730 2601.150 ;
        RECT 2309.830 2600.000 2310.130 2600.850 ;
        RECT 2305.815 2593.015 2306.145 2593.345 ;
        RECT 2310.430 2587.905 2310.730 2600.850 ;
        RECT 2312.270 2600.850 2315.350 2601.150 ;
        RECT 2312.270 2592.665 2312.570 2600.850 ;
        RECT 2315.050 2600.000 2315.350 2600.850 ;
        RECT 2315.670 2601.150 2315.970 2604.600 ;
        RECT 2320.890 2601.150 2321.190 2604.600 ;
        RECT 2315.670 2600.850 2318.090 2601.150 ;
        RECT 2315.670 2600.000 2315.970 2600.850 ;
        RECT 2312.255 2592.335 2312.585 2592.665 ;
        RECT 2317.790 2587.905 2318.090 2600.850 ;
        RECT 2319.630 2600.850 2321.190 2601.150 ;
        RECT 2319.630 2592.665 2319.930 2600.850 ;
        RECT 2320.890 2600.000 2321.190 2600.850 ;
        RECT 2321.510 2601.150 2321.810 2604.600 ;
        RECT 2326.730 2601.150 2327.030 2604.600 ;
        RECT 2321.510 2600.850 2324.530 2601.150 ;
        RECT 2321.510 2600.000 2321.810 2600.850 ;
        RECT 2319.615 2592.335 2319.945 2592.665 ;
        RECT 2324.230 2587.905 2324.530 2600.850 ;
        RECT 2326.070 2600.850 2327.030 2601.150 ;
        RECT 2326.070 2591.985 2326.370 2600.850 ;
        RECT 2326.730 2600.000 2327.030 2600.850 ;
        RECT 2327.350 2601.150 2327.650 2604.600 ;
        RECT 2332.570 2601.150 2332.870 2604.600 ;
        RECT 2327.350 2600.850 2330.970 2601.150 ;
        RECT 2327.350 2600.000 2327.650 2600.850 ;
        RECT 2326.055 2591.655 2326.385 2591.985 ;
        RECT 2330.670 2587.905 2330.970 2600.850 ;
        RECT 2332.510 2600.000 2332.870 2601.150 ;
        RECT 2333.190 2601.150 2333.490 2604.600 ;
        RECT 2338.410 2601.150 2338.710 2604.600 ;
        RECT 2333.190 2600.850 2336.490 2601.150 ;
        RECT 2333.190 2600.000 2333.490 2600.850 ;
        RECT 2332.510 2594.025 2332.810 2600.000 ;
        RECT 2332.495 2593.695 2332.825 2594.025 ;
        RECT 2336.190 2587.905 2336.490 2600.850 ;
        RECT 2337.110 2600.850 2338.710 2601.150 ;
        RECT 2337.110 2592.665 2337.410 2600.850 ;
        RECT 2338.410 2600.000 2338.710 2600.850 ;
        RECT 2339.030 2601.150 2339.330 2604.600 ;
        RECT 2344.250 2601.150 2344.550 2604.600 ;
        RECT 2339.030 2600.850 2342.010 2601.150 ;
        RECT 2339.030 2600.000 2339.330 2600.850 ;
        RECT 2337.095 2592.335 2337.425 2592.665 ;
        RECT 2341.710 2588.585 2342.010 2600.850 ;
        RECT 2342.630 2600.850 2344.550 2601.150 ;
        RECT 2342.630 2591.305 2342.930 2600.850 ;
        RECT 2344.250 2600.000 2344.550 2600.850 ;
        RECT 2344.870 2599.450 2345.170 2604.600 ;
        RECT 2344.870 2599.150 2345.690 2599.450 ;
        RECT 2342.615 2590.975 2342.945 2591.305 ;
        RECT 2341.695 2588.255 2342.025 2588.585 ;
        RECT 2345.390 2587.905 2345.690 2599.150 ;
        RECT 1536.695 2587.575 1537.025 2587.905 ;
        RECT 1543.135 2587.575 1543.465 2587.905 ;
        RECT 1551.415 2587.575 1551.745 2587.905 ;
        RECT 1558.775 2587.575 1559.105 2587.905 ;
        RECT 1627.775 2587.575 1628.105 2587.905 ;
        RECT 2191.735 2587.575 2192.065 2587.905 ;
        RECT 2193.575 2587.575 2193.905 2587.905 ;
        RECT 2198.175 2587.575 2198.505 2587.905 ;
        RECT 2200.015 2587.575 2200.345 2587.905 ;
        RECT 2207.375 2587.575 2207.705 2587.905 ;
        RECT 2213.815 2587.575 2214.145 2587.905 ;
        RECT 2248.775 2587.575 2249.105 2587.905 ;
        RECT 2254.295 2587.575 2254.625 2587.905 ;
        RECT 2259.815 2587.575 2260.145 2587.905 ;
        RECT 2269.015 2587.575 2269.345 2587.905 ;
        RECT 2276.375 2587.575 2276.705 2587.905 ;
        RECT 2281.895 2587.575 2282.225 2587.905 ;
        RECT 2289.255 2587.575 2289.585 2587.905 ;
        RECT 2295.695 2587.575 2296.025 2587.905 ;
        RECT 2303.975 2587.575 2304.305 2587.905 ;
        RECT 2310.415 2587.575 2310.745 2587.905 ;
        RECT 2317.775 2587.575 2318.105 2587.905 ;
        RECT 2324.215 2587.575 2324.545 2587.905 ;
        RECT 2330.655 2587.575 2330.985 2587.905 ;
        RECT 2336.175 2587.575 2336.505 2587.905 ;
        RECT 2345.375 2587.575 2345.705 2587.905 ;
        RECT 1498.020 2415.000 1501.020 2585.000 ;
        RECT 1678.020 2415.000 1681.020 2585.000 ;
        RECT 1858.020 2415.000 1861.020 2585.000 ;
        RECT 2169.655 2477.415 2169.985 2477.745 ;
        RECT 2169.670 2463.465 2169.970 2477.415 ;
        RECT 2169.655 2463.135 2169.985 2463.465 ;
        RECT 2218.020 2415.000 2221.020 2585.000 ;
        RECT 2398.020 2415.000 2401.020 2585.000 ;
      LAYER met4 ;
        RECT 1316.855 1210.240 1320.640 2388.880 ;
        RECT 1323.040 1210.240 1397.440 2388.880 ;
        RECT 1399.840 1210.240 2678.785 2388.880 ;
        RECT 1316.855 1206.295 2678.785 1210.240 ;
      LAYER met4 ;
        RECT 1552.020 1021.235 1555.020 1185.000 ;
        RECT 1732.020 1021.235 1735.020 1185.000 ;
        RECT 2092.020 1021.235 2095.020 1185.000 ;
        RECT 2272.020 1021.235 2275.020 1185.000 ;
        RECT 2370.215 1038.535 2370.545 1038.865 ;
        RECT 1796.135 1020.855 1796.465 1021.185 ;
        RECT 1830.175 1020.855 1830.505 1021.185 ;
        RECT 1855.015 1020.855 1855.345 1021.185 ;
        RECT 2282.815 1020.855 2283.145 1021.185 ;
        RECT 2340.775 1020.855 2341.105 1021.185 ;
        RECT 2351.815 1020.855 2352.145 1021.185 ;
        RECT 1640.655 1018.135 1640.985 1018.465 ;
        RECT 1647.095 1018.135 1647.425 1018.465 ;
        RECT 1653.535 1018.135 1653.865 1018.465 ;
        RECT 1674.695 1018.135 1675.025 1018.465 ;
        RECT 1714.255 1018.135 1714.585 1018.465 ;
        RECT 1719.775 1018.135 1720.105 1018.465 ;
        RECT 1745.535 1018.135 1745.865 1018.465 ;
        RECT 1755.655 1018.135 1755.985 1018.465 ;
        RECT 1640.670 1004.850 1640.970 1018.135 ;
        RECT 1641.575 1016.775 1641.905 1017.105 ;
        RECT 1641.590 1008.250 1641.890 1016.775 ;
        RECT 1641.590 1007.950 1642.230 1008.250 ;
        RECT 1641.310 1004.850 1641.610 1006.235 ;
        RECT 1640.670 1004.550 1641.610 1004.850 ;
        RECT 1641.310 1001.635 1641.610 1004.550 ;
        RECT 1641.930 1001.635 1642.230 1007.950 ;
        RECT 1647.110 1006.235 1647.410 1018.135 ;
        RECT 1648.015 1015.415 1648.345 1015.745 ;
        RECT 1648.030 1006.235 1648.330 1015.415 ;
        RECT 1653.550 1008.250 1653.850 1018.135 ;
        RECT 1661.815 1016.775 1662.145 1017.105 ;
        RECT 1664.575 1016.775 1664.905 1017.105 ;
        RECT 1655.375 1016.095 1655.705 1016.425 ;
        RECT 1658.135 1016.095 1658.465 1016.425 ;
        RECT 1647.110 1004.550 1647.450 1006.235 ;
        RECT 1647.150 1001.635 1647.450 1004.550 ;
        RECT 1647.770 1004.550 1648.330 1006.235 ;
        RECT 1652.990 1007.950 1653.850 1008.250 ;
        RECT 1647.770 1001.635 1648.070 1004.550 ;
        RECT 1652.990 1001.635 1653.290 1007.950 ;
        RECT 1653.610 1004.850 1653.910 1006.235 ;
        RECT 1655.390 1004.850 1655.690 1016.095 ;
        RECT 1653.610 1004.550 1655.690 1004.850 ;
        RECT 1658.150 1004.850 1658.450 1016.095 ;
        RECT 1658.830 1004.850 1659.130 1006.235 ;
        RECT 1658.150 1004.550 1659.130 1004.850 ;
        RECT 1653.610 1001.635 1653.910 1004.550 ;
        RECT 1658.830 1001.635 1659.130 1004.550 ;
        RECT 1659.450 1004.850 1659.750 1006.235 ;
        RECT 1661.830 1004.850 1662.130 1016.775 ;
        RECT 1659.450 1004.550 1662.130 1004.850 ;
        RECT 1664.590 1006.235 1664.890 1016.775 ;
        RECT 1670.095 1016.095 1670.425 1016.425 ;
        RECT 1668.255 1015.415 1668.585 1015.745 ;
        RECT 1664.590 1004.550 1664.970 1006.235 ;
        RECT 1659.450 1001.635 1659.750 1004.550 ;
        RECT 1664.670 1001.635 1664.970 1004.550 ;
        RECT 1665.290 1004.850 1665.590 1006.235 ;
        RECT 1668.270 1004.850 1668.570 1015.415 ;
        RECT 1670.110 1008.250 1670.410 1016.095 ;
        RECT 1673.775 1015.415 1674.105 1015.745 ;
        RECT 1670.110 1007.950 1670.810 1008.250 ;
        RECT 1665.290 1004.550 1668.570 1004.850 ;
        RECT 1665.290 1001.635 1665.590 1004.550 ;
        RECT 1670.510 1001.635 1670.810 1007.950 ;
        RECT 1671.130 1004.850 1671.430 1006.235 ;
        RECT 1673.790 1004.850 1674.090 1015.415 ;
        RECT 1671.130 1004.550 1674.090 1004.850 ;
        RECT 1674.710 1004.850 1675.010 1018.135 ;
        RECT 1700.455 1017.455 1700.785 1017.785 ;
        RECT 1704.135 1017.455 1704.465 1017.785 ;
        RECT 1682.975 1016.775 1683.305 1017.105 ;
        RECT 1691.255 1016.775 1691.585 1017.105 ;
        RECT 1681.135 1016.095 1681.465 1016.425 ;
        RECT 1680.215 1014.735 1680.545 1015.065 ;
        RECT 1676.350 1004.850 1676.650 1006.235 ;
        RECT 1674.710 1004.550 1676.650 1004.850 ;
        RECT 1671.130 1001.635 1671.430 1004.550 ;
        RECT 1676.350 1001.635 1676.650 1004.550 ;
        RECT 1676.970 1004.850 1677.270 1006.235 ;
        RECT 1680.230 1004.850 1680.530 1014.735 ;
        RECT 1676.970 1004.550 1680.530 1004.850 ;
        RECT 1681.150 1004.850 1681.450 1016.095 ;
        RECT 1682.990 1006.235 1683.290 1016.775 ;
        RECT 1684.815 1016.095 1685.145 1016.425 ;
        RECT 1682.190 1004.850 1682.490 1006.235 ;
        RECT 1681.150 1004.550 1682.490 1004.850 ;
        RECT 1676.970 1001.635 1677.270 1004.550 ;
        RECT 1682.190 1001.635 1682.490 1004.550 ;
        RECT 1682.810 1004.550 1683.290 1006.235 ;
        RECT 1684.830 1004.850 1685.130 1016.095 ;
        RECT 1689.415 1014.735 1689.745 1015.065 ;
        RECT 1688.030 1004.850 1688.330 1006.235 ;
        RECT 1684.830 1004.550 1688.330 1004.850 ;
        RECT 1682.810 1001.635 1683.110 1004.550 ;
        RECT 1688.030 1001.635 1688.330 1004.550 ;
        RECT 1688.650 1004.850 1688.950 1006.235 ;
        RECT 1689.430 1004.850 1689.730 1014.735 ;
        RECT 1688.650 1004.550 1689.730 1004.850 ;
        RECT 1691.270 1004.850 1691.570 1016.775 ;
        RECT 1697.695 1016.095 1698.025 1016.425 ;
        RECT 1695.855 1014.735 1696.185 1015.065 ;
        RECT 1693.870 1004.850 1694.170 1006.235 ;
        RECT 1691.270 1004.550 1694.170 1004.850 ;
        RECT 1688.650 1001.635 1688.950 1004.550 ;
        RECT 1693.870 1001.635 1694.170 1004.550 ;
        RECT 1694.490 1004.085 1694.790 1006.235 ;
        RECT 1695.870 1004.085 1696.170 1014.735 ;
        RECT 1697.710 1004.850 1698.010 1016.095 ;
        RECT 1700.470 1006.235 1700.770 1017.455 ;
        RECT 1699.710 1004.850 1700.010 1006.235 ;
        RECT 1697.710 1004.550 1700.010 1004.850 ;
        RECT 1694.490 1003.785 1696.170 1004.085 ;
        RECT 1694.490 1001.635 1694.790 1003.785 ;
        RECT 1699.710 1001.635 1700.010 1004.550 ;
        RECT 1700.330 1004.550 1700.770 1006.235 ;
        RECT 1700.330 1001.635 1700.630 1004.550 ;
        RECT 1704.150 1004.085 1704.450 1017.455 ;
        RECT 1708.735 1015.415 1709.065 1015.745 ;
        RECT 1705.550 1004.085 1705.850 1006.235 ;
        RECT 1704.150 1003.785 1705.850 1004.085 ;
        RECT 1705.550 1001.635 1705.850 1003.785 ;
        RECT 1706.170 1004.850 1706.470 1006.235 ;
        RECT 1708.750 1004.850 1709.050 1015.415 ;
        RECT 1711.495 1014.735 1711.825 1015.065 ;
        RECT 1712.415 1014.735 1712.745 1015.065 ;
        RECT 1711.510 1008.945 1711.810 1014.735 ;
        RECT 1711.495 1008.615 1711.825 1008.945 ;
        RECT 1712.430 1008.250 1712.730 1014.735 ;
        RECT 1712.010 1007.950 1712.730 1008.250 ;
        RECT 1711.375 1007.255 1711.705 1007.585 ;
        RECT 1706.170 1004.550 1709.050 1004.850 ;
        RECT 1706.170 1001.635 1706.470 1004.550 ;
        RECT 1711.390 1001.635 1711.690 1007.255 ;
        RECT 1712.010 1001.635 1712.310 1007.950 ;
        RECT 1714.270 1004.850 1714.570 1018.135 ;
        RECT 1717.935 1014.735 1718.265 1015.065 ;
        RECT 1717.950 1006.235 1718.250 1014.735 ;
        RECT 1717.230 1004.850 1717.530 1006.235 ;
        RECT 1714.270 1004.550 1717.530 1004.850 ;
        RECT 1717.230 1001.635 1717.530 1004.550 ;
        RECT 1717.850 1004.550 1718.250 1006.235 ;
        RECT 1719.790 1004.850 1720.090 1018.135 ;
        RECT 1726.215 1016.095 1726.545 1016.425 ;
        RECT 1724.375 1014.735 1724.705 1015.065 ;
        RECT 1723.070 1004.850 1723.370 1006.235 ;
        RECT 1719.790 1004.550 1723.370 1004.850 ;
        RECT 1717.850 1001.635 1718.150 1004.550 ;
        RECT 1723.070 1001.635 1723.370 1004.550 ;
        RECT 1723.690 1004.850 1723.990 1006.235 ;
        RECT 1724.390 1004.850 1724.690 1014.735 ;
        RECT 1723.690 1004.550 1724.690 1004.850 ;
        RECT 1726.230 1004.850 1726.530 1016.095 ;
        RECT 1732.655 1015.415 1732.985 1015.745 ;
        RECT 1739.095 1015.415 1739.425 1015.745 ;
        RECT 1729.895 1014.735 1730.225 1015.065 ;
        RECT 1729.910 1008.250 1730.210 1014.735 ;
        RECT 1729.530 1007.950 1730.210 1008.250 ;
        RECT 1728.910 1004.850 1729.210 1006.235 ;
        RECT 1726.230 1004.550 1729.210 1004.850 ;
        RECT 1723.690 1001.635 1723.990 1004.550 ;
        RECT 1728.910 1001.635 1729.210 1004.550 ;
        RECT 1729.530 1001.635 1729.830 1007.950 ;
        RECT 1732.670 1004.850 1732.970 1015.415 ;
        RECT 1735.415 1014.735 1735.745 1015.065 ;
        RECT 1735.430 1006.235 1735.730 1014.735 ;
        RECT 1734.750 1004.850 1735.050 1006.235 ;
        RECT 1732.670 1004.550 1735.050 1004.850 ;
        RECT 1734.750 1001.635 1735.050 1004.550 ;
        RECT 1735.370 1004.550 1735.730 1006.235 ;
        RECT 1739.110 1004.850 1739.410 1015.415 ;
        RECT 1741.855 1014.735 1742.185 1015.065 ;
        RECT 1740.590 1004.850 1740.890 1006.235 ;
        RECT 1739.110 1004.550 1740.890 1004.850 ;
        RECT 1735.370 1001.635 1735.670 1004.550 ;
        RECT 1740.590 1001.635 1740.890 1004.550 ;
        RECT 1741.210 1004.850 1741.510 1006.235 ;
        RECT 1741.870 1004.850 1742.170 1014.735 ;
        RECT 1741.210 1004.550 1742.170 1004.850 ;
        RECT 1745.550 1004.850 1745.850 1018.135 ;
        RECT 1749.215 1016.095 1749.545 1016.425 ;
        RECT 1748.295 1014.735 1748.625 1015.065 ;
        RECT 1746.430 1004.850 1746.730 1006.235 ;
        RECT 1745.550 1004.550 1746.730 1004.850 ;
        RECT 1741.210 1001.635 1741.510 1004.550 ;
        RECT 1746.430 1001.635 1746.730 1004.550 ;
        RECT 1747.050 1004.085 1747.350 1006.235 ;
        RECT 1748.310 1004.085 1748.610 1014.735 ;
        RECT 1749.230 1004.850 1749.530 1016.095 ;
        RECT 1754.735 1014.735 1755.065 1015.065 ;
        RECT 1752.270 1004.850 1752.570 1006.235 ;
        RECT 1749.230 1004.550 1752.570 1004.850 ;
        RECT 1747.050 1003.785 1748.610 1004.085 ;
        RECT 1747.050 1001.635 1747.350 1003.785 ;
        RECT 1752.270 1001.635 1752.570 1004.550 ;
        RECT 1752.890 1004.850 1753.190 1006.235 ;
        RECT 1754.750 1004.850 1755.050 1014.735 ;
        RECT 1752.890 1004.550 1755.050 1004.850 ;
        RECT 1755.670 1004.850 1755.970 1018.135 ;
        RECT 1786.935 1016.775 1787.265 1017.105 ;
        RECT 1763.935 1015.415 1764.265 1015.745 ;
        RECT 1765.775 1015.415 1766.105 1015.745 ;
        RECT 1774.055 1015.415 1774.385 1015.745 ;
        RECT 1780.495 1015.415 1780.825 1015.745 ;
        RECT 1758.415 1014.735 1758.745 1015.065 ;
        RECT 1758.430 1008.250 1758.730 1014.735 ;
        RECT 1758.430 1007.950 1759.030 1008.250 ;
        RECT 1758.110 1004.850 1758.410 1006.235 ;
        RECT 1755.670 1004.550 1758.410 1004.850 ;
        RECT 1752.890 1001.635 1753.190 1004.550 ;
        RECT 1758.110 1001.635 1758.410 1004.550 ;
        RECT 1758.730 1001.635 1759.030 1007.950 ;
        RECT 1763.950 1001.635 1764.250 1015.415 ;
        RECT 1764.570 1004.850 1764.870 1006.235 ;
        RECT 1765.790 1004.850 1766.090 1015.415 ;
        RECT 1766.695 1014.735 1767.025 1015.065 ;
        RECT 1771.295 1014.735 1771.625 1015.065 ;
        RECT 1764.570 1004.550 1766.090 1004.850 ;
        RECT 1766.710 1004.850 1767.010 1014.735 ;
        RECT 1769.790 1004.850 1770.090 1006.235 ;
        RECT 1766.710 1004.550 1770.090 1004.850 ;
        RECT 1764.570 1001.635 1764.870 1004.550 ;
        RECT 1769.790 1001.635 1770.090 1004.550 ;
        RECT 1770.410 1004.850 1770.710 1006.235 ;
        RECT 1771.310 1004.850 1771.610 1014.735 ;
        RECT 1770.410 1004.550 1771.610 1004.850 ;
        RECT 1774.070 1004.850 1774.370 1015.415 ;
        RECT 1777.735 1014.735 1778.065 1015.065 ;
        RECT 1775.630 1004.850 1775.930 1006.235 ;
        RECT 1774.070 1004.550 1775.930 1004.850 ;
        RECT 1770.410 1001.635 1770.710 1004.550 ;
        RECT 1775.630 1001.635 1775.930 1004.550 ;
        RECT 1776.250 1004.085 1776.550 1006.235 ;
        RECT 1777.750 1004.085 1778.050 1014.735 ;
        RECT 1780.510 1004.850 1780.810 1015.415 ;
        RECT 1782.335 1014.735 1782.665 1015.065 ;
        RECT 1782.350 1006.235 1782.650 1014.735 ;
        RECT 1786.950 1008.250 1787.250 1016.775 ;
        RECT 1788.775 1015.415 1789.105 1015.745 ;
        RECT 1786.950 1007.950 1787.610 1008.250 ;
        RECT 1781.470 1004.850 1781.770 1006.235 ;
        RECT 1780.510 1004.550 1781.770 1004.850 ;
        RECT 1776.250 1003.785 1778.050 1004.085 ;
        RECT 1776.250 1001.635 1776.550 1003.785 ;
        RECT 1781.470 1001.635 1781.770 1004.550 ;
        RECT 1782.090 1004.550 1782.650 1006.235 ;
        RECT 1782.090 1001.635 1782.390 1004.550 ;
        RECT 1787.310 1001.635 1787.610 1007.950 ;
        RECT 1787.930 1004.850 1788.230 1006.235 ;
        RECT 1788.790 1004.850 1789.090 1015.415 ;
        RECT 1789.695 1014.735 1790.025 1015.065 ;
        RECT 1793.375 1014.735 1793.705 1015.065 ;
        RECT 1787.930 1004.550 1789.090 1004.850 ;
        RECT 1789.710 1004.850 1790.010 1014.735 ;
        RECT 1793.390 1008.250 1793.690 1014.735 ;
        RECT 1793.390 1007.950 1794.070 1008.250 ;
        RECT 1793.150 1004.850 1793.450 1006.235 ;
        RECT 1789.710 1004.550 1793.450 1004.850 ;
        RECT 1787.930 1001.635 1788.230 1004.550 ;
        RECT 1793.150 1001.635 1793.450 1004.550 ;
        RECT 1793.770 1001.635 1794.070 1007.950 ;
        RECT 1796.150 1004.850 1796.450 1020.855 ;
        RECT 1801.655 1020.175 1801.985 1020.505 ;
        RECT 1799.815 1014.735 1800.145 1015.065 ;
        RECT 1799.830 1006.235 1800.130 1014.735 ;
        RECT 1798.990 1004.850 1799.290 1006.235 ;
        RECT 1796.150 1004.550 1799.290 1004.850 ;
        RECT 1798.990 1001.635 1799.290 1004.550 ;
        RECT 1799.610 1004.550 1800.130 1006.235 ;
        RECT 1801.670 1004.850 1801.970 1020.175 ;
        RECT 1808.095 1019.495 1808.425 1019.825 ;
        RECT 1806.255 1014.735 1806.585 1015.065 ;
        RECT 1804.830 1004.850 1805.130 1006.235 ;
        RECT 1801.670 1004.550 1805.130 1004.850 ;
        RECT 1799.610 1001.635 1799.910 1004.550 ;
        RECT 1804.830 1001.635 1805.130 1004.550 ;
        RECT 1805.450 1004.850 1805.750 1006.235 ;
        RECT 1806.270 1004.850 1806.570 1014.735 ;
        RECT 1805.450 1004.550 1806.570 1004.850 ;
        RECT 1808.110 1004.850 1808.410 1019.495 ;
        RECT 1814.535 1018.815 1814.865 1019.145 ;
        RECT 1821.895 1018.815 1822.225 1019.145 ;
        RECT 1812.695 1014.735 1813.025 1015.065 ;
        RECT 1810.670 1004.850 1810.970 1006.235 ;
        RECT 1808.110 1004.550 1810.970 1004.850 ;
        RECT 1805.450 1001.635 1805.750 1004.550 ;
        RECT 1810.670 1001.635 1810.970 1004.550 ;
        RECT 1811.290 1004.085 1811.590 1006.235 ;
        RECT 1812.710 1004.085 1813.010 1014.735 ;
        RECT 1814.550 1004.850 1814.850 1018.815 ;
        RECT 1817.295 1014.735 1817.625 1015.065 ;
        RECT 1817.310 1006.235 1817.610 1014.735 ;
        RECT 1821.910 1008.250 1822.210 1018.815 ;
        RECT 1823.735 1014.735 1824.065 1015.065 ;
        RECT 1821.910 1007.950 1822.650 1008.250 ;
        RECT 1816.510 1004.850 1816.810 1006.235 ;
        RECT 1814.550 1004.550 1816.810 1004.850 ;
        RECT 1811.290 1003.785 1813.010 1004.085 ;
        RECT 1811.290 1001.635 1811.590 1003.785 ;
        RECT 1816.510 1001.635 1816.810 1004.550 ;
        RECT 1817.130 1004.550 1817.610 1006.235 ;
        RECT 1817.130 1001.635 1817.430 1004.550 ;
        RECT 1822.350 1001.635 1822.650 1007.950 ;
        RECT 1822.970 1004.850 1823.270 1006.235 ;
        RECT 1823.750 1004.850 1824.050 1014.735 ;
        RECT 1822.970 1004.550 1824.050 1004.850 ;
        RECT 1828.810 1004.850 1829.110 1006.235 ;
        RECT 1830.190 1004.850 1830.490 1020.855 ;
        RECT 1837.535 1020.175 1837.865 1020.505 ;
        RECT 1832.015 1019.495 1832.345 1019.825 ;
        RECT 1828.810 1004.550 1830.490 1004.850 ;
        RECT 1832.030 1004.850 1832.330 1019.495 ;
        RECT 1834.650 1004.850 1834.950 1006.235 ;
        RECT 1832.030 1004.550 1834.950 1004.850 ;
        RECT 1837.550 1004.850 1837.850 1020.175 ;
        RECT 1843.055 1016.095 1843.385 1016.425 ;
        RECT 1840.490 1004.850 1840.790 1006.235 ;
        RECT 1837.550 1004.550 1840.790 1004.850 ;
        RECT 1843.070 1004.850 1843.370 1016.095 ;
        RECT 1846.330 1004.850 1846.630 1006.235 ;
        RECT 1843.070 1004.550 1846.630 1004.850 ;
        RECT 1822.970 1001.635 1823.270 1004.550 ;
        RECT 1828.810 1001.635 1829.110 1004.550 ;
        RECT 1834.650 1001.635 1834.950 1004.550 ;
        RECT 1840.490 1001.635 1840.790 1004.550 ;
        RECT 1846.330 1001.635 1846.630 1004.550 ;
        RECT 1852.170 1004.850 1852.470 1006.235 ;
        RECT 1855.030 1004.850 1855.330 1020.855 ;
        RECT 2246.935 1020.175 2247.265 1020.505 ;
        RECT 2241.415 1018.815 2241.745 1019.145 ;
        RECT 2241.430 1008.250 2241.730 1018.815 ;
        RECT 1852.170 1004.550 1855.330 1004.850 ;
        RECT 2241.310 1007.950 2241.730 1008.250 ;
        RECT 1852.170 1001.635 1852.470 1004.550 ;
        RECT 2241.310 1001.635 2241.610 1007.950 ;
        RECT 2241.915 1007.255 2242.245 1007.585 ;
        RECT 2241.930 1001.635 2242.230 1007.255 ;
        RECT 2246.950 1006.235 2247.250 1020.175 ;
        RECT 2247.855 1016.775 2248.185 1017.105 ;
        RECT 2254.295 1016.775 2254.625 1017.105 ;
        RECT 2260.735 1016.775 2261.065 1017.105 ;
        RECT 2266.255 1016.775 2266.585 1017.105 ;
        RECT 2280.055 1016.775 2280.385 1017.105 ;
        RECT 2247.870 1006.235 2248.170 1016.775 ;
        RECT 2253.375 1016.095 2253.705 1016.425 ;
        RECT 2253.390 1008.250 2253.690 1016.095 ;
        RECT 2246.950 1004.550 2247.450 1006.235 ;
        RECT 2247.150 1001.635 2247.450 1004.550 ;
        RECT 2247.770 1004.550 2248.170 1006.235 ;
        RECT 2252.990 1007.950 2253.690 1008.250 ;
        RECT 2247.770 1001.635 2248.070 1004.550 ;
        RECT 2252.990 1001.635 2253.290 1007.950 ;
        RECT 2253.610 1004.850 2253.910 1006.235 ;
        RECT 2254.310 1004.850 2254.610 1016.775 ;
        RECT 2258.895 1014.735 2259.225 1015.065 ;
        RECT 2258.910 1008.250 2259.210 1014.735 ;
        RECT 2253.610 1004.550 2254.610 1004.850 ;
        RECT 2258.830 1007.950 2259.210 1008.250 ;
        RECT 2253.610 1001.635 2253.910 1004.550 ;
        RECT 2258.830 1001.635 2259.130 1007.950 ;
        RECT 2259.450 1004.085 2259.750 1006.235 ;
        RECT 2260.750 1004.085 2261.050 1016.775 ;
        RECT 2264.415 1016.095 2264.745 1016.425 ;
        RECT 2264.430 1006.235 2264.730 1016.095 ;
        RECT 2264.430 1004.550 2264.970 1006.235 ;
        RECT 2259.450 1003.785 2261.050 1004.085 ;
        RECT 2259.450 1001.635 2259.750 1003.785 ;
        RECT 2264.670 1001.635 2264.970 1004.550 ;
        RECT 2265.290 1004.850 2265.590 1006.235 ;
        RECT 2266.270 1004.850 2266.570 1016.775 ;
        RECT 2274.535 1016.095 2274.865 1016.425 ;
        RECT 2276.375 1016.095 2276.705 1016.425 ;
        RECT 2270.855 1014.735 2271.185 1015.065 ;
        RECT 2270.870 1008.250 2271.170 1014.735 ;
        RECT 2265.290 1004.550 2266.570 1004.850 ;
        RECT 2270.510 1007.950 2271.170 1008.250 ;
        RECT 2265.290 1001.635 2265.590 1004.550 ;
        RECT 2270.510 1001.635 2270.810 1007.950 ;
        RECT 2271.130 1004.850 2271.430 1006.235 ;
        RECT 2274.550 1004.850 2274.850 1016.095 ;
        RECT 2276.390 1008.250 2276.690 1016.095 ;
        RECT 2271.130 1004.550 2274.850 1004.850 ;
        RECT 2276.350 1007.950 2276.690 1008.250 ;
        RECT 2271.130 1001.635 2271.430 1004.550 ;
        RECT 2276.350 1001.635 2276.650 1007.950 ;
        RECT 2276.970 1004.850 2277.270 1006.235 ;
        RECT 2280.070 1004.850 2280.370 1016.775 ;
        RECT 2281.895 1014.735 2282.225 1015.065 ;
        RECT 2276.970 1004.550 2280.370 1004.850 ;
        RECT 2281.910 1006.235 2282.210 1014.735 ;
        RECT 2282.830 1006.235 2283.130 1020.855 ;
        RECT 2335.255 1020.175 2335.585 1020.505 ;
        RECT 2293.855 1016.775 2294.185 1017.105 ;
        RECT 2304.895 1016.775 2305.225 1017.105 ;
        RECT 2311.335 1016.775 2311.665 1017.105 ;
        RECT 2287.415 1016.095 2287.745 1016.425 ;
        RECT 2281.910 1004.550 2282.490 1006.235 ;
        RECT 2276.970 1001.635 2277.270 1004.550 ;
        RECT 2282.190 1001.635 2282.490 1004.550 ;
        RECT 2282.810 1004.550 2283.130 1006.235 ;
        RECT 2287.430 1004.850 2287.730 1016.095 ;
        RECT 2289.255 1014.735 2289.585 1015.065 ;
        RECT 2288.030 1004.850 2288.330 1006.235 ;
        RECT 2287.430 1004.550 2288.330 1004.850 ;
        RECT 2282.810 1001.635 2283.110 1004.550 ;
        RECT 2288.030 1001.635 2288.330 1004.550 ;
        RECT 2288.650 1004.850 2288.950 1006.235 ;
        RECT 2289.270 1004.850 2289.570 1014.735 ;
        RECT 2288.650 1004.550 2289.570 1004.850 ;
        RECT 2288.650 1001.635 2288.950 1004.550 ;
        RECT 2293.870 1001.635 2294.170 1016.775 ;
        RECT 2300.295 1016.095 2300.625 1016.425 ;
        RECT 2294.775 1014.735 2295.105 1015.065 ;
        RECT 2294.790 1006.235 2295.090 1014.735 ;
        RECT 2300.310 1008.250 2300.610 1016.095 ;
        RECT 2302.135 1014.735 2302.465 1015.065 ;
        RECT 2294.490 1004.550 2295.090 1006.235 ;
        RECT 2299.710 1007.950 2300.610 1008.250 ;
        RECT 2294.490 1001.635 2294.790 1004.550 ;
        RECT 2299.710 1001.635 2300.010 1007.950 ;
        RECT 2300.330 1004.850 2300.630 1006.235 ;
        RECT 2302.150 1004.850 2302.450 1014.735 ;
        RECT 2300.330 1004.550 2302.450 1004.850 ;
        RECT 2304.910 1004.850 2305.210 1016.775 ;
        RECT 2307.655 1014.735 2307.985 1015.065 ;
        RECT 2305.550 1004.850 2305.850 1006.235 ;
        RECT 2304.910 1004.550 2305.850 1004.850 ;
        RECT 2300.330 1001.635 2300.630 1004.550 ;
        RECT 2305.550 1001.635 2305.850 1004.550 ;
        RECT 2306.170 1004.085 2306.470 1006.235 ;
        RECT 2307.670 1004.085 2307.970 1014.735 ;
        RECT 2311.350 1006.235 2311.650 1016.775 ;
        RECT 2315.935 1016.095 2316.265 1016.425 ;
        RECT 2323.295 1016.095 2323.625 1016.425 ;
        RECT 2329.735 1016.095 2330.065 1016.425 ;
        RECT 2312.255 1014.735 2312.585 1015.065 ;
        RECT 2312.270 1006.235 2312.570 1014.735 ;
        RECT 2311.350 1004.550 2311.690 1006.235 ;
        RECT 2306.170 1003.785 2307.970 1004.085 ;
        RECT 2306.170 1001.635 2306.470 1003.785 ;
        RECT 2311.390 1001.635 2311.690 1004.550 ;
        RECT 2312.010 1004.550 2312.570 1006.235 ;
        RECT 2312.010 1001.635 2312.310 1004.550 ;
        RECT 2315.950 1004.085 2316.250 1016.095 ;
        RECT 2317.775 1014.735 2318.105 1015.065 ;
        RECT 2322.375 1014.735 2322.705 1015.065 ;
        RECT 2317.790 1008.250 2318.090 1014.735 ;
        RECT 2317.790 1007.950 2318.150 1008.250 ;
        RECT 2317.230 1004.085 2317.530 1006.235 ;
        RECT 2315.950 1003.785 2317.530 1004.085 ;
        RECT 2317.230 1001.635 2317.530 1003.785 ;
        RECT 2317.850 1001.635 2318.150 1007.950 ;
        RECT 2322.390 1004.850 2322.690 1014.735 ;
        RECT 2323.310 1008.250 2323.610 1016.095 ;
        RECT 2328.815 1014.735 2329.145 1015.065 ;
        RECT 2323.310 1007.950 2323.990 1008.250 ;
        RECT 2323.070 1004.850 2323.370 1006.235 ;
        RECT 2322.390 1004.550 2323.370 1004.850 ;
        RECT 2323.070 1001.635 2323.370 1004.550 ;
        RECT 2323.690 1001.635 2323.990 1007.950 ;
        RECT 2328.830 1006.235 2329.130 1014.735 ;
        RECT 2329.750 1006.235 2330.050 1016.095 ;
        RECT 2335.270 1008.250 2335.570 1020.175 ;
        RECT 2336.175 1014.735 2336.505 1015.065 ;
        RECT 2328.830 1004.550 2329.210 1006.235 ;
        RECT 2328.910 1001.635 2329.210 1004.550 ;
        RECT 2329.530 1004.550 2330.050 1006.235 ;
        RECT 2334.750 1007.950 2335.570 1008.250 ;
        RECT 2329.530 1001.635 2329.830 1004.550 ;
        RECT 2334.750 1001.635 2335.050 1007.950 ;
        RECT 2335.370 1004.850 2335.670 1006.235 ;
        RECT 2336.190 1004.850 2336.490 1014.735 ;
        RECT 2340.790 1008.250 2341.090 1020.855 ;
        RECT 2346.295 1020.175 2346.625 1020.505 ;
        RECT 2342.615 1014.735 2342.945 1015.065 ;
        RECT 2335.370 1004.550 2336.490 1004.850 ;
        RECT 2340.590 1007.950 2341.090 1008.250 ;
        RECT 2335.370 1001.635 2335.670 1004.550 ;
        RECT 2340.590 1001.635 2340.890 1007.950 ;
        RECT 2341.210 1004.085 2341.510 1006.235 ;
        RECT 2342.630 1004.085 2342.930 1014.735 ;
        RECT 2346.310 1006.235 2346.610 1020.175 ;
        RECT 2347.215 1014.735 2347.545 1015.065 ;
        RECT 2347.230 1006.235 2347.530 1014.735 ;
        RECT 2351.830 1008.250 2352.130 1020.855 ;
        RECT 2358.255 1016.095 2358.585 1016.425 ;
        RECT 2363.775 1016.095 2364.105 1016.425 ;
        RECT 2353.655 1014.735 2353.985 1015.065 ;
        RECT 2351.830 1007.950 2352.570 1008.250 ;
        RECT 2346.310 1004.550 2346.730 1006.235 ;
        RECT 2341.210 1003.785 2342.930 1004.085 ;
        RECT 2341.210 1001.635 2341.510 1003.785 ;
        RECT 2346.430 1001.635 2346.730 1004.550 ;
        RECT 2347.050 1004.550 2347.530 1006.235 ;
        RECT 2347.050 1001.635 2347.350 1004.550 ;
        RECT 2352.270 1001.635 2352.570 1007.950 ;
        RECT 2352.890 1004.850 2353.190 1006.235 ;
        RECT 2353.670 1004.850 2353.970 1014.735 ;
        RECT 2358.270 1008.250 2358.570 1016.095 ;
        RECT 2359.175 1014.735 2359.505 1015.065 ;
        RECT 2352.890 1004.550 2353.970 1004.850 ;
        RECT 2358.110 1007.950 2358.570 1008.250 ;
        RECT 2359.190 1008.250 2359.490 1014.735 ;
        RECT 2359.190 1007.950 2360.410 1008.250 ;
        RECT 2352.890 1001.635 2353.190 1004.550 ;
        RECT 2358.110 1001.635 2358.410 1007.950 ;
        RECT 2358.730 1004.085 2359.030 1006.235 ;
        RECT 2360.110 1004.085 2360.410 1007.950 ;
        RECT 2363.790 1006.235 2364.090 1016.095 ;
        RECT 2364.695 1014.735 2365.025 1015.065 ;
        RECT 2364.710 1006.235 2365.010 1014.735 ;
        RECT 2370.230 1008.250 2370.530 1038.535 ;
        RECT 2452.020 1021.235 2455.020 1185.000 ;
        RECT 2387.695 1020.855 2388.025 1021.185 ;
        RECT 2395.975 1020.855 2396.305 1021.185 ;
        RECT 2408.855 1020.855 2409.185 1021.185 ;
        RECT 2451.175 1020.855 2451.505 1021.185 ;
        RECT 2381.255 1020.175 2381.585 1020.505 ;
        RECT 2375.735 1016.095 2376.065 1016.425 ;
        RECT 2371.135 1014.735 2371.465 1015.065 ;
        RECT 2363.790 1004.550 2364.250 1006.235 ;
        RECT 2358.730 1003.785 2360.410 1004.085 ;
        RECT 2358.730 1001.635 2359.030 1003.785 ;
        RECT 2363.950 1001.635 2364.250 1004.550 ;
        RECT 2364.570 1004.550 2365.010 1006.235 ;
        RECT 2369.790 1007.950 2370.530 1008.250 ;
        RECT 2364.570 1001.635 2364.870 1004.550 ;
        RECT 2369.790 1001.635 2370.090 1007.950 ;
        RECT 2370.410 1004.850 2370.710 1006.235 ;
        RECT 2371.150 1004.850 2371.450 1014.735 ;
        RECT 2375.750 1008.250 2376.050 1016.095 ;
        RECT 2377.575 1014.735 2377.905 1015.065 ;
        RECT 2370.410 1004.550 2371.450 1004.850 ;
        RECT 2375.630 1007.950 2376.050 1008.250 ;
        RECT 2370.410 1001.635 2370.710 1004.550 ;
        RECT 2375.630 1001.635 2375.930 1007.950 ;
        RECT 2376.250 1004.085 2376.550 1006.235 ;
        RECT 2377.590 1004.085 2377.890 1014.735 ;
        RECT 2381.270 1006.235 2381.570 1020.175 ;
        RECT 2382.175 1014.735 2382.505 1015.065 ;
        RECT 2382.190 1006.235 2382.490 1014.735 ;
        RECT 2387.710 1007.570 2388.010 1020.855 ;
        RECT 2390.455 1020.175 2390.785 1020.505 ;
        RECT 2388.615 1016.095 2388.945 1016.425 ;
        RECT 2381.270 1004.550 2381.770 1006.235 ;
        RECT 2376.250 1003.785 2377.890 1004.085 ;
        RECT 2376.250 1001.635 2376.550 1003.785 ;
        RECT 2381.470 1001.635 2381.770 1004.550 ;
        RECT 2382.090 1004.550 2382.490 1006.235 ;
        RECT 2387.310 1007.270 2388.010 1007.570 ;
        RECT 2382.090 1001.635 2382.390 1004.550 ;
        RECT 2387.310 1001.635 2387.610 1007.270 ;
        RECT 2387.930 1004.850 2388.230 1006.235 ;
        RECT 2388.630 1004.850 2388.930 1016.095 ;
        RECT 2387.930 1004.550 2388.930 1004.850 ;
        RECT 2390.470 1004.850 2390.770 1020.175 ;
        RECT 2393.215 1016.775 2393.545 1017.105 ;
        RECT 2393.230 1007.570 2393.530 1016.775 ;
        RECT 2393.230 1007.270 2394.070 1007.570 ;
        RECT 2393.150 1004.850 2393.450 1006.235 ;
        RECT 2390.470 1004.550 2393.450 1004.850 ;
        RECT 2387.930 1001.635 2388.230 1004.550 ;
        RECT 2393.150 1001.635 2393.450 1004.550 ;
        RECT 2393.770 1001.635 2394.070 1007.270 ;
        RECT 2395.990 1004.850 2396.290 1020.855 ;
        RECT 2402.415 1019.495 2402.745 1019.825 ;
        RECT 2399.655 1014.735 2399.985 1015.065 ;
        RECT 2399.670 1006.235 2399.970 1014.735 ;
        RECT 2398.990 1004.850 2399.290 1006.235 ;
        RECT 2395.990 1004.550 2399.290 1004.850 ;
        RECT 2398.990 1001.635 2399.290 1004.550 ;
        RECT 2399.610 1004.550 2399.970 1006.235 ;
        RECT 2402.430 1004.850 2402.730 1019.495 ;
        RECT 2406.095 1014.735 2406.425 1015.065 ;
        RECT 2404.830 1004.850 2405.130 1006.235 ;
        RECT 2402.430 1004.550 2405.130 1004.850 ;
        RECT 2399.610 1001.635 2399.910 1004.550 ;
        RECT 2404.830 1001.635 2405.130 1004.550 ;
        RECT 2405.450 1004.850 2405.750 1006.235 ;
        RECT 2406.110 1004.850 2406.410 1014.735 ;
        RECT 2405.450 1004.550 2406.410 1004.850 ;
        RECT 2408.870 1004.850 2409.170 1020.855 ;
        RECT 2429.095 1020.175 2429.425 1020.505 ;
        RECT 2415.295 1018.135 2415.625 1018.465 ;
        RECT 2410.695 1014.735 2411.025 1015.065 ;
        RECT 2410.710 1008.250 2411.010 1014.735 ;
        RECT 2410.710 1007.950 2411.590 1008.250 ;
        RECT 2410.670 1004.850 2410.970 1006.235 ;
        RECT 2408.870 1004.550 2410.970 1004.850 ;
        RECT 2405.450 1001.635 2405.750 1004.550 ;
        RECT 2410.670 1001.635 2410.970 1004.550 ;
        RECT 2411.290 1001.635 2411.590 1007.950 ;
        RECT 2415.310 1004.850 2415.610 1018.135 ;
        RECT 2421.735 1017.455 2422.065 1017.785 ;
        RECT 2417.135 1014.735 2417.465 1015.065 ;
        RECT 2417.150 1006.235 2417.450 1014.735 ;
        RECT 2416.510 1004.850 2416.810 1006.235 ;
        RECT 2415.310 1004.550 2416.810 1004.850 ;
        RECT 2416.510 1001.635 2416.810 1004.550 ;
        RECT 2417.130 1004.550 2417.450 1006.235 ;
        RECT 2421.750 1004.850 2422.050 1017.455 ;
        RECT 2423.575 1014.735 2423.905 1015.065 ;
        RECT 2422.350 1004.850 2422.650 1006.235 ;
        RECT 2421.750 1004.550 2422.650 1004.850 ;
        RECT 2417.130 1001.635 2417.430 1004.550 ;
        RECT 2422.350 1001.635 2422.650 1004.550 ;
        RECT 2422.970 1004.850 2423.270 1006.235 ;
        RECT 2423.590 1004.850 2423.890 1014.735 ;
        RECT 2429.110 1006.235 2429.410 1020.175 ;
        RECT 2437.375 1018.135 2437.705 1018.465 ;
        RECT 2431.855 1016.095 2432.185 1016.425 ;
        RECT 2422.970 1004.550 2423.890 1004.850 ;
        RECT 2428.810 1004.550 2429.410 1006.235 ;
        RECT 2431.870 1004.850 2432.170 1016.095 ;
        RECT 2434.650 1004.850 2434.950 1006.235 ;
        RECT 2431.870 1004.550 2434.950 1004.850 ;
        RECT 2437.390 1004.850 2437.690 1018.135 ;
        RECT 2442.895 1017.455 2443.225 1017.785 ;
        RECT 2440.490 1004.850 2440.790 1006.235 ;
        RECT 2437.390 1004.550 2440.790 1004.850 ;
        RECT 2442.910 1004.850 2443.210 1017.455 ;
        RECT 2446.330 1004.850 2446.630 1006.235 ;
        RECT 2442.910 1004.550 2446.630 1004.850 ;
        RECT 2451.190 1004.850 2451.490 1020.855 ;
        RECT 2452.170 1004.850 2452.470 1006.235 ;
        RECT 2451.190 1004.550 2452.470 1004.850 ;
        RECT 2422.970 1001.635 2423.270 1004.550 ;
        RECT 2428.810 1001.635 2429.110 1004.550 ;
        RECT 2434.650 1001.635 2434.950 1004.550 ;
        RECT 2440.490 1001.635 2440.790 1004.550 ;
        RECT 2446.330 1001.635 2446.630 1004.550 ;
        RECT 2452.170 1001.635 2452.470 1004.550 ;
      LAYER met4 ;
        RECT 1505.000 555.000 1881.480 1001.235 ;
        RECT 2105.000 555.000 2481.480 1001.235 ;
      LAYER met4 ;
        RECT 1598.715 550.000 1599.015 554.600 ;
        RECT 1604.955 550.000 1605.255 554.600 ;
        RECT 1611.195 550.000 1611.495 554.600 ;
        RECT 1617.435 550.000 1617.735 554.600 ;
        RECT 1623.675 550.000 1623.975 554.600 ;
        RECT 1629.915 550.000 1630.215 554.600 ;
        RECT 1636.155 550.000 1636.455 554.600 ;
        RECT 1642.395 550.000 1642.695 554.600 ;
        RECT 1648.635 550.000 1648.935 554.600 ;
        RECT 1654.875 550.000 1655.175 554.600 ;
        RECT 1661.115 550.000 1661.415 554.600 ;
        RECT 1667.355 550.000 1667.655 554.600 ;
        RECT 1673.595 550.000 1673.895 554.600 ;
        RECT 1679.835 550.000 1680.135 554.600 ;
        RECT 1686.075 550.000 1686.375 554.600 ;
        RECT 1692.315 550.000 1692.615 554.600 ;
        RECT 1698.555 550.000 1698.855 554.600 ;
        RECT 1704.795 550.000 1705.095 554.600 ;
        RECT 1711.035 550.000 1711.335 554.600 ;
        RECT 1717.275 550.000 1717.575 554.600 ;
        RECT 1723.515 550.000 1723.815 554.600 ;
        RECT 1729.755 550.000 1730.055 554.600 ;
        RECT 1735.995 550.000 1736.295 554.600 ;
        RECT 1742.235 550.000 1742.535 554.600 ;
        RECT 1748.475 550.000 1748.775 554.600 ;
        RECT 1754.715 550.000 1755.015 554.600 ;
        RECT 1760.955 550.000 1761.255 554.600 ;
        RECT 1767.195 550.000 1767.495 554.600 ;
        RECT 1773.435 550.000 1773.735 554.600 ;
        RECT 1779.675 550.000 1779.975 554.600 ;
        RECT 1785.915 550.000 1786.215 554.600 ;
        RECT 1792.155 550.000 1792.455 554.600 ;
        RECT 2198.715 550.000 2199.015 554.600 ;
        RECT 2204.955 550.000 2205.255 554.600 ;
        RECT 2211.195 550.000 2211.495 554.600 ;
        RECT 2217.435 550.000 2217.735 554.600 ;
        RECT 2223.675 550.000 2223.975 554.600 ;
        RECT 2229.915 550.000 2230.215 554.600 ;
        RECT 2236.155 550.000 2236.455 554.600 ;
        RECT 2242.395 550.000 2242.695 554.600 ;
        RECT 2248.635 550.000 2248.935 554.600 ;
        RECT 2254.875 550.000 2255.175 554.600 ;
        RECT 2261.115 550.000 2261.415 554.600 ;
        RECT 2267.355 550.000 2267.655 554.600 ;
        RECT 2273.595 550.000 2273.895 554.600 ;
        RECT 2279.835 550.000 2280.135 554.600 ;
        RECT 2286.075 550.000 2286.375 554.600 ;
        RECT 2292.315 550.000 2292.615 554.600 ;
        RECT 2298.555 550.000 2298.855 554.600 ;
        RECT 2304.795 550.000 2305.095 554.600 ;
        RECT 2311.035 550.000 2311.335 554.600 ;
        RECT 2317.275 550.000 2317.575 554.600 ;
        RECT 2323.515 550.000 2323.815 554.600 ;
        RECT 2329.755 550.000 2330.055 554.600 ;
        RECT 2335.995 550.000 2336.295 554.600 ;
        RECT 2342.235 550.000 2342.535 554.600 ;
        RECT 2348.475 550.000 2348.775 554.600 ;
        RECT 2354.715 550.000 2355.015 554.600 ;
        RECT 2360.955 550.000 2361.255 554.600 ;
        RECT 2367.195 550.000 2367.495 554.600 ;
        RECT 2373.435 550.000 2373.735 554.600 ;
        RECT 2379.675 550.000 2379.975 554.600 ;
        RECT 2385.915 550.000 2386.215 554.600 ;
        RECT 2392.155 550.000 2392.455 554.600 ;
  END
END user_project_wrapper
END LIBRARY

